<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Michał Derewecki" version="11.75236">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="Zimowe Otwarte Mistrzostwa Polski w Pływaniu w Kategoriach MASTERS POZNAŃ 2022" course="SCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2022-12-18" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Poznań" nation="POL" />
      <POINTTABLE pointtableid="1126" name="DSV Master Performance Table" version="2022" />
      <QUALIFY from="2021-09-01" until="2022-12-15" />
      <SESSIONS>
        <SESSION date="2022-12-16" daytime="15:00" endtime="21:05" number="1">
          <EVENTS>
            <EVENT eventid="6059" daytime="15:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6060" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7133" />
                    <RANKING order="2" place="2" resultid="7501" />
                    <RANKING order="3" place="3" resultid="8483" />
                    <RANKING order="4" place="4" resultid="8184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6062" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9450" />
                    <RANKING order="2" place="2" resultid="7789" />
                    <RANKING order="3" place="3" resultid="7604" />
                    <RANKING order="4" place="4" resultid="8349" />
                    <RANKING order="5" place="5" resultid="9768" />
                    <RANKING order="6" place="6" resultid="8932" />
                    <RANKING order="7" place="7" resultid="7667" />
                    <RANKING order="8" place="8" resultid="9573" />
                    <RANKING order="9" place="9" resultid="8404" />
                    <RANKING order="10" place="10" resultid="8192" />
                    <RANKING order="11" place="11" resultid="9580" />
                    <RANKING order="12" place="12" resultid="7463" />
                    <RANKING order="13" place="13" resultid="7612" />
                    <RANKING order="14" place="14" resultid="8179" />
                    <RANKING order="15" place="15" resultid="9932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6063" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7576" />
                    <RANKING order="2" place="2" resultid="9550" />
                    <RANKING order="3" place="3" resultid="7756" />
                    <RANKING order="4" place="4" resultid="8292" />
                    <RANKING order="5" place="5" resultid="8526" />
                    <RANKING order="6" place="-1" resultid="9813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6064" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9440" />
                    <RANKING order="2" place="2" resultid="9472" />
                    <RANKING order="3" place="3" resultid="7340" />
                    <RANKING order="4" place="4" resultid="7652" />
                    <RANKING order="5" place="5" resultid="8412" />
                    <RANKING order="6" place="6" resultid="7768" />
                    <RANKING order="7" place="7" resultid="7673" />
                    <RANKING order="8" place="8" resultid="9568" />
                    <RANKING order="9" place="-1" resultid="7902" />
                    <RANKING order="10" place="-1" resultid="8078" />
                    <RANKING order="11" place="-1" resultid="8660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6065" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9193" />
                    <RANKING order="2" place="2" resultid="6944" />
                    <RANKING order="3" place="3" resultid="8805" />
                    <RANKING order="4" place="4" resultid="9873" />
                    <RANKING order="5" place="5" resultid="9556" />
                    <RANKING order="6" place="6" resultid="8591" />
                    <RANKING order="7" place="7" resultid="9201" />
                    <RANKING order="8" place="8" resultid="9479" />
                    <RANKING order="9" place="9" resultid="9257" />
                    <RANKING order="10" place="-1" resultid="8084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6066" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8417" />
                    <RANKING order="2" place="2" resultid="8313" />
                    <RANKING order="3" place="3" resultid="8210" />
                    <RANKING order="4" place="4" resultid="9234" />
                    <RANKING order="5" place="5" resultid="9266" />
                    <RANKING order="6" place="6" resultid="9243" />
                    <RANKING order="7" place="7" resultid="8992" />
                    <RANKING order="8" place="8" resultid="9001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6067" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9273" />
                    <RANKING order="2" place="2" resultid="8547" />
                    <RANKING order="3" place="3" resultid="7350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6068" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8009" />
                    <RANKING order="2" place="2" resultid="8798" />
                    <RANKING order="3" place="3" resultid="7763" />
                    <RANKING order="4" place="4" resultid="9786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6069" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9249" />
                    <RANKING order="2" place="2" resultid="8048" />
                    <RANKING order="3" place="3" resultid="7307" />
                    <RANKING order="4" place="4" resultid="8152" />
                    <RANKING order="5" place="5" resultid="8317" />
                    <RANKING order="6" place="6" resultid="8147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6070" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9007" />
                    <RANKING order="2" place="2" resultid="7103" />
                    <RANKING order="3" place="3" resultid="6964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6071" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7931" />
                    <RANKING order="2" place="2" resultid="7544" />
                    <RANKING order="3" place="3" resultid="9465" />
                    <RANKING order="4" place="4" resultid="7536" />
                    <RANKING order="5" place="5" resultid="9563" />
                    <RANKING order="6" place="6" resultid="7381" />
                    <RANKING order="7" place="7" resultid="7368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6072" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7388" />
                    <RANKING order="2" place="2" resultid="7160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6073" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6074" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6075" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6076" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11393" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11394" daytime="15:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11395" daytime="15:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11396" daytime="15:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11397" daytime="15:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11398" daytime="15:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11399" daytime="15:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11400" daytime="15:12" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11401" daytime="15:12" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6077" daytime="15:14" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6078" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8922" />
                    <RANKING order="2" place="1" resultid="8941" />
                    <RANKING order="3" place="3" resultid="8466" />
                    <RANKING order="4" place="4" resultid="7189" />
                    <RANKING order="5" place="5" resultid="8473" />
                    <RANKING order="6" place="-1" resultid="7987" />
                    <RANKING order="7" place="-1" resultid="8794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6079" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9218" />
                    <RANKING order="2" place="2" resultid="7844" />
                    <RANKING order="3" place="3" resultid="9027" />
                    <RANKING order="4" place="4" resultid="8986" />
                    <RANKING order="5" place="5" resultid="6974" />
                    <RANKING order="6" place="6" resultid="9775" />
                    <RANKING order="7" place="7" resultid="7595" />
                    <RANKING order="8" place="8" resultid="8824" />
                    <RANKING order="9" place="9" resultid="8818" />
                    <RANKING order="10" place="10" resultid="9722" />
                    <RANKING order="11" place="11" resultid="7646" />
                    <RANKING order="12" place="12" resultid="8424" />
                    <RANKING order="13" place="13" resultid="8534" />
                    <RANKING order="14" place="14" resultid="6799" />
                    <RANKING order="15" place="15" resultid="7621" />
                    <RANKING order="16" place="16" resultid="7143" />
                    <RANKING order="17" place="17" resultid="9746" />
                    <RANKING order="18" place="18" resultid="9605" />
                    <RANKING order="19" place="19" resultid="7123" />
                    <RANKING order="20" place="20" resultid="7249" />
                    <RANKING order="21" place="21" resultid="8397" />
                    <RANKING order="22" place="-1" resultid="8169" />
                    <RANKING order="23" place="-1" resultid="8500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6080" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9781" />
                    <RANKING order="2" place="2" resultid="9737" />
                    <RANKING order="3" place="3" resultid="8363" />
                    <RANKING order="4" place="4" resultid="9677" />
                    <RANKING order="5" place="5" resultid="9021" />
                    <RANKING order="6" place="6" resultid="8173" />
                    <RANKING order="7" place="7" resultid="8599" />
                    <RANKING order="8" place="8" resultid="11345" />
                    <RANKING order="9" place="9" resultid="8269" />
                    <RANKING order="10" place="10" resultid="7071" />
                    <RANKING order="11" place="11" resultid="8727" />
                    <RANKING order="12" place="12" resultid="7357" />
                    <RANKING order="13" place="13" resultid="8391" />
                    <RANKING order="14" place="14" resultid="9132" />
                    <RANKING order="15" place="15" resultid="7234" />
                    <RANKING order="16" place="16" resultid="9795" />
                    <RANKING order="17" place="-1" resultid="7291" />
                    <RANKING order="18" place="-1" resultid="8190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6081" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9798" />
                    <RANKING order="2" place="2" resultid="6961" />
                    <RANKING order="3" place="3" resultid="11364" />
                    <RANKING order="4" place="4" resultid="7430" />
                    <RANKING order="5" place="5" resultid="9115" />
                    <RANKING order="6" place="6" resultid="7974" />
                    <RANKING order="7" place="7" resultid="9617" />
                    <RANKING order="8" place="8" resultid="7283" />
                    <RANKING order="9" place="9" resultid="7472" />
                    <RANKING order="10" place="10" resultid="9140" />
                    <RANKING order="11" place="11" resultid="8669" />
                    <RANKING order="12" place="12" resultid="8245" />
                    <RANKING order="13" place="13" resultid="6915" />
                    <RANKING order="14" place="14" resultid="8377" />
                    <RANKING order="15" place="15" resultid="8515" />
                    <RANKING order="16" place="16" resultid="7927" />
                    <RANKING order="17" place="17" resultid="9319" />
                    <RANKING order="18" place="-1" resultid="7477" />
                    <RANKING order="19" place="-1" resultid="6907" />
                    <RANKING order="20" place="-1" resultid="8384" />
                    <RANKING order="21" place="-1" resultid="9593" />
                    <RANKING order="22" place="-1" resultid="9690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6082" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9585" />
                    <RANKING order="2" place="2" resultid="7702" />
                    <RANKING order="3" place="3" resultid="9032" />
                    <RANKING order="4" place="4" resultid="6951" />
                    <RANKING order="5" place="5" resultid="8813" />
                    <RANKING order="6" place="6" resultid="7939" />
                    <RANKING order="7" place="7" resultid="9296" />
                    <RANKING order="8" place="8" resultid="11381" />
                    <RANKING order="9" place="9" resultid="9430" />
                    <RANKING order="10" place="10" resultid="7967" />
                    <RANKING order="11" place="11" resultid="8616" />
                    <RANKING order="12" place="12" resultid="9626" />
                    <RANKING order="13" place="13" resultid="8638" />
                    <RANKING order="14" place="14" resultid="8722" />
                    <RANKING order="15" place="15" resultid="7014" />
                    <RANKING order="16" place="16" resultid="11391" />
                    <RANKING order="17" place="17" resultid="9684" />
                    <RANKING order="18" place="18" resultid="8506" />
                    <RANKING order="19" place="19" resultid="9753" />
                    <RANKING order="20" place="20" resultid="9338" />
                    <RANKING order="21" place="21" resultid="8629" />
                    <RANKING order="22" place="-1" resultid="7199" />
                    <RANKING order="23" place="-1" resultid="7861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6083" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7661" />
                    <RANKING order="2" place="2" resultid="8708" />
                    <RANKING order="3" place="3" resultid="9639" />
                    <RANKING order="4" place="4" resultid="7331" />
                    <RANKING order="5" place="5" resultid="9847" />
                    <RANKING order="6" place="6" resultid="9109" />
                    <RANKING order="7" place="7" resultid="8809" />
                    <RANKING order="8" place="8" resultid="7996" />
                    <RANKING order="9" place="9" resultid="7749" />
                    <RANKING order="10" place="10" resultid="9733" />
                    <RANKING order="11" place="11" resultid="7177" />
                    <RANKING order="12" place="12" resultid="7322" />
                    <RANKING order="13" place="13" resultid="7454" />
                    <RANKING order="14" place="13" resultid="8205" />
                    <RANKING order="15" place="15" resultid="9598" />
                    <RANKING order="16" place="16" resultid="9287" />
                    <RANKING order="17" place="17" resultid="8699" />
                    <RANKING order="18" place="18" resultid="8372" />
                    <RANKING order="19" place="19" resultid="8716" />
                    <RANKING order="20" place="20" resultid="9313" />
                    <RANKING order="21" place="21" resultid="9208" />
                    <RANKING order="22" place="22" resultid="8132" />
                    <RANKING order="23" place="-1" resultid="6934" />
                    <RANKING order="24" place="-1" resultid="7222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6084" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8063" />
                    <RANKING order="2" place="2" resultid="8867" />
                    <RANKING order="3" place="3" resultid="9101" />
                    <RANKING order="4" place="4" resultid="8958" />
                    <RANKING order="5" place="5" resultid="6998" />
                    <RANKING order="6" place="6" resultid="8273" />
                    <RANKING order="7" place="7" resultid="8732" />
                    <RANKING order="8" place="8" resultid="7780" />
                    <RANKING order="9" place="-1" resultid="6987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6085" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6789" />
                    <RANKING order="2" place="2" resultid="8647" />
                    <RANKING order="3" place="3" resultid="7682" />
                    <RANKING order="4" place="4" resultid="9014" />
                    <RANKING order="5" place="5" resultid="7298" />
                    <RANKING order="6" place="6" resultid="8462" />
                    <RANKING order="7" place="7" resultid="9841" />
                    <RANKING order="8" place="8" resultid="7048" />
                    <RANKING order="9" place="9" resultid="8202" />
                    <RANKING order="10" place="10" resultid="8197" />
                    <RANKING order="11" place="11" resultid="8039" />
                    <RANKING order="12" place="12" resultid="7117" />
                    <RANKING order="13" place="13" resultid="7210" />
                    <RANKING order="14" place="14" resultid="7728" />
                    <RANKING order="15" place="-1" resultid="8848" />
                    <RANKING order="16" place="-1" resultid="7870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6086" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9456" />
                    <RANKING order="2" place="2" resultid="7921" />
                    <RANKING order="3" place="3" resultid="7032" />
                    <RANKING order="4" place="4" resultid="9867" />
                    <RANKING order="5" place="5" resultid="9305" />
                    <RANKING order="6" place="6" resultid="6809" />
                    <RANKING order="7" place="7" resultid="7740" />
                    <RANKING order="8" place="8" resultid="8979" />
                    <RANKING order="9" place="9" resultid="8974" />
                    <RANKING order="10" place="10" resultid="9804" />
                    <RANKING order="11" place="11" resultid="8968" />
                    <RANKING order="12" place="12" resultid="9490" />
                    <RANKING order="13" place="13" resultid="9611" />
                    <RANKING order="14" place="14" resultid="8255" />
                    <RANKING order="15" place="-1" resultid="9631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6087" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9322" />
                    <RANKING order="2" place="2" resultid="9331" />
                    <RANKING order="3" place="3" resultid="6877" />
                    <RANKING order="4" place="4" resultid="7522" />
                    <RANKING order="5" place="5" resultid="7312" />
                    <RANKING order="6" place="6" resultid="6837" />
                    <RANKING order="7" place="-1" resultid="9421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6088" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7511" />
                    <RANKING order="2" place="2" resultid="7639" />
                    <RANKING order="3" place="3" resultid="9280" />
                    <RANKING order="4" place="4" resultid="7410" />
                    <RANKING order="5" place="5" resultid="7268" />
                    <RANKING order="6" place="-1" resultid="7586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6089" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8030" />
                    <RANKING order="2" place="2" resultid="7395" />
                    <RANKING order="3" place="3" resultid="6893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6090" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7516" />
                    <RANKING order="2" place="2" resultid="8070" />
                    <RANKING order="3" place="3" resultid="7913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6091" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6092" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6093" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11402" daytime="15:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11403" daytime="15:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11404" daytime="15:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11405" daytime="15:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11406" daytime="15:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11407" daytime="15:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11408" daytime="15:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11409" daytime="15:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11410" daytime="15:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11411" daytime="15:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11412" daytime="15:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="11413" daytime="15:32" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="11414" daytime="15:32" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="11415" daytime="15:34" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="11416" daytime="15:34" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="11417" daytime="15:36" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="11418" daytime="15:38" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="11419" daytime="15:38" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6094" daytime="15:40" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6095" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8610" />
                    <RANKING order="2" place="2" resultid="7134" />
                    <RANKING order="3" place="3" resultid="8484" />
                    <RANKING order="4" place="4" resultid="6863" />
                    <RANKING order="5" place="-1" resultid="7502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6096" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8933" />
                    <RANKING order="2" place="2" resultid="7605" />
                    <RANKING order="3" place="3" resultid="8555" />
                    <RANKING order="4" place="4" resultid="7464" />
                    <RANKING order="5" place="5" resultid="9933" />
                    <RANKING order="6" place="-1" resultid="9040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6097" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8358" />
                    <RANKING order="2" place="2" resultid="7577" />
                    <RANKING order="3" place="3" resultid="9648" />
                    <RANKING order="4" place="4" resultid="8739" />
                    <RANKING order="5" place="5" resultid="9926" />
                    <RANKING order="6" place="6" resultid="8307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6098" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7653" />
                    <RANKING order="2" place="2" resultid="9441" />
                    <RANKING order="3" place="3" resultid="7341" />
                    <RANKING order="4" place="4" resultid="8298" />
                    <RANKING order="5" place="5" resultid="8284" />
                    <RANKING order="6" place="6" resultid="8127" />
                    <RANKING order="7" place="7" resultid="7674" />
                    <RANKING order="8" place="-1" resultid="8559" />
                    <RANKING order="9" place="-1" resultid="7089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6099" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9194" />
                    <RANKING order="2" place="2" resultid="7112" />
                    <RANKING order="3" place="3" resultid="6945" />
                    <RANKING order="4" place="4" resultid="7004" />
                    <RANKING order="5" place="5" resultid="8161" />
                    <RANKING order="6" place="6" resultid="7093" />
                    <RANKING order="7" place="7" resultid="9874" />
                    <RANKING order="8" place="8" resultid="8876" />
                    <RANKING order="9" place="-1" resultid="8085" />
                    <RANKING order="10" place="-1" resultid="9258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6100" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8211" />
                    <RANKING order="2" place="2" resultid="9496" />
                    <RANKING order="3" place="3" resultid="9235" />
                    <RANKING order="4" place="4" resultid="9343" />
                    <RANKING order="5" place="5" resultid="8993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6101" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9274" />
                    <RANKING order="2" place="2" resultid="7719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6102" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6103" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9917" />
                    <RANKING order="2" place="2" resultid="8318" />
                    <RANKING order="3" place="3" resultid="8093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6104" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6105" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="6106" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6107" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6108" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6109" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6110" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11420" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11421" daytime="15:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11422" daytime="15:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11423" daytime="15:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11424" daytime="16:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6111" daytime="16:04" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6112" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9224" />
                    <RANKING order="2" place="2" resultid="8474" />
                    <RANKING order="3" place="-1" resultid="7988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6113" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7845" />
                    <RANKING order="2" place="2" resultid="9723" />
                    <RANKING order="3" place="3" resultid="8425" />
                    <RANKING order="4" place="4" resultid="7144" />
                    <RANKING order="5" place="5" resultid="7124" />
                    <RANKING order="6" place="-1" resultid="8501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6114" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9352" />
                    <RANKING order="2" place="2" resultid="9760" />
                    <RANKING order="3" place="3" resultid="8600" />
                    <RANKING order="4" place="4" resultid="7840" />
                    <RANKING order="5" place="5" resultid="11346" />
                    <RANKING order="6" place="6" resultid="8174" />
                    <RANKING order="7" place="7" resultid="7072" />
                    <RANKING order="8" place="8" resultid="9701" />
                    <RANKING order="9" place="9" resultid="7358" />
                    <RANKING order="10" place="10" resultid="8579" />
                    <RANKING order="11" place="11" resultid="6924" />
                    <RANKING order="12" place="-1" resultid="7255" />
                    <RANKING order="13" place="-1" resultid="7292" />
                    <RANKING order="14" place="-1" resultid="7834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6115" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9618" />
                    <RANKING order="2" place="2" resultid="7975" />
                    <RANKING order="3" place="3" resultid="7633" />
                    <RANKING order="4" place="4" resultid="9141" />
                    <RANKING order="5" place="5" resultid="8757" />
                    <RANKING order="6" place="6" resultid="9320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6116" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7703" />
                    <RANKING order="2" place="2" resultid="7567" />
                    <RANKING order="3" place="3" resultid="9033" />
                    <RANKING order="4" place="4" resultid="6952" />
                    <RANKING order="5" place="5" resultid="7968" />
                    <RANKING order="6" place="6" resultid="11382" />
                    <RANKING order="7" place="7" resultid="8748" />
                    <RANKING order="8" place="8" resultid="7711" />
                    <RANKING order="9" place="9" resultid="8639" />
                    <RANKING order="10" place="10" resultid="8899" />
                    <RANKING order="11" place="-1" resultid="7862" />
                    <RANKING order="12" place="-1" resultid="9297" />
                    <RANKING order="13" place="-1" resultid="9586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6117" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7041" />
                    <RANKING order="2" place="2" resultid="8264" />
                    <RANKING order="3" place="3" resultid="8892" />
                    <RANKING order="4" place="4" resultid="7332" />
                    <RANKING order="5" place="5" resultid="9655" />
                    <RANKING order="6" place="6" resultid="8017" />
                    <RANKING order="7" place="7" resultid="9288" />
                    <RANKING order="8" place="8" resultid="9209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6118" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6901" />
                    <RANKING order="2" place="2" resultid="6992" />
                    <RANKING order="3" place="3" resultid="8102" />
                    <RANKING order="4" place="4" resultid="9522" />
                    <RANKING order="5" place="5" resultid="8884" />
                    <RANKING order="6" place="6" resultid="7781" />
                    <RANKING order="7" place="7" resultid="6821" />
                    <RANKING order="8" place="-1" resultid="8829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6119" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8648" />
                    <RANKING order="2" place="2" resultid="6790" />
                    <RANKING order="3" place="3" resultid="8655" />
                    <RANKING order="4" place="4" resultid="7299" />
                    <RANKING order="5" place="5" resultid="8675" />
                    <RANKING order="6" place="6" resultid="8040" />
                    <RANKING order="7" place="7" resultid="7211" />
                    <RANKING order="8" place="8" resultid="6845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6120" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9057" />
                    <RANKING order="2" place="2" resultid="7033" />
                    <RANKING order="3" place="3" resultid="7441" />
                    <RANKING order="4" place="4" resultid="9805" />
                    <RANKING order="5" place="-1" resultid="8569" />
                    <RANKING order="6" place="-1" resultid="9306" />
                    <RANKING order="7" place="-1" resultid="9632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6121" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9323" />
                    <RANKING order="2" place="2" resultid="6878" />
                    <RANKING order="3" place="3" resultid="9332" />
                    <RANKING order="4" place="4" resultid="7424" />
                    <RANKING order="5" place="5" resultid="7151" />
                    <RANKING order="6" place="-1" resultid="7907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6122" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9661" />
                    <RANKING order="2" place="2" resultid="9281" />
                    <RANKING order="3" place="3" resultid="9048" />
                    <RANKING order="4" place="4" resultid="7022" />
                    <RANKING order="5" place="5" resultid="6828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6123" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6124" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6125" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6126" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6127" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11425" daytime="16:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11426" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11427" daytime="16:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11428" daytime="16:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11429" daytime="16:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11430" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11431" daytime="16:34" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11432" daytime="16:38" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11433" daytime="16:40" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6128" daytime="16:44" gender="X" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6129" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6130" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9864" />
                    <RANKING order="2" place="2" resultid="8236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6131" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9899" />
                    <RANKING order="2" place="2" resultid="9667" />
                    <RANKING order="3" place="3" resultid="9089" />
                    <RANKING order="4" place="4" resultid="8777" />
                    <RANKING order="5" place="5" resultid="9816" />
                    <RANKING order="6" place="6" resultid="9668" />
                    <RANKING order="7" place="7" resultid="9852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6132" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9854" />
                    <RANKING order="2" place="2" resultid="9901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6133" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9826" />
                    <RANKING order="2" place="2" resultid="9902" />
                    <RANKING order="3" place="3" resultid="8234" />
                    <RANKING order="4" place="4" resultid="8843" />
                    <RANKING order="5" place="5" resultid="8233" />
                    <RANKING order="6" place="6" resultid="9409" />
                    <RANKING order="7" place="7" resultid="9904" />
                    <RANKING order="8" place="8" resultid="9090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6134" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9408" />
                    <RANKING order="2" place="2" resultid="9518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6135" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11434" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11435" daytime="16:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11436" daytime="16:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6145" daytime="16:54" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6153" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6154" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7827" />
                    <RANKING order="2" place="2" resultid="8556" />
                    <RANKING order="3" place="3" resultid="9041" />
                    <RANKING order="4" place="4" resultid="7613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6155" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6156" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8299" />
                    <RANKING order="2" place="-1" resultid="8128" />
                    <RANKING order="3" place="-1" resultid="8661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6157" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8877" />
                    <RANKING order="2" place="-1" resultid="8592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6158" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9149" />
                    <RANKING order="2" place="-1" resultid="8835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6159" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7550" />
                    <RANKING order="2" place="2" resultid="7720" />
                    <RANKING order="3" place="3" resultid="8548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6160" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6161" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8049" />
                    <RANKING order="2" place="2" resultid="8153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6162" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="6163" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6164" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6165" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6166" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6167" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6168" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11643" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11644" daytime="17:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6169" daytime="17:28" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6170" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8923" />
                    <RANKING order="2" place="2" resultid="8942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6171" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7596" />
                    <RANKING order="2" place="2" resultid="9122" />
                    <RANKING order="3" place="3" resultid="9823" />
                    <RANKING order="4" place="-1" resultid="7622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6172" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6925" />
                    <RANKING order="2" place="-1" resultid="7235" />
                    <RANKING order="3" place="-1" resultid="7256" />
                    <RANKING order="4" place="-1" resultid="9740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6173" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8519" />
                    <RANKING order="2" place="-1" resultid="8217" />
                    <RANKING order="3" place="-1" resultid="8378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6174" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7568" />
                    <RANKING order="2" place="2" resultid="9069" />
                    <RANKING order="3" place="3" resultid="9685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6175" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8709" />
                    <RANKING order="2" place="2" resultid="9640" />
                    <RANKING order="3" place="3" resultid="8907" />
                    <RANKING order="4" place="4" resultid="8770" />
                    <RANKING order="5" place="5" resultid="7056" />
                    <RANKING order="6" place="6" resultid="9599" />
                    <RANKING order="7" place="7" resultid="7323" />
                    <RANKING order="8" place="8" resultid="9734" />
                    <RANKING order="9" place="-1" resultid="6935" />
                    <RANKING order="10" place="-1" resultid="8133" />
                    <RANKING order="11" place="-1" resultid="9314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6176" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8868" />
                    <RANKING order="2" place="2" resultid="8765" />
                    <RANKING order="3" place="3" resultid="8885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6177" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7184" />
                    <RANKING order="2" place="-1" resultid="6846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6178" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7741" />
                    <RANKING order="2" place="2" resultid="9612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6179" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7523" />
                    <RANKING order="2" place="2" resultid="6838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6180" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7640" />
                    <RANKING order="2" place="2" resultid="9359" />
                    <RANKING order="3" place="3" resultid="7411" />
                    <RANKING order="4" place="4" resultid="7023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6181" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6182" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6183" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6184" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6185" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11645" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11646" daytime="17:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11647" daytime="17:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11648" daytime="18:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11649" daytime="18:26" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6186" daytime="18:44" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6187" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6188" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="6189" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8354" />
                    <RANKING order="2" place="2" resultid="8740" />
                    <RANKING order="3" place="3" resultid="9649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6190" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7169" />
                    <RANKING order="2" place="2" resultid="8560" />
                    <RANKING order="3" place="3" resultid="9365" />
                    <RANKING order="4" place="4" resultid="8285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6191" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6192" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8694" />
                    <RANKING order="2" place="2" resultid="9344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6193" agemax="54" agemin="50" name="Kat. F" />
                <AGEGROUP agegroupid="6194" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7448" />
                    <RANKING order="2" place="2" resultid="9787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6195" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9918" />
                    <RANKING order="2" place="2" resultid="8094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6196" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="6197" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="6198" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6199" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6200" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6201" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6202" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11650" daytime="18:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11651" daytime="19:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6203" daytime="19:42" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6204" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6205" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7697" />
                    <RANKING order="2" place="2" resultid="8682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6206" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8688" />
                    <RANKING order="2" place="-1" resultid="9702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6207" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="6208" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8749" />
                    <RANKING order="2" place="2" resultid="7015" />
                    <RANKING order="3" place="3" resultid="9531" />
                    <RANKING order="4" place="4" resultid="8900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6209" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9656" />
                    <RANKING order="2" place="2" resultid="11386" />
                    <RANKING order="3" place="3" resultid="9378" />
                    <RANKING order="4" place="4" resultid="7223" />
                    <RANKING order="5" place="-1" resultid="9074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6210" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9102" />
                    <RANKING order="2" place="2" resultid="9523" />
                    <RANKING order="3" place="3" resultid="8959" />
                    <RANKING order="4" place="4" resultid="7265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6211" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="6212" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9373" />
                    <RANKING order="2" place="2" resultid="6810" />
                    <RANKING order="3" place="3" resultid="6855" />
                    <RANKING order="4" place="4" resultid="8570" />
                    <RANKING order="5" place="5" resultid="7218" />
                    <RANKING order="6" place="-1" resultid="8256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6213" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7152" />
                    <RANKING order="2" place="2" resultid="8913" />
                    <RANKING order="3" place="3" resultid="9422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6214" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9501" />
                    <RANKING order="2" place="2" resultid="9049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6215" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6216" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6217" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6218" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6219" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11652" daytime="19:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11653" daytime="20:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11654" daytime="20:34" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-12-17" daytime="08:30" endtime="12:14" number="2">
          <EVENTS>
            <EVENT eventid="6220" daytime="08:30" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6222" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9534" />
                    <RANKING order="2" place="2" resultid="8493" />
                    <RANKING order="3" place="3" resultid="7503" />
                    <RANKING order="4" place="4" resultid="8485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6223" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9451" />
                    <RANKING order="2" place="2" resultid="8193" />
                    <RANKING order="3" place="3" resultid="8228" />
                    <RANKING order="4" place="4" resultid="9574" />
                    <RANKING order="5" place="5" resultid="9581" />
                    <RANKING order="6" place="6" resultid="7498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6224" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9810" />
                    <RANKING order="2" place="2" resultid="8308" />
                    <RANKING order="3" place="3" resultid="8293" />
                    <RANKING order="4" place="4" resultid="8741" />
                    <RANKING order="5" place="5" resultid="8527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6225" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7654" />
                    <RANKING order="2" place="2" resultid="9442" />
                    <RANKING order="3" place="3" resultid="8300" />
                    <RANKING order="4" place="-1" resultid="8079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6226" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9195" />
                    <RANKING order="2" place="2" resultid="9437" />
                    <RANKING order="3" place="3" resultid="8086" />
                    <RANKING order="4" place="4" resultid="8162" />
                    <RANKING order="5" place="5" resultid="9480" />
                    <RANKING order="6" place="6" resultid="9202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6227" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6228" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6229" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8010" />
                    <RANKING order="2" place="2" resultid="8799" />
                    <RANKING order="3" place="3" resultid="7764" />
                    <RANKING order="4" place="4" resultid="9788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6230" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9250" />
                    <RANKING order="2" place="2" resultid="9919" />
                    <RANKING order="3" place="3" resultid="8095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6231" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9507" />
                    <RANKING order="2" place="2" resultid="6966" />
                    <RANKING order="3" place="3" resultid="7376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6232" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7537" />
                    <RANKING order="2" place="2" resultid="7382" />
                    <RANKING order="3" place="3" resultid="7369" />
                    <RANKING order="4" place="-1" resultid="7932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6233" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7389" />
                    <RANKING order="2" place="2" resultid="7161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6234" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6235" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6236" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6237" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11437" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11438" daytime="08:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11439" daytime="08:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11440" daytime="08:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11441" daytime="08:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6238" daytime="08:42" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6239" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8950" />
                    <RANKING order="2" place="2" resultid="8475" />
                    <RANKING order="3" place="3" resultid="9538" />
                    <RANKING order="4" place="4" resultid="8539" />
                    <RANKING order="5" place="-1" resultid="7989" />
                    <RANKING order="6" place="-1" resultid="8795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6240" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6975" />
                    <RANKING order="2" place="2" resultid="7735" />
                    <RANKING order="3" place="3" resultid="7846" />
                    <RANKING order="4" place="4" resultid="8819" />
                    <RANKING order="5" place="5" resultid="9179" />
                    <RANKING order="6" place="6" resultid="7145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6241" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9782" />
                    <RANKING order="2" place="2" resultid="8364" />
                    <RANKING order="3" place="3" resultid="7257" />
                    <RANKING order="4" place="4" resultid="9133" />
                    <RANKING order="5" place="5" resultid="8580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6242" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9799" />
                    <RANKING order="2" place="2" resultid="9771" />
                    <RANKING order="3" place="3" resultid="7431" />
                    <RANKING order="4" place="4" resultid="8520" />
                    <RANKING order="5" place="5" resultid="7284" />
                    <RANKING order="6" place="6" resultid="7478" />
                    <RANKING order="7" place="7" resultid="8246" />
                    <RANKING order="8" place="8" resultid="8670" />
                    <RANKING order="9" place="-1" resultid="9691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6243" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9587" />
                    <RANKING order="2" place="2" resultid="7704" />
                    <RANKING order="3" place="3" resultid="7946" />
                    <RANKING order="4" place="4" resultid="9627" />
                    <RANKING order="5" place="5" resultid="7863" />
                    <RANKING order="6" place="6" resultid="7712" />
                    <RANKING order="7" place="7" resultid="7078" />
                    <RANKING order="8" place="8" resultid="7485" />
                    <RANKING order="9" place="9" resultid="7958" />
                    <RANKING order="10" place="10" resultid="7490" />
                    <RANKING order="11" place="11" resultid="8630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6244" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7662" />
                    <RANKING order="2" place="2" resultid="9110" />
                    <RANKING order="3" place="3" resultid="7057" />
                    <RANKING order="4" place="4" resultid="9641" />
                    <RANKING order="5" place="5" resultid="8908" />
                    <RANKING order="6" place="6" resultid="8771" />
                    <RANKING order="7" place="7" resultid="9157" />
                    <RANKING order="8" place="8" resultid="7324" />
                    <RANKING order="9" place="9" resultid="7455" />
                    <RANKING order="10" place="10" resultid="8701" />
                    <RANKING order="11" place="-1" resultid="9075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6245" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8869" />
                    <RANKING order="2" place="2" resultid="6993" />
                    <RANKING order="3" place="3" resultid="8103" />
                    <RANKING order="4" place="4" resultid="8960" />
                    <RANKING order="5" place="5" resultid="8274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6246" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9015" />
                    <RANKING order="2" place="2" resultid="8463" />
                    <RANKING order="3" place="3" resultid="7118" />
                    <RANKING order="4" place="4" resultid="8849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6247" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9457" />
                    <RANKING order="2" place="2" resultid="7742" />
                    <RANKING order="3" place="3" resultid="9307" />
                    <RANKING order="4" place="4" resultid="8980" />
                    <RANKING order="5" place="5" resultid="9491" />
                    <RANKING order="6" place="6" resultid="8969" />
                    <RANKING order="7" place="-1" resultid="7922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6248" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9333" />
                    <RANKING order="2" place="2" resultid="7153" />
                    <RANKING order="3" place="3" resultid="9423" />
                    <RANKING order="4" place="4" resultid="7524" />
                    <RANKING order="5" place="5" resultid="7313" />
                    <RANKING order="6" place="-1" resultid="9324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6249" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9184" />
                    <RANKING order="2" place="2" resultid="9502" />
                    <RANKING order="3" place="3" resultid="7024" />
                    <RANKING order="4" place="4" resultid="9386" />
                    <RANKING order="5" place="-1" resultid="7587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6250" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7531" />
                    <RANKING order="2" place="2" resultid="7403" />
                    <RANKING order="3" place="3" resultid="7396" />
                    <RANKING order="4" place="4" resultid="6894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6251" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6252" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6253" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6254" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11442" daytime="08:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11443" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11444" daytime="08:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11445" daytime="08:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11446" daytime="08:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11447" daytime="08:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11448" daytime="08:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11449" daytime="08:56" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11450" daytime="08:58" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6255" daytime="09:00" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6256" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8611" />
                    <RANKING order="2" place="2" resultid="6865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6257" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9042" />
                    <RANKING order="2" place="2" resultid="7668" />
                    <RANKING order="3" place="3" resultid="9542" />
                    <RANKING order="4" place="4" resultid="7465" />
                    <RANKING order="5" place="5" resultid="9934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6258" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="6259" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9473" />
                    <RANKING order="2" place="2" resultid="7875" />
                    <RANKING order="3" place="3" resultid="9366" />
                    <RANKING order="4" place="4" resultid="7903" />
                    <RANKING order="5" place="-1" resultid="7090" />
                    <RANKING order="6" place="-1" resultid="8080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6260" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7881" />
                    <RANKING order="2" place="2" resultid="8878" />
                    <RANKING order="3" place="3" resultid="12233" />
                    <RANKING order="4" place="4" resultid="9259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6261" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9497" />
                    <RANKING order="2" place="2" resultid="9236" />
                    <RANKING order="3" place="3" resultid="9345" />
                    <RANKING order="4" place="4" resultid="7207" />
                    <RANKING order="5" place="5" resultid="8994" />
                    <RANKING order="6" place="6" resultid="9267" />
                    <RANKING order="7" place="7" resultid="9002" />
                    <RANKING order="8" place="8" resultid="9244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6262" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7721" />
                    <RANKING order="2" place="2" resultid="7351" />
                    <RANKING order="3" place="-1" resultid="7551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6263" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6264" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8154" />
                    <RANKING order="2" place="2" resultid="8319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6265" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9008" />
                    <RANKING order="2" place="2" resultid="7104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6266" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9466" />
                    <RANKING order="2" place="2" resultid="6919" />
                    <RANKING order="3" place="3" resultid="7545" />
                    <RANKING order="4" place="4" resultid="7383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6267" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6268" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6269" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6270" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6271" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11451" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11452" daytime="09:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11453" daytime="09:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11454" daytime="09:18" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6272" daytime="09:22" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6273" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9226" />
                    <RANKING order="2" place="2" resultid="8454" />
                    <RANKING order="3" place="3" resultid="8540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6274" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7698" />
                    <RANKING order="2" place="2" resultid="7125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6275" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9353" />
                    <RANKING order="2" place="2" resultid="8854" />
                    <RANKING order="3" place="3" resultid="9761" />
                    <RANKING order="4" place="4" resultid="7236" />
                    <RANKING order="5" place="-1" resultid="9703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6276" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8441" />
                    <RANKING order="2" place="2" resultid="7634" />
                    <RANKING order="3" place="3" resultid="9619" />
                    <RANKING order="4" place="4" resultid="7976" />
                    <RANKING order="5" place="5" resultid="9594" />
                    <RANKING order="6" place="6" resultid="8758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6277" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9034" />
                    <RANKING order="2" place="2" resultid="7569" />
                    <RANKING order="3" place="3" resultid="11377" />
                    <RANKING order="4" place="4" resultid="8723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6278" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8265" />
                    <RANKING order="2" place="2" resultid="9657" />
                    <RANKING order="3" place="3" resultid="7058" />
                    <RANKING order="4" place="4" resultid="8018" />
                    <RANKING order="5" place="5" resultid="8279" />
                    <RANKING order="6" place="6" resultid="7278" />
                    <RANKING order="7" place="7" resultid="8717" />
                    <RANKING order="8" place="8" resultid="9379" />
                    <RANKING order="9" place="9" resultid="9210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6279" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6902" />
                    <RANKING order="2" place="2" resultid="7854" />
                    <RANKING order="3" place="3" resultid="8104" />
                    <RANKING order="4" place="4" resultid="6999" />
                    <RANKING order="5" place="5" resultid="8886" />
                    <RANKING order="6" place="6" resultid="7782" />
                    <RANKING order="7" place="7" resultid="8002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6280" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7683" />
                    <RANKING order="2" place="2" resultid="7688" />
                    <RANKING order="3" place="3" resultid="8676" />
                    <RANKING order="4" place="4" resultid="8041" />
                    <RANKING order="5" place="5" resultid="8511" />
                    <RANKING order="6" place="6" resultid="8859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6281" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9868" />
                    <RANKING order="2" place="2" resultid="9058" />
                    <RANKING order="3" place="3" resultid="7272" />
                    <RANKING order="4" place="4" resultid="8023" />
                    <RANKING order="5" place="5" resultid="8975" />
                    <RANKING order="6" place="6" resultid="9391" />
                    <RANKING order="7" place="7" resultid="8257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6282" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6879" />
                    <RANKING order="2" place="2" resultid="7425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6283" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9662" />
                    <RANKING order="2" place="2" resultid="9360" />
                    <RANKING order="3" place="3" resultid="9050" />
                    <RANKING order="4" place="4" resultid="7412" />
                    <RANKING order="5" place="5" resultid="6829" />
                    <RANKING order="6" place="-1" resultid="7588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6284" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6285" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6286" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6287" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6288" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11455" daytime="09:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11456" daytime="09:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11457" daytime="09:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11458" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11459" daytime="09:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11460" daytime="09:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6289" daytime="09:52" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6290" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7135" />
                    <RANKING order="2" place="2" resultid="8494" />
                    <RANKING order="3" place="3" resultid="7504" />
                    <RANKING order="4" place="4" resultid="8186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6291" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7790" />
                    <RANKING order="2" place="2" resultid="8934" />
                    <RANKING order="3" place="3" resultid="7606" />
                    <RANKING order="4" place="4" resultid="8405" />
                    <RANKING order="5" place="5" resultid="9575" />
                    <RANKING order="6" place="6" resultid="7614" />
                    <RANKING order="7" place="7" resultid="9545" />
                    <RANKING order="8" place="8" resultid="8180" />
                    <RANKING order="9" place="-1" resultid="7194" />
                    <RANKING order="10" place="-1" resultid="8194" />
                    <RANKING order="11" place="-1" resultid="9582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6292" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7578" />
                    <RANKING order="2" place="2" resultid="9552" />
                    <RANKING order="3" place="3" resultid="7757" />
                    <RANKING order="4" place="4" resultid="8528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6293" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9443" />
                    <RANKING order="2" place="2" resultid="7342" />
                    <RANKING order="3" place="3" resultid="8413" />
                    <RANKING order="4" place="4" resultid="7769" />
                    <RANKING order="5" place="5" resultid="8662" />
                    <RANKING order="6" place="6" resultid="7170" />
                    <RANKING order="7" place="7" resultid="8286" />
                    <RANKING order="8" place="8" resultid="7675" />
                    <RANKING order="9" place="9" resultid="9569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6294" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6946" />
                    <RANKING order="2" place="2" resultid="8806" />
                    <RANKING order="3" place="3" resultid="9875" />
                    <RANKING order="4" place="4" resultid="9557" />
                    <RANKING order="5" place="5" resultid="8593" />
                    <RANKING order="6" place="6" resultid="9400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6295" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8418" />
                    <RANKING order="2" place="2" resultid="8314" />
                    <RANKING order="3" place="3" resultid="9268" />
                    <RANKING order="4" place="4" resultid="9245" />
                    <RANKING order="5" place="-1" resultid="8836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6296" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7552" />
                    <RANKING order="2" place="2" resultid="8325" />
                    <RANKING order="3" place="3" resultid="8331" />
                    <RANKING order="4" place="4" resultid="8549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6297" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7449" />
                    <RANKING order="2" place="2" resultid="8800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6298" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8050" />
                    <RANKING order="2" place="2" resultid="7308" />
                    <RANKING order="3" place="3" resultid="8148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6299" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9009" />
                    <RANKING order="2" place="2" resultid="6967" />
                    <RANKING order="3" place="3" resultid="7377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6300" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9565" />
                    <RANKING order="2" place="2" resultid="7538" />
                    <RANKING order="3" place="3" resultid="9467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6301" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7390" />
                    <RANKING order="2" place="2" resultid="7162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6302" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6303" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6304" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6305" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11461" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11462" daytime="09:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11463" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11464" daytime="10:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11465" daytime="10:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11466" daytime="10:06" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6306" daytime="10:08" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6307" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8943" />
                    <RANKING order="2" place="2" resultid="8924" />
                    <RANKING order="3" place="3" resultid="8951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6308" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6976" />
                    <RANKING order="2" place="2" resultid="9028" />
                    <RANKING order="3" place="3" resultid="8840" />
                    <RANKING order="4" place="4" resultid="9776" />
                    <RANKING order="5" place="5" resultid="9123" />
                    <RANKING order="6" place="6" resultid="7597" />
                    <RANKING order="7" place="7" resultid="9724" />
                    <RANKING order="8" place="8" resultid="8825" />
                    <RANKING order="9" place="9" resultid="8426" />
                    <RANKING order="10" place="10" resultid="9180" />
                    <RANKING order="11" place="11" resultid="7647" />
                    <RANKING order="12" place="12" resultid="7318" />
                    <RANKING order="13" place="13" resultid="7623" />
                    <RANKING order="14" place="14" resultid="8502" />
                    <RANKING order="15" place="15" resultid="9748" />
                    <RANKING order="16" place="16" resultid="9606" />
                    <RANKING order="17" place="17" resultid="8398" />
                    <RANKING order="18" place="-1" resultid="8683" />
                    <RANKING order="19" place="-1" resultid="8820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6309" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8365" />
                    <RANKING order="2" place="2" resultid="9022" />
                    <RANKING order="3" place="3" resultid="8175" />
                    <RANKING order="4" place="4" resultid="11347" />
                    <RANKING order="5" place="5" resultid="8601" />
                    <RANKING order="6" place="6" resultid="7073" />
                    <RANKING order="7" place="7" resultid="8728" />
                    <RANKING order="8" place="8" resultid="8450" />
                    <RANKING order="9" place="9" resultid="7359" />
                    <RANKING order="10" place="10" resultid="8392" />
                    <RANKING order="11" place="10" resultid="8689" />
                    <RANKING order="12" place="12" resultid="9741" />
                    <RANKING order="13" place="13" resultid="6926" />
                    <RANKING order="14" place="14" resultid="9796" />
                    <RANKING order="15" place="-1" resultid="7293" />
                    <RANKING order="16" place="-1" resultid="7835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6310" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9772" />
                    <RANKING order="2" place="2" resultid="9116" />
                    <RANKING order="3" place="3" resultid="9143" />
                    <RANKING order="4" place="4" resultid="9680" />
                    <RANKING order="5" place="5" resultid="8671" />
                    <RANKING order="6" place="6" resultid="6916" />
                    <RANKING order="7" place="7" resultid="8218" />
                    <RANKING order="8" place="8" resultid="8379" />
                    <RANKING order="9" place="9" resultid="7928" />
                    <RANKING order="10" place="10" resultid="8516" />
                    <RANKING order="11" place="11" resultid="7230" />
                    <RANKING order="12" place="-1" resultid="6909" />
                    <RANKING order="13" place="-1" resultid="8385" />
                    <RANKING order="14" place="-1" resultid="9692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6311" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6953" />
                    <RANKING order="2" place="2" resultid="9431" />
                    <RANKING order="3" place="3" resultid="7940" />
                    <RANKING order="4" place="4" resultid="8750" />
                    <RANKING order="5" place="5" resultid="9298" />
                    <RANKING order="6" place="6" resultid="8617" />
                    <RANKING order="7" place="7" resultid="7016" />
                    <RANKING order="8" place="8" resultid="8640" />
                    <RANKING order="9" place="9" resultid="8901" />
                    <RANKING order="10" place="10" resultid="11392" />
                    <RANKING order="11" place="11" resultid="9754" />
                    <RANKING order="12" place="12" resultid="8507" />
                    <RANKING order="13" place="13" resultid="9339" />
                    <RANKING order="14" place="14" resultid="7491" />
                    <RANKING order="15" place="15" resultid="8631" />
                    <RANKING order="16" place="-1" resultid="7083" />
                    <RANKING order="17" place="-1" resultid="7200" />
                    <RANKING order="18" place="-1" resultid="7969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6312" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9848" />
                    <RANKING order="2" place="2" resultid="9642" />
                    <RANKING order="3" place="3" resultid="7333" />
                    <RANKING order="4" place="4" resultid="7997" />
                    <RANKING order="5" place="5" resultid="7750" />
                    <RANKING order="6" place="6" resultid="7178" />
                    <RANKING order="7" place="7" resultid="8772" />
                    <RANKING order="8" place="8" resultid="9695" />
                    <RANKING order="9" place="9" resultid="9289" />
                    <RANKING order="10" place="10" resultid="7456" />
                    <RANKING order="11" place="11" resultid="8702" />
                    <RANKING order="12" place="12" resultid="8206" />
                    <RANKING order="13" place="13" resultid="6936" />
                    <RANKING order="14" place="14" resultid="9435" />
                    <RANKING order="15" place="15" resultid="9315" />
                    <RANKING order="16" place="16" resultid="8373" />
                    <RANKING order="17" place="17" resultid="8224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6313" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8064" />
                    <RANKING order="2" place="2" resultid="8870" />
                    <RANKING order="3" place="3" resultid="9103" />
                    <RANKING order="4" place="4" resultid="8434" />
                    <RANKING order="5" place="5" resultid="8275" />
                    <RANKING order="6" place="6" resultid="8733" />
                    <RANKING order="7" place="-1" resultid="6988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6314" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6791" />
                    <RANKING order="2" place="2" resultid="8649" />
                    <RANKING order="3" place="3" resultid="7300" />
                    <RANKING order="4" place="4" resultid="9842" />
                    <RANKING order="5" place="5" resultid="7119" />
                    <RANKING order="6" place="6" resultid="7871" />
                    <RANKING order="7" place="7" resultid="6847" />
                    <RANKING order="8" place="8" resultid="8850" />
                    <RANKING order="9" place="9" resultid="7729" />
                    <RANKING order="10" place="-1" resultid="7049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6315" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7923" />
                    <RANKING order="2" place="2" resultid="7034" />
                    <RANKING order="3" place="3" resultid="7743" />
                    <RANKING order="4" place="4" resultid="9308" />
                    <RANKING order="5" place="5" resultid="9613" />
                    <RANKING order="6" place="6" resultid="7243" />
                    <RANKING order="7" place="7" resultid="8258" />
                    <RANKING order="8" place="-1" resultid="8970" />
                    <RANKING order="9" place="-1" resultid="9374" />
                    <RANKING order="10" place="-1" resultid="9633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6316" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7525" />
                    <RANKING order="2" place="2" resultid="9424" />
                    <RANKING order="3" place="3" resultid="8914" />
                    <RANKING order="4" place="4" resultid="6839" />
                    <RANKING order="5" place="-1" resultid="7908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6317" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7641" />
                    <RANKING order="2" place="2" resultid="7512" />
                    <RANKING order="3" place="3" resultid="9282" />
                    <RANKING order="4" place="4" resultid="7413" />
                    <RANKING order="5" place="5" resultid="7269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6318" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8032" />
                    <RANKING order="2" place="2" resultid="7397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6319" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7517" />
                    <RANKING order="2" place="2" resultid="8072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6320" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6321" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6322" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11467" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11468" daytime="10:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11469" daytime="10:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11470" daytime="10:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11471" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11472" daytime="10:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11473" daytime="10:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11474" daytime="10:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11475" daytime="10:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11476" daytime="10:28" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11477" daytime="10:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="11478" daytime="10:32" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="11479" daytime="10:34" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6323" daytime="10:36" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6324" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7136" />
                    <RANKING order="2" place="2" resultid="8612" />
                    <RANKING order="3" place="3" resultid="8486" />
                    <RANKING order="4" place="4" resultid="9535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6325" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8935" />
                    <RANKING order="2" place="2" resultid="8350" />
                    <RANKING order="3" place="3" resultid="9043" />
                    <RANKING order="4" place="4" resultid="7791" />
                    <RANKING order="5" place="5" resultid="7607" />
                    <RANKING order="6" place="6" resultid="7669" />
                    <RANKING order="7" place="7" resultid="7466" />
                    <RANKING order="8" place="8" resultid="9081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6326" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7579" />
                    <RANKING order="2" place="2" resultid="7962" />
                    <RANKING order="3" place="3" resultid="8309" />
                    <RANKING order="4" place="4" resultid="9928" />
                    <RANKING order="5" place="5" resultid="7758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6327" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7655" />
                    <RANKING order="2" place="2" resultid="7343" />
                    <RANKING order="3" place="3" resultid="9474" />
                    <RANKING order="4" place="4" resultid="7876" />
                    <RANKING order="5" place="5" resultid="9367" />
                    <RANKING order="6" place="6" resultid="8287" />
                    <RANKING order="7" place="7" resultid="8561" />
                    <RANKING order="8" place="8" resultid="7676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6328" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9196" />
                    <RANKING order="2" place="2" resultid="6947" />
                    <RANKING order="3" place="3" resultid="7005" />
                    <RANKING order="4" place="4" resultid="7882" />
                    <RANKING order="5" place="5" resultid="8087" />
                    <RANKING order="6" place="6" resultid="8163" />
                    <RANKING order="7" place="7" resultid="9876" />
                    <RANKING order="8" place="8" resultid="8594" />
                    <RANKING order="9" place="9" resultid="9203" />
                    <RANKING order="10" place="-1" resultid="8879" />
                    <RANKING order="11" place="-1" resultid="9260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6329" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8212" />
                    <RANKING order="2" place="2" resultid="9498" />
                    <RANKING order="3" place="3" resultid="8419" />
                    <RANKING order="4" place="4" resultid="8786" />
                    <RANKING order="5" place="5" resultid="9151" />
                    <RANKING order="6" place="6" resultid="9237" />
                    <RANKING order="7" place="7" resultid="9003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6330" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9276" />
                    <RANKING order="2" place="2" resultid="7722" />
                    <RANKING order="3" place="3" resultid="8332" />
                    <RANKING order="4" place="4" resultid="8326" />
                    <RANKING order="5" place="5" resultid="8550" />
                    <RANKING order="6" place="6" resultid="8057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6331" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8011" />
                    <RANKING order="2" place="2" resultid="8138" />
                    <RANKING order="3" place="3" resultid="7765" />
                    <RANKING order="4" place="4" resultid="9789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6332" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9251" />
                    <RANKING order="2" place="2" resultid="8155" />
                    <RANKING order="3" place="3" resultid="9920" />
                    <RANKING order="4" place="4" resultid="8320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6333" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6334" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7933" />
                    <RANKING order="2" place="2" resultid="7546" />
                    <RANKING order="3" place="3" resultid="7370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6335" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6336" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6337" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6338" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6339" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11480" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11481" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11482" daytime="10:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11483" daytime="10:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11484" daytime="10:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11485" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11486" daytime="10:52" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6340" daytime="10:54" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6341" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8467" />
                    <RANKING order="2" place="2" resultid="8455" />
                    <RANKING order="3" place="3" resultid="8476" />
                    <RANKING order="4" place="4" resultid="9539" />
                    <RANKING order="5" place="5" resultid="8587" />
                    <RANKING order="6" place="-1" resultid="7990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6342" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7847" />
                    <RANKING order="2" place="2" resultid="9219" />
                    <RANKING order="3" place="3" resultid="8987" />
                    <RANKING order="4" place="4" resultid="9171" />
                    <RANKING order="5" place="5" resultid="8427" />
                    <RANKING order="6" place="6" resultid="7250" />
                    <RANKING order="7" place="7" resultid="7598" />
                    <RANKING order="8" place="8" resultid="8535" />
                    <RANKING order="9" place="9" resultid="7146" />
                    <RANKING order="10" place="10" resultid="7624" />
                    <RANKING order="11" place="11" resultid="8503" />
                    <RANKING order="12" place="12" resultid="9607" />
                    <RANKING order="13" place="-1" resultid="7126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6343" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8855" />
                    <RANKING order="2" place="2" resultid="9354" />
                    <RANKING order="3" place="3" resultid="9762" />
                    <RANKING order="4" place="4" resultid="8602" />
                    <RANKING order="5" place="5" resultid="7841" />
                    <RANKING order="6" place="6" resultid="8270" />
                    <RANKING order="7" place="7" resultid="8176" />
                    <RANKING order="8" place="8" resultid="7258" />
                    <RANKING order="9" place="9" resultid="8581" />
                    <RANKING order="10" place="10" resultid="9134" />
                    <RANKING order="11" place="11" resultid="7237" />
                    <RANKING order="12" place="-1" resultid="8729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6344" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9800" />
                    <RANKING order="2" place="2" resultid="8521" />
                    <RANKING order="3" place="3" resultid="7432" />
                    <RANKING order="4" place="4" resultid="7977" />
                    <RANKING order="5" place="5" resultid="7635" />
                    <RANKING order="6" place="6" resultid="7473" />
                    <RANKING order="7" place="7" resultid="9144" />
                    <RANKING order="8" place="8" resultid="7285" />
                    <RANKING order="9" place="9" resultid="8247" />
                    <RANKING order="10" place="10" resultid="6887" />
                    <RANKING order="11" place="11" resultid="8672" />
                    <RANKING order="12" place="12" resultid="8219" />
                    <RANKING order="13" place="-1" resultid="7479" />
                    <RANKING order="14" place="-1" resultid="9620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6345" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9588" />
                    <RANKING order="2" place="2" resultid="7705" />
                    <RANKING order="3" place="3" resultid="9035" />
                    <RANKING order="4" place="4" resultid="6954" />
                    <RANKING order="5" place="5" resultid="7970" />
                    <RANKING order="6" place="6" resultid="9299" />
                    <RANKING order="7" place="7" resultid="11383" />
                    <RANKING order="8" place="8" resultid="7947" />
                    <RANKING order="9" place="9" resultid="9461" />
                    <RANKING order="10" place="10" resultid="7713" />
                    <RANKING order="11" place="11" resultid="9628" />
                    <RANKING order="12" place="12" resultid="7067" />
                    <RANKING order="13" place="13" resultid="7959" />
                    <RANKING order="14" place="14" resultid="7486" />
                    <RANKING order="15" place="15" resultid="7079" />
                    <RANKING order="16" place="16" resultid="8902" />
                    <RANKING order="17" place="17" resultid="9686" />
                    <RANKING order="18" place="18" resultid="9755" />
                    <RANKING order="19" place="19" resultid="7227" />
                    <RANKING order="20" place="-1" resultid="7017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6346" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7042" />
                    <RANKING order="2" place="2" resultid="8893" />
                    <RANKING order="3" place="3" resultid="7334" />
                    <RANKING order="4" place="4" resultid="9111" />
                    <RANKING order="5" place="5" resultid="7998" />
                    <RANKING order="6" place="6" resultid="9600" />
                    <RANKING order="7" place="7" resultid="9158" />
                    <RANKING order="8" place="8" resultid="9290" />
                    <RANKING order="9" place="9" resultid="9380" />
                    <RANKING order="10" place="10" resultid="6937" />
                    <RANKING order="11" place="11" resultid="9211" />
                    <RANKING order="12" place="12" resultid="8225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6347" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8065" />
                    <RANKING order="2" place="2" resultid="9104" />
                    <RANKING order="3" place="3" resultid="9524" />
                    <RANKING order="4" place="4" resultid="8887" />
                    <RANKING order="5" place="5" resultid="7783" />
                    <RANKING order="6" place="6" resultid="8003" />
                    <RANKING order="7" place="7" resultid="8276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6348" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6792" />
                    <RANKING order="2" place="2" resultid="7684" />
                    <RANKING order="3" place="3" resultid="8650" />
                    <RANKING order="4" place="4" resultid="7301" />
                    <RANKING order="5" place="5" resultid="8656" />
                    <RANKING order="6" place="6" resultid="8042" />
                    <RANKING order="7" place="7" resultid="7730" />
                    <RANKING order="8" place="-1" resultid="8198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6349" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9869" />
                    <RANKING order="2" place="2" resultid="7442" />
                    <RANKING order="3" place="3" resultid="9806" />
                    <RANKING order="4" place="4" resultid="9492" />
                    <RANKING order="5" place="5" resultid="6857" />
                    <RANKING order="6" place="6" resultid="8571" />
                    <RANKING order="7" place="-1" resultid="7273" />
                    <RANKING order="8" place="-1" resultid="8981" />
                    <RANKING order="9" place="-1" resultid="9634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6350" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9334" />
                    <RANKING order="2" place="2" resultid="7314" />
                    <RANKING order="3" place="3" resultid="8144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6351" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9663" />
                    <RANKING order="2" place="2" resultid="9283" />
                    <RANKING order="3" place="-1" resultid="9051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6352" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8033" />
                    <RANKING order="2" place="2" resultid="7404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6353" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6354" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6355" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6356" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11487" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11488" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11489" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11490" daytime="11:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11491" daytime="11:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11492" daytime="11:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11493" daytime="11:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11494" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11495" daytime="11:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11496" daytime="11:14" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11497" daytime="11:16" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6357" daytime="11:18" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6358" agemax="24" agemin="20" name="Kat. 0" />
                <AGEGROUP agegroupid="6359" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7828" />
                    <RANKING order="2" place="2" resultid="7615" />
                    <RANKING order="3" place="3" resultid="9546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6360" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8742" />
                    <RANKING order="2" place="2" resultid="8355" />
                    <RANKING order="3" place="3" resultid="9650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6361" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8301" />
                    <RANKING order="2" place="2" resultid="8663" />
                    <RANKING order="3" place="3" resultid="8562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6362" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7113" />
                    <RANKING order="2" place="-1" resultid="7204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6363" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8787" />
                    <RANKING order="2" place="2" resultid="9346" />
                    <RANKING order="3" place="3" resultid="8995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6364" agemax="54" agemin="50" name="Kat. F" />
                <AGEGROUP agegroupid="6365" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="6366" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8051" />
                    <RANKING order="2" place="2" resultid="8096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6367" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="6368" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="6369" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6370" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6371" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6372" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6373" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11498" daytime="11:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11499" daytime="11:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6374" daytime="11:30" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6375" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8925" />
                    <RANKING order="2" place="2" resultid="9227" />
                    <RANKING order="3" place="3" resultid="9718" />
                    <RANKING order="4" place="4" resultid="8944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6376" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="6377" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11348" />
                    <RANKING order="2" place="2" resultid="9704" />
                    <RANKING order="3" place="3" resultid="6927" />
                    <RANKING order="4" place="-1" resultid="7836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6378" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6379" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7570" />
                    <RANKING order="2" place="2" resultid="7941" />
                    <RANKING order="3" place="3" resultid="8251" />
                    <RANKING order="4" place="4" resultid="7864" />
                    <RANKING order="5" place="5" resultid="9070" />
                    <RANKING order="6" place="6" resultid="8751" />
                    <RANKING order="7" place="-1" resultid="8641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6380" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8710" />
                    <RANKING order="2" place="2" resultid="9486" />
                    <RANKING order="3" place="3" resultid="8894" />
                    <RANKING order="4" place="4" resultid="7325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6381" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9525" />
                    <RANKING order="2" place="2" resultid="8961" />
                    <RANKING order="3" place="3" resultid="8437" />
                    <RANKING order="4" place="4" resultid="8766" />
                    <RANKING order="5" place="5" resultid="9163" />
                    <RANKING order="6" place="6" resultid="8446" />
                    <RANKING order="7" place="7" resultid="6822" />
                    <RANKING order="8" place="8" resultid="7215" />
                    <RANKING order="9" place="9" resultid="8830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6382" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8677" />
                    <RANKING order="2" place="2" resultid="7050" />
                    <RANKING order="3" place="3" resultid="7212" />
                    <RANKING order="4" place="4" resultid="8860" />
                    <RANKING order="5" place="-1" resultid="6848" />
                    <RANKING order="6" place="-1" resultid="6872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6383" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7035" />
                    <RANKING order="2" place="2" resultid="8572" />
                    <RANKING order="3" place="3" resultid="8024" />
                    <RANKING order="4" place="4" resultid="6856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6384" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6880" />
                    <RANKING order="2" place="2" resultid="7154" />
                    <RANKING order="3" place="-1" resultid="9325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6385" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7025" />
                    <RANKING order="2" place="2" resultid="6830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6386" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6387" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6388" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6389" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6390" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11500" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11501" daytime="11:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11502" daytime="11:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11503" daytime="11:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11504" daytime="11:52" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6391" daytime="11:56" gender="X" number="20" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6408" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6409" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8232" />
                    <RANKING order="2" place="2" resultid="9865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6410" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9898" />
                    <RANKING order="2" place="2" resultid="9818" />
                    <RANKING order="3" place="3" resultid="9669" />
                    <RANKING order="4" place="4" resultid="9091" />
                    <RANKING order="5" place="5" resultid="8778" />
                    <RANKING order="6" place="6" resultid="9670" />
                    <RANKING order="7" place="7" resultid="9853" />
                    <RANKING order="8" place="8" resultid="11366" />
                    <RANKING order="9" place="9" resultid="9855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6411" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9900" />
                    <RANKING order="2" place="2" resultid="9905" />
                    <RANKING order="3" place="3" resultid="7246" />
                    <RANKING order="4" place="-1" resultid="8844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6412" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9903" />
                    <RANKING order="2" place="2" resultid="9827" />
                    <RANKING order="3" place="3" resultid="8917" />
                    <RANKING order="4" place="4" resultid="9856" />
                    <RANKING order="5" place="5" resultid="8235" />
                    <RANKING order="6" place="6" resultid="9092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6413" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9410" />
                    <RANKING order="2" place="2" resultid="9828" />
                    <RANKING order="3" place="3" resultid="9851" />
                    <RANKING order="4" place="4" resultid="9519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6414" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11505" daytime="11:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11506" daytime="12:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11507" daytime="12:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-12-17" daytime="15:10" endtime="19:36" number="3">
          <EVENTS>
            <EVENT eventid="6415" daytime="15:10" gender="F" number="21" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6417" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6418" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9044" />
                    <RANKING order="2" place="2" resultid="7670" />
                    <RANKING order="3" place="3" resultid="7467" />
                    <RANKING order="4" place="4" resultid="9543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6419" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7963" />
                    <RANKING order="2" place="2" resultid="7580" />
                    <RANKING order="3" place="3" resultid="8529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6420" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9475" />
                    <RANKING order="2" place="2" resultid="7344" />
                    <RANKING order="3" place="3" resultid="7877" />
                    <RANKING order="4" place="4" resultid="9368" />
                    <RANKING order="5" place="5" resultid="7904" />
                    <RANKING order="6" place="-1" resultid="7770" />
                    <RANKING order="7" place="-1" resultid="8081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6421" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7006" />
                    <RANKING order="2" place="2" resultid="7883" />
                    <RANKING order="3" place="3" resultid="9204" />
                    <RANKING order="4" place="4" resultid="9481" />
                    <RANKING order="5" place="5" resultid="9261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6422" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9499" />
                    <RANKING order="2" place="2" resultid="9238" />
                    <RANKING order="3" place="3" resultid="7208" />
                    <RANKING order="4" place="4" resultid="9269" />
                    <RANKING order="5" place="5" resultid="8996" />
                    <RANKING order="6" place="6" resultid="9004" />
                    <RANKING order="7" place="7" resultid="9246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6423" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7723" />
                    <RANKING order="2" place="2" resultid="7352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6424" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8012" />
                    <RANKING order="2" place="2" resultid="8139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6425" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8156" />
                    <RANKING order="2" place="2" resultid="8321" />
                    <RANKING order="3" place="3" resultid="8149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6426" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9010" />
                    <RANKING order="2" place="2" resultid="7105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6427" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7934" />
                    <RANKING order="2" place="2" resultid="6920" />
                    <RANKING order="3" place="3" resultid="7547" />
                    <RANKING order="4" place="4" resultid="7384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6428" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6429" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6430" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6431" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6432" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11508" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11509" daytime="15:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11510" daytime="15:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11511" daytime="15:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11512" daytime="15:22" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6433" daytime="15:26" gender="M" number="22" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6434" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9821" />
                    <RANKING order="2" place="2" resultid="8456" />
                    <RANKING order="3" place="3" resultid="8468" />
                    <RANKING order="4" place="4" resultid="8541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6435" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8988" />
                    <RANKING order="2" place="2" resultid="9172" />
                    <RANKING order="3" place="3" resultid="7251" />
                    <RANKING order="4" place="4" resultid="8428" />
                    <RANKING order="5" place="5" resultid="7127" />
                    <RANKING order="6" place="-1" resultid="8170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6436" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9175" />
                    <RANKING order="2" place="2" resultid="9355" />
                    <RANKING order="3" place="3" resultid="8856" />
                    <RANKING order="4" place="4" resultid="9763" />
                    <RANKING order="5" place="5" resultid="7238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6437" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8442" />
                    <RANKING order="2" place="2" resultid="7636" />
                    <RANKING order="3" place="3" resultid="9595" />
                    <RANKING order="4" place="4" resultid="7978" />
                    <RANKING order="5" place="5" resultid="9621" />
                    <RANKING order="6" place="6" resultid="8760" />
                    <RANKING order="7" place="7" resultid="7231" />
                    <RANKING order="8" place="-1" resultid="6888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6438" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9036" />
                    <RANKING order="2" place="2" resultid="9300" />
                    <RANKING order="3" place="3" resultid="7068" />
                    <RANKING order="4" place="4" resultid="8724" />
                    <RANKING order="5" place="5" resultid="9756" />
                    <RANKING order="6" place="6" resultid="9340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6439" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9643" />
                    <RANKING order="2" place="2" resultid="7335" />
                    <RANKING order="3" place="3" resultid="8266" />
                    <RANKING order="4" place="4" resultid="9601" />
                    <RANKING order="5" place="5" resultid="8019" />
                    <RANKING order="6" place="6" resultid="7279" />
                    <RANKING order="7" place="7" resultid="8280" />
                    <RANKING order="8" place="8" resultid="9159" />
                    <RANKING order="9" place="9" resultid="8718" />
                    <RANKING order="10" place="10" resultid="9212" />
                    <RANKING order="11" place="11" resultid="9316" />
                    <RANKING order="12" place="-1" resultid="9658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6440" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6903" />
                    <RANKING order="2" place="2" resultid="7855" />
                    <RANKING order="3" place="3" resultid="8105" />
                    <RANKING order="4" place="4" resultid="7000" />
                    <RANKING order="5" place="5" resultid="7419" />
                    <RANKING order="6" place="6" resultid="8888" />
                    <RANKING order="7" place="7" resultid="7784" />
                    <RANKING order="8" place="8" resultid="8734" />
                    <RANKING order="9" place="9" resultid="8004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6441" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7685" />
                    <RANKING order="2" place="2" resultid="8114" />
                    <RANKING order="3" place="3" resultid="8043" />
                    <RANKING order="4" place="4" resultid="8512" />
                    <RANKING order="5" place="5" resultid="7731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6442" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9870" />
                    <RANKING order="2" place="2" resultid="9059" />
                    <RANKING order="3" place="3" resultid="7443" />
                    <RANKING order="4" place="4" resultid="8976" />
                    <RANKING order="5" place="5" resultid="9309" />
                    <RANKING order="6" place="6" resultid="9392" />
                    <RANKING order="7" place="7" resultid="8025" />
                    <RANKING order="8" place="8" resultid="8259" />
                    <RANKING order="9" place="-1" resultid="7274" />
                    <RANKING order="10" place="-1" resultid="8971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6443" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7315" />
                    <RANKING order="2" place="2" resultid="6881" />
                    <RANKING order="3" place="3" resultid="7426" />
                    <RANKING order="4" place="4" resultid="9335" />
                    <RANKING order="5" place="-1" resultid="7909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6444" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9664" />
                    <RANKING order="2" place="2" resultid="9361" />
                    <RANKING order="3" place="3" resultid="7414" />
                    <RANKING order="4" place="4" resultid="9052" />
                    <RANKING order="5" place="5" resultid="9387" />
                    <RANKING order="6" place="-1" resultid="7589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6445" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7405" />
                    <RANKING order="2" place="2" resultid="7398" />
                    <RANKING order="3" place="3" resultid="6898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6446" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7917" />
                    <RANKING order="2" place="2" resultid="8073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6447" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6448" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6449" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11513" daytime="15:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11514" daytime="15:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11515" daytime="15:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11516" daytime="15:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11517" daytime="15:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11518" daytime="15:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11519" daytime="15:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11520" daytime="15:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11521" daytime="15:46" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6450" daytime="15:50" gender="F" number="23" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6451" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7137" />
                    <RANKING order="2" place="2" resultid="7505" />
                    <RANKING order="3" place="3" resultid="9536" />
                    <RANKING order="4" place="4" resultid="8487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6452" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8351" />
                    <RANKING order="2" place="2" resultid="9769" />
                    <RANKING order="3" place="3" resultid="8936" />
                    <RANKING order="4" place="4" resultid="7792" />
                    <RANKING order="5" place="5" resultid="7608" />
                    <RANKING order="6" place="6" resultid="9576" />
                    <RANKING order="7" place="7" resultid="7829" />
                    <RANKING order="8" place="8" resultid="7468" />
                    <RANKING order="9" place="9" resultid="7616" />
                    <RANKING order="10" place="-1" resultid="7195" />
                    <RANKING order="11" place="-1" resultid="8406" />
                    <RANKING order="12" place="-1" resultid="9082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6453" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8356" />
                    <RANKING order="2" place="2" resultid="7964" />
                    <RANKING order="3" place="3" resultid="9651" />
                    <RANKING order="4" place="4" resultid="8743" />
                    <RANKING order="5" place="5" resultid="8294" />
                    <RANKING order="6" place="6" resultid="8110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6454" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7656" />
                    <RANKING order="2" place="2" resultid="8302" />
                    <RANKING order="3" place="3" resultid="8664" />
                    <RANKING order="4" place="4" resultid="8414" />
                    <RANKING order="5" place="5" resultid="7878" />
                    <RANKING order="6" place="6" resultid="7677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6455" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9197" />
                    <RANKING order="2" place="2" resultid="6948" />
                    <RANKING order="3" place="3" resultid="7007" />
                    <RANKING order="4" place="4" resultid="7884" />
                    <RANKING order="5" place="5" resultid="8088" />
                    <RANKING order="6" place="6" resultid="8807" />
                    <RANKING order="7" place="7" resultid="9558" />
                    <RANKING order="8" place="8" resultid="9877" />
                    <RANKING order="9" place="9" resultid="9401" />
                    <RANKING order="10" place="-1" resultid="9205" />
                    <RANKING order="11" place="-1" resultid="9482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6456" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8213" />
                    <RANKING order="2" place="2" resultid="8315" />
                    <RANKING order="3" place="3" resultid="8788" />
                    <RANKING order="4" place="4" resultid="8420" />
                    <RANKING order="5" place="5" resultid="8997" />
                    <RANKING order="6" place="-1" resultid="8837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6457" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9277" />
                    <RANKING order="2" place="2" resultid="8058" />
                    <RANKING order="3" place="3" resultid="8333" />
                    <RANKING order="4" place="4" resultid="8327" />
                    <RANKING order="5" place="5" resultid="8551" />
                    <RANKING order="6" place="6" resultid="7353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6458" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8140" />
                    <RANKING order="2" place="2" resultid="9790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6459" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9252" />
                    <RANKING order="2" place="2" resultid="8322" />
                    <RANKING order="3" place="-1" resultid="8052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6460" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9509" />
                    <RANKING order="2" place="2" resultid="6968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6461" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7935" />
                    <RANKING order="2" place="2" resultid="7371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6462" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6463" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6464" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6465" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6466" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11522" daytime="15:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11523" daytime="15:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11524" daytime="15:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11525" daytime="15:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11526" daytime="15:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11527" daytime="15:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11528" daytime="16:00" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6467" daytime="16:00" gender="M" number="24" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6468" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8926" />
                    <RANKING order="2" place="2" resultid="7190" />
                    <RANKING order="3" place="2" resultid="8945" />
                    <RANKING order="4" place="4" resultid="8952" />
                    <RANKING order="5" place="5" resultid="8457" />
                    <RANKING order="6" place="6" resultid="9540" />
                    <RANKING order="7" place="7" resultid="8588" />
                    <RANKING order="8" place="-1" resultid="7991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6469" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9220" />
                    <RANKING order="2" place="2" resultid="7848" />
                    <RANKING order="3" place="3" resultid="9029" />
                    <RANKING order="4" place="4" resultid="7599" />
                    <RANKING order="5" place="5" resultid="8826" />
                    <RANKING order="6" place="6" resultid="8429" />
                    <RANKING order="7" place="7" resultid="9725" />
                    <RANKING order="8" place="8" resultid="7648" />
                    <RANKING order="9" place="9" resultid="8625" />
                    <RANKING order="10" place="10" resultid="8536" />
                    <RANKING order="11" place="11" resultid="7147" />
                    <RANKING order="12" place="12" resultid="7625" />
                    <RANKING order="13" place="13" resultid="7128" />
                    <RANKING order="14" place="14" resultid="9608" />
                    <RANKING order="15" place="15" resultid="8399" />
                    <RANKING order="16" place="-1" resultid="7319" />
                    <RANKING order="17" place="-1" resultid="9777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6470" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9783" />
                    <RANKING order="2" place="2" resultid="8366" />
                    <RANKING order="3" place="3" resultid="7837" />
                    <RANKING order="4" place="4" resultid="9939" />
                    <RANKING order="5" place="5" resultid="9023" />
                    <RANKING order="6" place="6" resultid="8177" />
                    <RANKING order="7" place="7" resultid="8603" />
                    <RANKING order="8" place="8" resultid="8271" />
                    <RANKING order="9" place="9" resultid="7074" />
                    <RANKING order="10" place="10" resultid="9705" />
                    <RANKING order="11" place="11" resultid="7360" />
                    <RANKING order="12" place="12" resultid="8730" />
                    <RANKING order="13" place="13" resultid="8393" />
                    <RANKING order="14" place="14" resultid="6928" />
                    <RANKING order="15" place="-1" resultid="7294" />
                    <RANKING order="16" place="-1" resultid="8582" />
                    <RANKING order="17" place="-1" resultid="11349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6471" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9801" />
                    <RANKING order="2" place="2" resultid="9117" />
                    <RANKING order="3" place="3" resultid="9085" />
                    <RANKING order="4" place="4" resultid="7286" />
                    <RANKING order="5" place="5" resultid="7979" />
                    <RANKING order="6" place="6" resultid="9514" />
                    <RANKING order="7" place="7" resultid="9145" />
                    <RANKING order="8" place="8" resultid="9681" />
                    <RANKING order="9" place="9" resultid="6889" />
                    <RANKING order="10" place="10" resultid="8761" />
                    <RANKING order="11" place="11" resultid="8220" />
                    <RANKING order="12" place="12" resultid="7929" />
                    <RANKING order="13" place="13" resultid="7232" />
                    <RANKING order="14" place="-1" resultid="6908" />
                    <RANKING order="15" place="-1" resultid="7474" />
                    <RANKING order="16" place="-1" resultid="7692" />
                    <RANKING order="17" place="-1" resultid="8386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6472" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9589" />
                    <RANKING order="2" place="2" resultid="7706" />
                    <RANKING order="3" place="3" resultid="6955" />
                    <RANKING order="4" place="4" resultid="9037" />
                    <RANKING order="5" place="5" resultid="11384" />
                    <RANKING order="6" place="6" resultid="8252" />
                    <RANKING order="7" place="7" resultid="7942" />
                    <RANKING order="8" place="8" resultid="9462" />
                    <RANKING order="9" place="9" resultid="7971" />
                    <RANKING order="10" place="10" resultid="7948" />
                    <RANKING order="11" place="11" resultid="9629" />
                    <RANKING order="12" place="12" resultid="9301" />
                    <RANKING order="13" place="13" resultid="7960" />
                    <RANKING order="14" place="14" resultid="11363" />
                    <RANKING order="15" place="15" resultid="7865" />
                    <RANKING order="16" place="16" resultid="7487" />
                    <RANKING order="17" place="17" resultid="8642" />
                    <RANKING order="18" place="18" resultid="8903" />
                    <RANKING order="19" place="19" resultid="9687" />
                    <RANKING order="20" place="20" resultid="7228" />
                    <RANKING order="21" place="-1" resultid="8815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6473" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7663" />
                    <RANKING order="2" place="2" resultid="8711" />
                    <RANKING order="3" place="3" resultid="8895" />
                    <RANKING order="4" place="4" resultid="7043" />
                    <RANKING order="5" place="5" resultid="9644" />
                    <RANKING order="6" place="6" resultid="8810" />
                    <RANKING order="7" place="7" resultid="7179" />
                    <RANKING order="8" place="7" resultid="7999" />
                    <RANKING order="9" place="9" resultid="7751" />
                    <RANKING order="10" place="10" resultid="8207" />
                    <RANKING order="11" place="11" resultid="9291" />
                    <RANKING order="12" place="12" resultid="9696" />
                    <RANKING order="13" place="13" resultid="7224" />
                    <RANKING order="14" place="14" resultid="8703" />
                    <RANKING order="15" place="15" resultid="8374" />
                    <RANKING order="16" place="16" resultid="9213" />
                    <RANKING order="17" place="17" resultid="8226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6474" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8066" />
                    <RANKING order="2" place="2" resultid="8436" />
                    <RANKING order="3" place="3" resultid="8962" />
                    <RANKING order="4" place="4" resultid="9526" />
                    <RANKING order="5" place="5" resultid="9105" />
                    <RANKING order="6" place="6" resultid="9164" />
                    <RANKING order="7" place="7" resultid="6823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6475" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6793" />
                    <RANKING order="2" place="2" resultid="8657" />
                    <RANKING order="3" place="3" resultid="7302" />
                    <RANKING order="4" place="4" resultid="8203" />
                    <RANKING order="5" place="5" resultid="9843" />
                    <RANKING order="6" place="6" resultid="7051" />
                    <RANKING order="7" place="7" resultid="8199" />
                    <RANKING order="8" place="8" resultid="8044" />
                    <RANKING order="9" place="9" resultid="8861" />
                    <RANKING order="10" place="-1" resultid="6873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6476" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7924" />
                    <RANKING order="2" place="2" resultid="9807" />
                    <RANKING order="3" place="3" resultid="8026" />
                    <RANKING order="4" place="4" resultid="9614" />
                    <RANKING order="5" place="5" resultid="7244" />
                    <RANKING order="6" place="-1" resultid="8573" />
                    <RANKING order="7" place="-1" resultid="9635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6477" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9326" />
                    <RANKING order="2" place="2" resultid="7316" />
                    <RANKING order="3" place="3" resultid="7427" />
                    <RANKING order="4" place="4" resultid="7155" />
                    <RANKING order="5" place="5" resultid="6840" />
                    <RANKING order="6" place="6" resultid="8145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6478" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7513" />
                    <RANKING order="2" place="2" resultid="7642" />
                    <RANKING order="3" place="3" resultid="6831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6479" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6480" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6481" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6482" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6483" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11529" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11530" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11531" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11532" daytime="16:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11533" daytime="16:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11534" daytime="16:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11535" daytime="16:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11536" daytime="16:12" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11537" daytime="16:14" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11538" daytime="16:14" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11539" daytime="16:16" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="11540" daytime="16:16" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="11541" daytime="16:18" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="11542" daytime="16:18" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6484" daytime="16:20" gender="F" number="25" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6485" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6486" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9452" />
                    <RANKING order="2" place="2" resultid="8195" />
                    <RANKING order="3" place="3" resultid="9583" />
                    <RANKING order="4" place="4" resultid="9577" />
                    <RANKING order="5" place="5" resultid="7499" />
                    <RANKING order="6" place="-1" resultid="9083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6487" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8310" />
                    <RANKING order="2" place="2" resultid="8295" />
                    <RANKING order="3" place="3" resultid="7759" />
                    <RANKING order="4" place="4" resultid="8530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6488" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7657" />
                    <RANKING order="2" place="2" resultid="9444" />
                    <RANKING order="3" place="3" resultid="8303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6489" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9198" />
                    <RANKING order="2" place="2" resultid="8164" />
                    <RANKING order="3" place="3" resultid="8089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6490" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9152" />
                    <RANKING order="2" place="2" resultid="9239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6491" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6492" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8013" />
                    <RANKING order="2" place="2" resultid="8801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6493" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9253" />
                    <RANKING order="2" place="2" resultid="9921" />
                    <RANKING order="3" place="3" resultid="8157" />
                    <RANKING order="4" place="-1" resultid="8097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6494" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9510" />
                    <RANKING order="2" place="2" resultid="6969" />
                    <RANKING order="3" place="3" resultid="7378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6495" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7539" />
                    <RANKING order="2" place="2" resultid="7372" />
                    <RANKING order="3" place="-1" resultid="7385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6496" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7391" />
                    <RANKING order="2" place="2" resultid="7163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6497" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6498" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6499" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6500" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11543" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11544" daytime="16:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11545" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11546" daytime="16:32" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6501" daytime="16:36" gender="M" number="26" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6502" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8953" />
                    <RANKING order="2" place="2" resultid="8469" />
                    <RANKING order="3" place="3" resultid="8477" />
                    <RANKING order="4" place="4" resultid="8542" />
                    <RANKING order="5" place="-1" resultid="7992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6503" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6977" />
                    <RANKING order="2" place="2" resultid="7849" />
                    <RANKING order="3" place="3" resultid="8821" />
                    <RANKING order="4" place="4" resultid="9181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6504" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6505" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9773" />
                    <RANKING order="2" place="2" resultid="8522" />
                    <RANKING order="3" place="3" resultid="8248" />
                    <RANKING order="4" place="4" resultid="7287" />
                    <RANKING order="5" place="-1" resultid="7480" />
                    <RANKING order="6" place="-1" resultid="8673" />
                    <RANKING order="7" place="-1" resultid="9693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6506" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9590" />
                    <RANKING order="2" place="2" resultid="7707" />
                    <RANKING order="3" place="3" resultid="7949" />
                    <RANKING order="4" place="4" resultid="7714" />
                    <RANKING order="5" place="5" resultid="7080" />
                    <RANKING order="6" place="6" resultid="7492" />
                    <RANKING order="7" place="7" resultid="8632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6507" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7664" />
                    <RANKING order="2" place="2" resultid="9112" />
                    <RANKING order="3" place="3" resultid="7059" />
                    <RANKING order="4" place="4" resultid="8909" />
                    <RANKING order="5" place="5" resultid="8773" />
                    <RANKING order="6" place="6" resultid="9160" />
                    <RANKING order="7" place="7" resultid="7326" />
                    <RANKING order="8" place="8" resultid="7457" />
                    <RANKING order="9" place="9" resultid="6938" />
                    <RANKING order="10" place="-1" resultid="9076" />
                    <RANKING order="11" place="-1" resultid="9381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6508" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6994" />
                    <RANKING order="2" place="2" resultid="8106" />
                    <RANKING order="3" place="3" resultid="8963" />
                    <RANKING order="4" place="4" resultid="7420" />
                    <RANKING order="5" place="5" resultid="9188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6509" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9016" />
                    <RANKING order="2" place="2" resultid="7303" />
                    <RANKING order="3" place="3" resultid="7052" />
                    <RANKING order="4" place="4" resultid="7120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6510" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9458" />
                    <RANKING order="2" place="2" resultid="7444" />
                    <RANKING order="3" place="3" resultid="7744" />
                    <RANKING order="4" place="4" resultid="9310" />
                    <RANKING order="5" place="5" resultid="9493" />
                    <RANKING order="6" place="-1" resultid="8982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6511" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9336" />
                    <RANKING order="2" place="2" resultid="7526" />
                    <RANKING order="3" place="3" resultid="9425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6512" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9185" />
                    <RANKING order="2" place="2" resultid="9503" />
                    <RANKING order="3" place="3" resultid="7026" />
                    <RANKING order="4" place="4" resultid="9388" />
                    <RANKING order="5" place="-1" resultid="7590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6513" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7533" />
                    <RANKING order="2" place="2" resultid="7406" />
                    <RANKING order="3" place="3" resultid="7399" />
                    <RANKING order="4" place="4" resultid="6895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6514" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6515" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6516" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6517" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11547" daytime="16:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11548" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11549" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11550" daytime="16:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11551" daytime="16:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11552" daytime="16:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11553" daytime="16:56" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6518" daytime="16:58" gender="F" number="27" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6519" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7138" />
                    <RANKING order="2" place="2" resultid="8614" />
                    <RANKING order="3" place="3" resultid="8495" />
                    <RANKING order="4" place="4" resultid="6866" />
                    <RANKING order="5" place="5" resultid="8187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6520" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7793" />
                    <RANKING order="2" place="2" resultid="8937" />
                    <RANKING order="3" place="3" resultid="8407" />
                    <RANKING order="4" place="4" resultid="7617" />
                    <RANKING order="5" place="5" resultid="9547" />
                    <RANKING order="6" place="6" resultid="8181" />
                    <RANKING order="7" place="-1" resultid="9935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6521" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9553" />
                    <RANKING order="2" place="2" resultid="8111" />
                    <RANKING order="3" place="3" resultid="7760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6522" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9445" />
                    <RANKING order="2" place="2" resultid="7345" />
                    <RANKING order="3" place="3" resultid="7771" />
                    <RANKING order="4" place="4" resultid="7171" />
                    <RANKING order="5" place="5" resultid="8665" />
                    <RANKING order="6" place="6" resultid="9476" />
                    <RANKING order="7" place="7" resultid="8288" />
                    <RANKING order="8" place="8" resultid="8563" />
                    <RANKING order="9" place="9" resultid="7678" />
                    <RANKING order="10" place="-1" resultid="9369" />
                    <RANKING order="11" place="-1" resultid="9570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6523" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7114" />
                    <RANKING order="2" place="2" resultid="9878" />
                    <RANKING order="3" place="3" resultid="8165" />
                    <RANKING order="4" place="4" resultid="9559" />
                    <RANKING order="5" place="5" resultid="8595" />
                    <RANKING order="6" place="6" resultid="9402" />
                    <RANKING order="7" place="-1" resultid="9262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6524" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8214" />
                    <RANKING order="2" place="2" resultid="8695" />
                    <RANKING order="3" place="3" resultid="9347" />
                    <RANKING order="4" place="4" resultid="9270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6525" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7553" />
                    <RANKING order="2" place="2" resultid="7724" />
                    <RANKING order="3" place="3" resultid="8334" />
                    <RANKING order="4" place="4" resultid="8328" />
                    <RANKING order="5" place="5" resultid="8552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6526" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7450" />
                    <RANKING order="2" place="2" resultid="8802" />
                    <RANKING order="3" place="3" resultid="9791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6527" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8053" />
                    <RANKING order="2" place="2" resultid="7309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6528" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6529" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9468" />
                    <RANKING order="2" place="2" resultid="7540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6530" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6531" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6532" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6533" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6534" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11554" daytime="16:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11555" daytime="17:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11556" daytime="17:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11557" daytime="17:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11558" daytime="17:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11559" daytime="17:24" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6535" daytime="17:28" gender="M" number="28" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6536" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8927" />
                    <RANKING order="2" place="2" resultid="9228" />
                    <RANKING order="3" place="3" resultid="8946" />
                    <RANKING order="4" place="4" resultid="9719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6537" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9778" />
                    <RANKING order="2" place="2" resultid="8841" />
                    <RANKING order="3" place="3" resultid="9726" />
                    <RANKING order="4" place="4" resultid="9124" />
                    <RANKING order="5" place="5" resultid="7600" />
                    <RANKING order="6" place="6" resultid="9749" />
                    <RANKING order="7" place="7" resultid="7626" />
                    <RANKING order="8" place="8" resultid="9609" />
                    <RANKING order="9" place="9" resultid="8400" />
                    <RANKING order="10" place="-1" resultid="11388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6538" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8367" />
                    <RANKING order="2" place="2" resultid="9024" />
                    <RANKING order="3" place="3" resultid="11350" />
                    <RANKING order="4" place="4" resultid="7838" />
                    <RANKING order="5" place="5" resultid="7075" />
                    <RANKING order="6" place="6" resultid="7259" />
                    <RANKING order="7" place="7" resultid="8690" />
                    <RANKING order="8" place="8" resultid="8583" />
                    <RANKING order="9" place="9" resultid="8451" />
                    <RANKING order="10" place="10" resultid="7361" />
                    <RANKING order="11" place="11" resultid="9742" />
                    <RANKING order="12" place="12" resultid="9136" />
                    <RANKING order="13" place="13" resultid="7239" />
                    <RANKING order="14" place="-1" resultid="7295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6539" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7693" />
                    <RANKING order="2" place="2" resultid="9118" />
                    <RANKING order="3" place="3" resultid="7433" />
                    <RANKING order="4" place="4" resultid="9086" />
                    <RANKING order="5" place="5" resultid="9515" />
                    <RANKING order="6" place="6" resultid="9622" />
                    <RANKING order="7" place="7" resultid="7481" />
                    <RANKING order="8" place="8" resultid="9146" />
                    <RANKING order="9" place="9" resultid="9682" />
                    <RANKING order="10" place="10" resultid="8380" />
                    <RANKING order="11" place="11" resultid="8221" />
                    <RANKING order="12" place="-1" resultid="6910" />
                    <RANKING order="13" place="-1" resultid="8387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6540" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7571" />
                    <RANKING order="2" place="2" resultid="6956" />
                    <RANKING order="3" place="3" resultid="7084" />
                    <RANKING order="4" place="4" resultid="8752" />
                    <RANKING order="5" place="5" resultid="7018" />
                    <RANKING order="6" place="6" resultid="7866" />
                    <RANKING order="7" place="7" resultid="8618" />
                    <RANKING order="8" place="8" resultid="7943" />
                    <RANKING order="9" place="9" resultid="8904" />
                    <RANKING order="10" place="10" resultid="9688" />
                    <RANKING order="11" place="11" resultid="9757" />
                    <RANKING order="12" place="12" resultid="8508" />
                    <RANKING order="13" place="13" resultid="8633" />
                    <RANKING order="14" place="-1" resultid="7201" />
                    <RANKING order="15" place="-1" resultid="7493" />
                    <RANKING order="16" place="-1" resultid="9071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6541" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7044" />
                    <RANKING order="2" place="2" resultid="9849" />
                    <RANKING order="3" place="3" resultid="7336" />
                    <RANKING order="4" place="4" resultid="8774" />
                    <RANKING order="5" place="5" resultid="7752" />
                    <RANKING order="6" place="6" resultid="9602" />
                    <RANKING order="7" place="7" resultid="8704" />
                    <RANKING order="8" place="8" resultid="7327" />
                    <RANKING order="9" place="9" resultid="8281" />
                    <RANKING order="10" place="10" resultid="9292" />
                    <RANKING order="11" place="11" resultid="7458" />
                    <RANKING order="12" place="12" resultid="6939" />
                    <RANKING order="13" place="13" resultid="9822" />
                    <RANKING order="14" place="14" resultid="8719" />
                    <RANKING order="15" place="15" resultid="8622" />
                    <RANKING order="16" place="-1" resultid="9077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6542" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8871" />
                    <RANKING order="2" place="2" resultid="9106" />
                    <RANKING order="3" place="3" resultid="7856" />
                    <RANKING order="4" place="4" resultid="8435" />
                    <RANKING order="5" place="5" resultid="8767" />
                    <RANKING order="6" place="6" resultid="7001" />
                    <RANKING order="7" place="7" resultid="8277" />
                    <RANKING order="8" place="8" resultid="8735" />
                    <RANKING order="9" place="9" resultid="7785" />
                    <RANKING order="10" place="-1" resultid="6989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6543" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6794" />
                    <RANKING order="2" place="2" resultid="8651" />
                    <RANKING order="3" place="3" resultid="9017" />
                    <RANKING order="4" place="4" resultid="9844" />
                    <RANKING order="5" place="5" resultid="6849" />
                    <RANKING order="6" place="6" resultid="8851" />
                    <RANKING order="7" place="7" resultid="7732" />
                    <RANKING order="8" place="8" resultid="9915" />
                    <RANKING order="9" place="-1" resultid="7185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6544" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7036" />
                    <RANKING order="2" place="2" resultid="9375" />
                    <RANKING order="3" place="3" resultid="7745" />
                    <RANKING order="4" place="4" resultid="9615" />
                    <RANKING order="5" place="5" resultid="9808" />
                    <RANKING order="6" place="6" resultid="8260" />
                    <RANKING order="7" place="-1" resultid="7925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6545" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7527" />
                    <RANKING order="2" place="2" resultid="9426" />
                    <RANKING order="3" place="3" resultid="8915" />
                    <RANKING order="4" place="4" resultid="6841" />
                    <RANKING order="5" place="-1" resultid="9327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6546" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7643" />
                    <RANKING order="2" place="2" resultid="9284" />
                    <RANKING order="3" place="3" resultid="9053" />
                    <RANKING order="4" place="-1" resultid="7415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6547" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6548" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7519" />
                    <RANKING order="2" place="2" resultid="8074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6549" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6550" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6551" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11560" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11561" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11562" daytime="17:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11563" daytime="17:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11564" daytime="17:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11565" daytime="17:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11566" daytime="18:02" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11567" daytime="18:06" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11568" daytime="18:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11569" daytime="18:12" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11570" daytime="18:16" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="11571" daytime="18:18" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6552" daytime="18:22" gender="F" number="29" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6553" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6867" />
                    <RANKING order="2" place="2" resultid="8488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6554" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9045" />
                    <RANKING order="2" place="2" resultid="7830" />
                    <RANKING order="3" place="3" resultid="9936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6555" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7581" />
                    <RANKING order="2" place="2" resultid="8359" />
                    <RANKING order="3" place="3" resultid="9929" />
                    <RANKING order="4" place="4" resultid="8744" />
                    <RANKING order="5" place="-1" resultid="9652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6556" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7174" />
                    <RANKING order="2" place="2" resultid="8289" />
                    <RANKING order="3" place="3" resultid="8564" />
                    <RANKING order="4" place="4" resultid="8129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6557" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8880" />
                    <RANKING order="2" place="-1" resultid="7205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6558" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8789" />
                    <RANKING order="2" place="2" resultid="8696" />
                    <RANKING order="3" place="3" resultid="9348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6559" agemax="54" agemin="50" name="Kat. F" />
                <AGEGROUP agegroupid="6560" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="6561" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9922" />
                    <RANKING order="2" place="2" resultid="8098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6562" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="6563" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="6564" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6565" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6566" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6567" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6568" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11572" daytime="18:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11573" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11574" daytime="18:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6569" daytime="18:48" gender="M" number="30" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6570" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9229" />
                    <RANKING order="2" place="2" resultid="8478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6571" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6572" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9356" />
                    <RANKING order="2" place="2" resultid="9764" />
                    <RANKING order="3" place="3" resultid="7842" />
                    <RANKING order="4" place="4" resultid="8604" />
                    <RANKING order="5" place="5" resultid="9706" />
                    <RANKING order="6" place="6" resultid="6929" />
                    <RANKING order="7" place="-1" resultid="7260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6573" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="6574" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7572" />
                    <RANKING order="2" place="2" resultid="8753" />
                    <RANKING order="3" place="3" resultid="7715" />
                    <RANKING order="4" place="4" resultid="8643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6575" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8712" />
                    <RANKING order="2" place="2" resultid="9487" />
                    <RANKING order="3" place="3" resultid="7060" />
                    <RANKING order="4" place="4" resultid="8910" />
                    <RANKING order="5" place="5" resultid="9382" />
                    <RANKING order="6" place="-1" resultid="9659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6576" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6995" />
                    <RANKING order="2" place="2" resultid="9527" />
                    <RANKING order="3" place="3" resultid="8447" />
                    <RANKING order="4" place="4" resultid="8831" />
                    <RANKING order="5" place="5" resultid="6824" />
                    <RANKING order="6" place="-1" resultid="7216" />
                    <RANKING order="7" place="-1" resultid="8872" />
                    <RANKING order="8" place="-1" resultid="9839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6577" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8652" />
                    <RANKING order="2" place="2" resultid="7689" />
                    <RANKING order="3" place="3" resultid="8678" />
                    <RANKING order="4" place="4" resultid="8862" />
                    <RANKING order="5" place="-1" resultid="6850" />
                    <RANKING order="6" place="-1" resultid="7213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6578" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7037" />
                    <RANKING order="2" place="2" resultid="6858" />
                    <RANKING order="3" place="3" resultid="8574" />
                    <RANKING order="4" place="-1" resultid="9636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6579" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6882" />
                    <RANKING order="2" place="2" resultid="7156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6580" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9665" />
                    <RANKING order="2" place="2" resultid="7027" />
                    <RANKING order="3" place="3" resultid="6832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6581" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6582" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6583" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6584" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6585" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11575" daytime="18:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11576" daytime="19:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11577" daytime="19:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11578" daytime="19:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11579" daytime="19:30" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6586" daytime="19:36" gender="F" number="31" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6603" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6604" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6605" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8360" />
                    <RANKING order="2" place="2" resultid="9671" />
                    <RANKING order="3" place="3" resultid="8230" />
                    <RANKING order="4" place="4" resultid="9859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6606" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6607" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9830" />
                    <RANKING order="2" place="2" resultid="9861" />
                    <RANKING order="3" place="3" resultid="9411" />
                    <RANKING order="4" place="4" resultid="8238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6608" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="6609" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11580" daytime="19:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11581" daytime="19:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6610" daytime="19:44" gender="M" number="32" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6611" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6612" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="6613" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11371" />
                    <RANKING order="2" place="2" resultid="9094" />
                    <RANKING order="3" place="3" resultid="8779" />
                    <RANKING order="4" place="4" resultid="9863" />
                    <RANKING order="5" place="5" resultid="9857" />
                    <RANKING order="6" place="6" resultid="11372" />
                    <RANKING order="7" place="-1" resultid="8845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6614" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9907" />
                    <RANKING order="2" place="2" resultid="9672" />
                    <RANKING order="3" place="3" resultid="9128" />
                    <RANKING order="4" place="4" resultid="8918" />
                    <RANKING order="5" place="5" resultid="9835" />
                    <RANKING order="6" place="6" resultid="8780" />
                    <RANKING order="7" place="7" resultid="9414" />
                    <RANKING order="8" place="8" resultid="8240" />
                    <RANKING order="9" place="9" resultid="8006" />
                    <RANKING order="10" place="-1" resultid="7245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6615" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9837" />
                    <RANKING order="2" place="2" resultid="9908" />
                    <RANKING order="3" place="3" resultid="8242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6616" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9829" />
                    <RANKING order="2" place="-1" resultid="9413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6617" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9912" />
                    <RANKING order="2" place="2" resultid="9412" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11582" daytime="19:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11583" daytime="19:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11584" daytime="19:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-12-18" daytime="08:30" endtime="12:31" number="4">
          <EVENTS>
            <EVENT eventid="6618" daytime="08:30" gender="F" number="33" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6620" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7139" />
                    <RANKING order="2" place="2" resultid="7507" />
                    <RANKING order="3" place="3" resultid="8489" />
                    <RANKING order="4" place="-1" resultid="8615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6621" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8938" />
                    <RANKING order="2" place="2" resultid="7609" />
                    <RANKING order="3" place="3" resultid="7831" />
                    <RANKING order="4" place="4" resultid="7618" />
                    <RANKING order="5" place="-1" resultid="7196" />
                    <RANKING order="6" place="-1" resultid="8408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6622" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8745" />
                    <RANKING order="2" place="2" resultid="9653" />
                    <RANKING order="3" place="3" resultid="8296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6623" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8304" />
                    <RANKING order="2" place="2" resultid="8666" />
                    <RANKING order="3" place="3" resultid="7173" />
                    <RANKING order="4" place="4" resultid="8565" />
                    <RANKING order="5" place="5" resultid="7679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6624" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9199" />
                    <RANKING order="2" place="2" resultid="7008" />
                    <RANKING order="3" place="3" resultid="7095" />
                    <RANKING order="4" place="4" resultid="8881" />
                    <RANKING order="5" place="5" resultid="9560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6625" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8790" />
                    <RANKING order="2" place="2" resultid="8998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6626" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9278" />
                    <RANKING order="2" place="2" resultid="8329" />
                    <RANKING order="3" place="3" resultid="8060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6627" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6628" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9254" />
                    <RANKING order="2" place="2" resultid="8054" />
                    <RANKING order="3" place="3" resultid="8099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6629" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6630" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="6631" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="6632" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6633" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6634" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6635" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11585" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11586" daytime="08:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11587" daytime="08:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11588" daytime="08:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6636" daytime="08:40" gender="M" number="34" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6637" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8928" />
                    <RANKING order="2" place="2" resultid="8947" />
                    <RANKING order="3" place="3" resultid="7191" />
                    <RANKING order="4" place="4" resultid="8954" />
                    <RANKING order="5" place="5" resultid="9720" />
                    <RANKING order="6" place="6" resultid="8479" />
                    <RANKING order="7" place="-1" resultid="7993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6638" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9221" />
                    <RANKING order="2" place="2" resultid="9030" />
                    <RANKING order="3" place="3" resultid="9779" />
                    <RANKING order="4" place="4" resultid="8827" />
                    <RANKING order="5" place="5" resultid="7601" />
                    <RANKING order="6" place="6" resultid="8430" />
                    <RANKING order="7" place="7" resultid="7649" />
                    <RANKING order="8" place="-1" resultid="7850" />
                    <RANKING order="9" place="-1" resultid="9750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6639" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9940" />
                    <RANKING order="2" place="2" resultid="8368" />
                    <RANKING order="3" place="3" resultid="9025" />
                    <RANKING order="4" place="4" resultid="8605" />
                    <RANKING order="5" place="5" resultid="9765" />
                    <RANKING order="6" place="6" resultid="11351" />
                    <RANKING order="7" place="7" resultid="7076" />
                    <RANKING order="8" place="8" resultid="9707" />
                    <RANKING order="9" place="9" resultid="8394" />
                    <RANKING order="10" place="10" resultid="9743" />
                    <RANKING order="11" place="11" resultid="6930" />
                    <RANKING order="12" place="-1" resultid="7261" />
                    <RANKING order="13" place="-1" resultid="9784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6640" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7694" />
                    <RANKING order="2" place="2" resultid="9119" />
                    <RANKING order="3" place="3" resultid="9087" />
                    <RANKING order="4" place="4" resultid="9147" />
                    <RANKING order="5" place="5" resultid="8762" />
                    <RANKING order="6" place="6" resultid="7288" />
                    <RANKING order="7" place="-1" resultid="6911" />
                    <RANKING order="8" place="-1" resultid="9516" />
                    <RANKING order="9" place="-1" resultid="9623" />
                    <RANKING order="10" place="-1" resultid="9802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6641" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7708" />
                    <RANKING order="2" place="2" resultid="6957" />
                    <RANKING order="3" place="3" resultid="7573" />
                    <RANKING order="4" place="4" resultid="8253" />
                    <RANKING order="5" place="5" resultid="11385" />
                    <RANKING order="6" place="6" resultid="7944" />
                    <RANKING order="7" place="7" resultid="7867" />
                    <RANKING order="8" place="8" resultid="7085" />
                    <RANKING order="9" place="-1" resultid="8619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6642" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7665" />
                    <RANKING order="2" place="2" resultid="8713" />
                    <RANKING order="3" place="3" resultid="7045" />
                    <RANKING order="4" place="4" resultid="8896" />
                    <RANKING order="5" place="5" resultid="7737" />
                    <RANKING order="6" place="6" resultid="9488" />
                    <RANKING order="7" place="7" resultid="7180" />
                    <RANKING order="8" place="8" resultid="7753" />
                    <RANKING order="9" place="9" resultid="9214" />
                    <RANKING order="10" place="-1" resultid="6940" />
                    <RANKING order="11" place="-1" resultid="7337" />
                    <RANKING order="12" place="-1" resultid="9293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6643" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8067" />
                    <RANKING order="2" place="2" resultid="9528" />
                    <RANKING order="3" place="3" resultid="8964" />
                    <RANKING order="4" place="4" resultid="8438" />
                    <RANKING order="5" place="5" resultid="8107" />
                    <RANKING order="6" place="6" resultid="9165" />
                    <RANKING order="7" place="7" resultid="6825" />
                    <RANKING order="8" place="-1" resultid="6990" />
                    <RANKING order="9" place="-1" resultid="8832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6644" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6795" />
                    <RANKING order="2" place="2" resultid="7304" />
                    <RANKING order="3" place="3" resultid="8658" />
                    <RANKING order="4" place="4" resultid="8679" />
                    <RANKING order="5" place="5" resultid="8863" />
                    <RANKING order="6" place="6" resultid="6851" />
                    <RANKING order="7" place="-1" resultid="6874" />
                    <RANKING order="8" place="-1" resultid="7053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6645" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7445" />
                    <RANKING order="2" place="2" resultid="8575" />
                    <RANKING order="3" place="3" resultid="8027" />
                    <RANKING order="4" place="-1" resultid="6859" />
                    <RANKING order="5" place="-1" resultid="9637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6646" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9328" />
                    <RANKING order="2" place="2" resultid="6883" />
                    <RANKING order="3" place="3" resultid="7157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6647" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6833" />
                    <RANKING order="2" place="2" resultid="9054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6648" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6649" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6650" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6651" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6652" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11589" daytime="08:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11590" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11591" daytime="08:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11592" daytime="08:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11593" daytime="08:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11594" daytime="08:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11595" daytime="08:56" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11596" daytime="08:58" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11597" daytime="09:00" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6653" daytime="09:02" gender="F" number="35" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6654" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8496" />
                    <RANKING order="2" place="2" resultid="6868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6655" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9578" />
                    <RANKING order="2" place="-1" resultid="9453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6656" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6657" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7658" />
                    <RANKING order="2" place="2" resultid="9446" />
                    <RANKING order="3" place="3" resultid="8305" />
                    <RANKING order="4" place="4" resultid="7346" />
                    <RANKING order="5" place="-1" resultid="7772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6658" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8166" />
                    <RANKING order="2" place="2" resultid="8090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6659" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8791" />
                    <RANKING order="2" place="2" resultid="9153" />
                    <RANKING order="3" place="3" resultid="9240" />
                    <RANKING order="4" place="4" resultid="9349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6660" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6661" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8803" />
                    <RANKING order="2" place="-1" resultid="8014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6662" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6663" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6970" />
                    <RANKING order="2" place="2" resultid="7379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6664" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7541" />
                    <RANKING order="2" place="2" resultid="7373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6665" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7392" />
                    <RANKING order="2" place="2" resultid="7165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6666" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6667" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6668" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6669" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11598" daytime="09:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11599" daytime="09:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11600" daytime="09:16" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6670" daytime="09:20" gender="M" number="36" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6671" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8955" />
                    <RANKING order="2" place="2" resultid="9230" />
                    <RANKING order="3" place="3" resultid="8480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6672" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6978" />
                    <RANKING order="2" place="2" resultid="9182" />
                    <RANKING order="3" place="3" resultid="8822" />
                    <RANKING order="4" place="-1" resultid="7129" />
                    <RANKING order="5" place="-1" resultid="8684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6673" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6674" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8523" />
                    <RANKING order="2" place="2" resultid="8249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6675" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7709" />
                    <RANKING order="2" place="2" resultid="7950" />
                    <RANKING order="3" place="3" resultid="7716" />
                    <RANKING order="4" place="4" resultid="8754" />
                    <RANKING order="5" place="5" resultid="7081" />
                    <RANKING order="6" place="6" resultid="8634" />
                    <RANKING order="7" place="-1" resultid="7494" />
                    <RANKING order="8" place="-1" resultid="8644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6676" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7738" />
                    <RANKING order="2" place="2" resultid="7061" />
                    <RANKING order="3" place="3" resultid="9113" />
                    <RANKING order="4" place="4" resultid="8775" />
                    <RANKING order="5" place="5" resultid="8911" />
                    <RANKING order="6" place="6" resultid="7328" />
                    <RANKING order="7" place="7" resultid="7459" />
                    <RANKING order="8" place="-1" resultid="8020" />
                    <RANKING order="9" place="-1" resultid="8705" />
                    <RANKING order="10" place="-1" resultid="9078" />
                    <RANKING order="11" place="-1" resultid="9697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6677" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6996" />
                    <RANKING order="2" place="2" resultid="8108" />
                    <RANKING order="3" place="3" resultid="8965" />
                    <RANKING order="4" place="4" resultid="9189" />
                    <RANKING order="5" place="-1" resultid="8873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6678" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9018" />
                    <RANKING order="2" place="2" resultid="7054" />
                    <RANKING order="3" place="3" resultid="7121" />
                    <RANKING order="4" place="4" resultid="8045" />
                    <RANKING order="5" place="5" resultid="8852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6679" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9459" />
                    <RANKING order="2" place="2" resultid="7038" />
                    <RANKING order="3" place="3" resultid="7746" />
                    <RANKING order="4" place="4" resultid="9494" />
                    <RANKING order="5" place="-1" resultid="7219" />
                    <RANKING order="6" place="-1" resultid="8983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6680" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7158" />
                    <RANKING order="2" place="2" resultid="7528" />
                    <RANKING order="3" place="3" resultid="9427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6681" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9362" />
                    <RANKING order="2" place="2" resultid="9186" />
                    <RANKING order="3" place="3" resultid="9504" />
                    <RANKING order="4" place="4" resultid="7028" />
                    <RANKING order="5" place="-1" resultid="7591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6682" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7534" />
                    <RANKING order="2" place="2" resultid="7407" />
                    <RANKING order="3" place="3" resultid="6896" />
                    <RANKING order="4" place="-1" resultid="7400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6683" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6684" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6685" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6686" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11601" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11602" daytime="09:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11603" daytime="09:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11604" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11605" daytime="09:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11606" daytime="09:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6687" daytime="09:52" gender="F" number="37" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6688" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7508" />
                    <RANKING order="2" place="2" resultid="8490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6689" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7671" />
                    <RANKING order="2" place="2" resultid="7469" />
                    <RANKING order="3" place="3" resultid="7794" />
                    <RANKING order="4" place="4" resultid="7610" />
                    <RANKING order="5" place="-1" resultid="9046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6690" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7965" />
                    <RANKING order="2" place="2" resultid="7582" />
                    <RANKING order="3" place="3" resultid="8531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6691" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9477" />
                    <RANKING order="2" place="2" resultid="7659" />
                    <RANKING order="3" place="3" resultid="7347" />
                    <RANKING order="4" place="4" resultid="9370" />
                    <RANKING order="5" place="5" resultid="7905" />
                    <RANKING order="6" place="-1" resultid="8082" />
                    <RANKING order="7" place="-1" resultid="9571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6692" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7009" />
                    <RANKING order="2" place="2" resultid="7885" />
                    <RANKING order="3" place="3" resultid="8091" />
                    <RANKING order="4" place="4" resultid="9206" />
                    <RANKING order="5" place="5" resultid="9483" />
                    <RANKING order="6" place="6" resultid="9263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6693" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8421" />
                    <RANKING order="2" place="2" resultid="9154" />
                    <RANKING order="3" place="3" resultid="9241" />
                    <RANKING order="4" place="4" resultid="9271" />
                    <RANKING order="5" place="5" resultid="9005" />
                    <RANKING order="6" place="6" resultid="8999" />
                    <RANKING order="7" place="7" resultid="9247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6694" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7725" />
                    <RANKING order="2" place="2" resultid="8335" />
                    <RANKING order="3" place="3" resultid="7354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6695" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8015" />
                    <RANKING order="2" place="2" resultid="8142" />
                    <RANKING order="3" place="3" resultid="7766" />
                    <RANKING order="4" place="-1" resultid="9792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6696" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8158" />
                    <RANKING order="2" place="2" resultid="9255" />
                    <RANKING order="3" place="3" resultid="8323" />
                    <RANKING order="4" place="4" resultid="8150" />
                    <RANKING order="5" place="5" resultid="7310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6697" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9012" />
                    <RANKING order="2" place="2" resultid="9512" />
                    <RANKING order="3" place="3" resultid="7106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6698" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7936" />
                    <RANKING order="2" place="2" resultid="7548" />
                    <RANKING order="3" place="3" resultid="6921" />
                    <RANKING order="4" place="4" resultid="9469" />
                    <RANKING order="5" place="5" resultid="7386" />
                    <RANKING order="6" place="6" resultid="7374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6699" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7393" />
                    <RANKING order="2" place="-1" resultid="7109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6700" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6701" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6702" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6703" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11607" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11608" daytime="09:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11609" daytime="09:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11610" daytime="09:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11611" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11612" daytime="10:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6704" daytime="10:02" gender="M" number="38" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6705" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9820" />
                    <RANKING order="2" place="2" resultid="8458" />
                    <RANKING order="3" place="3" resultid="8470" />
                    <RANKING order="4" place="4" resultid="8543" />
                    <RANKING order="5" place="-1" resultid="7994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6706" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8989" />
                    <RANKING order="2" place="2" resultid="7461" />
                    <RANKING order="3" place="3" resultid="8171" />
                    <RANKING order="4" place="4" resultid="9173" />
                    <RANKING order="5" place="5" resultid="7252" />
                    <RANKING order="6" place="6" resultid="8626" />
                    <RANKING order="7" place="7" resultid="8431" />
                    <RANKING order="8" place="8" resultid="7148" />
                    <RANKING order="9" place="9" resultid="7627" />
                    <RANKING order="10" place="-1" resultid="7851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6707" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9176" />
                    <RANKING order="2" place="2" resultid="8857" />
                    <RANKING order="3" place="3" resultid="9357" />
                    <RANKING order="4" place="4" resultid="9766" />
                    <RANKING order="5" place="5" resultid="8606" />
                    <RANKING order="6" place="6" resultid="9138" />
                    <RANKING order="7" place="-1" resultid="7240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6708" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8443" />
                    <RANKING order="2" place="2" resultid="9596" />
                    <RANKING order="3" place="3" resultid="7637" />
                    <RANKING order="4" place="4" resultid="9127" />
                    <RANKING order="5" place="5" resultid="7980" />
                    <RANKING order="6" place="6" resultid="6890" />
                    <RANKING order="7" place="7" resultid="7289" />
                    <RANKING order="8" place="8" resultid="8763" />
                    <RANKING order="9" place="9" resultid="11378" />
                    <RANKING order="10" place="-1" resultid="6912" />
                    <RANKING order="11" place="-1" resultid="9624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6709" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9038" />
                    <RANKING order="2" place="2" resultid="9591" />
                    <RANKING order="3" place="3" resultid="9302" />
                    <RANKING order="4" place="4" resultid="8816" />
                    <RANKING order="5" place="5" resultid="8725" />
                    <RANKING order="6" place="6" resultid="7069" />
                    <RANKING order="7" place="7" resultid="9758" />
                    <RANKING order="8" place="8" resultid="9341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6710" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9645" />
                    <RANKING order="2" place="2" resultid="7338" />
                    <RANKING order="3" place="3" resultid="8811" />
                    <RANKING order="4" place="4" resultid="8897" />
                    <RANKING order="5" place="5" resultid="8267" />
                    <RANKING order="6" place="6" resultid="7280" />
                    <RANKING order="7" place="7" resultid="8282" />
                    <RANKING order="8" place="8" resultid="8208" />
                    <RANKING order="9" place="9" resultid="8021" />
                    <RANKING order="10" place="10" resultid="9383" />
                    <RANKING order="11" place="11" resultid="9161" />
                    <RANKING order="12" place="12" resultid="9215" />
                    <RANKING order="13" place="13" resultid="9317" />
                    <RANKING order="14" place="-1" resultid="7062" />
                    <RANKING order="15" place="-1" resultid="8000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6711" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6904" />
                    <RANKING order="2" place="2" resultid="8068" />
                    <RANKING order="3" place="3" resultid="7857" />
                    <RANKING order="4" place="4" resultid="7002" />
                    <RANKING order="5" place="5" resultid="7421" />
                    <RANKING order="6" place="6" resultid="7786" />
                    <RANKING order="7" place="7" resultid="8889" />
                    <RANKING order="8" place="8" resultid="8736" />
                    <RANKING order="9" place="9" resultid="9166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6712" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7686" />
                    <RANKING order="2" place="2" resultid="6796" />
                    <RANKING order="3" place="3" resultid="7305" />
                    <RANKING order="4" place="4" resultid="8115" />
                    <RANKING order="5" place="5" resultid="8046" />
                    <RANKING order="6" place="6" resultid="8200" />
                    <RANKING order="7" place="7" resultid="7733" />
                    <RANKING order="8" place="8" resultid="8864" />
                    <RANKING order="9" place="-1" resultid="7872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6713" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9871" />
                    <RANKING order="2" place="2" resultid="9060" />
                    <RANKING order="3" place="3" resultid="7446" />
                    <RANKING order="4" place="4" resultid="7275" />
                    <RANKING order="5" place="5" resultid="9393" />
                    <RANKING order="6" place="6" resultid="8977" />
                    <RANKING order="7" place="7" resultid="9311" />
                    <RANKING order="8" place="8" resultid="8028" />
                    <RANKING order="9" place="9" resultid="8972" />
                    <RANKING order="10" place="10" resultid="8261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6714" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7317" />
                    <RANKING order="2" place="2" resultid="7428" />
                    <RANKING order="3" place="3" resultid="6884" />
                    <RANKING order="4" place="-1" resultid="7910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6715" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9666" />
                    <RANKING order="2" place="2" resultid="9363" />
                    <RANKING order="3" place="3" resultid="7514" />
                    <RANKING order="4" place="4" resultid="7416" />
                    <RANKING order="5" place="5" resultid="9389" />
                    <RANKING order="6" place="6" resultid="6834" />
                    <RANKING order="7" place="-1" resultid="7592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6716" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7408" />
                    <RANKING order="2" place="2" resultid="6897" />
                    <RANKING order="3" place="3" resultid="7401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6717" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7919" />
                    <RANKING order="2" place="2" resultid="8075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6718" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6719" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6720" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11613" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11614" daytime="10:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11615" daytime="10:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11616" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11617" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11618" daytime="10:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11619" daytime="10:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11620" daytime="10:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11621" daytime="10:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11622" daytime="10:16" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="11623" daytime="10:18" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6721" daytime="10:20" gender="F" number="39" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6722" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7140" />
                    <RANKING order="2" place="2" resultid="8497" />
                    <RANKING order="3" place="3" resultid="6869" />
                    <RANKING order="4" place="4" resultid="8188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6723" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7795" />
                    <RANKING order="2" place="2" resultid="8939" />
                    <RANKING order="3" place="3" resultid="7832" />
                    <RANKING order="4" place="4" resultid="7619" />
                    <RANKING order="5" place="5" resultid="8409" />
                    <RANKING order="6" place="6" resultid="9937" />
                    <RANKING order="7" place="7" resultid="8182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6724" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7583" />
                    <RANKING order="2" place="2" resultid="9554" />
                    <RANKING order="3" place="3" resultid="9930" />
                    <RANKING order="4" place="4" resultid="8746" />
                    <RANKING order="5" place="5" resultid="8112" />
                    <RANKING order="6" place="6" resultid="7761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6725" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9447" />
                    <RANKING order="2" place="2" resultid="7172" />
                    <RANKING order="3" place="3" resultid="7773" />
                    <RANKING order="4" place="4" resultid="8667" />
                    <RANKING order="5" place="5" resultid="9371" />
                    <RANKING order="6" place="6" resultid="8290" />
                    <RANKING order="7" place="7" resultid="7680" />
                    <RANKING order="8" place="8" resultid="8130" />
                    <RANKING order="9" place="-1" resultid="8566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6726" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9879" />
                    <RANKING order="2" place="2" resultid="7096" />
                    <RANKING order="3" place="3" resultid="9561" />
                    <RANKING order="4" place="4" resultid="8882" />
                    <RANKING order="5" place="5" resultid="8596" />
                    <RANKING order="6" place="6" resultid="9403" />
                    <RANKING order="7" place="7" resultid="9264" />
                    <RANKING order="8" place="-1" resultid="8167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6727" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9350" />
                    <RANKING order="2" place="-1" resultid="8215" />
                    <RANKING order="3" place="-1" resultid="8838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6728" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7554" />
                    <RANKING order="2" place="2" resultid="7726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6729" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7451" />
                    <RANKING order="2" place="2" resultid="9793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6730" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8055" />
                    <RANKING order="2" place="2" resultid="9924" />
                    <RANKING order="3" place="3" resultid="8159" />
                    <RANKING order="4" place="4" resultid="8100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6731" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6732" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9566" />
                    <RANKING order="2" place="2" resultid="7542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6733" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6734" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="6735" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6736" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6737" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11624" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11625" daytime="10:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11626" daytime="10:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11627" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11628" daytime="10:56" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6738" daytime="11:04" gender="M" number="40" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6739" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9231" />
                    <RANKING order="2" place="2" resultid="8929" />
                    <RANKING order="3" place="-1" resultid="8459" />
                    <RANKING order="4" place="-1" resultid="8544" />
                    <RANKING order="5" place="-1" resultid="8948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6740" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7700" />
                    <RANKING order="2" place="2" resultid="8842" />
                    <RANKING order="3" place="3" resultid="9125" />
                    <RANKING order="4" place="4" resultid="7602" />
                    <RANKING order="5" place="5" resultid="9751" />
                    <RANKING order="6" place="6" resultid="7628" />
                    <RANKING order="7" place="7" resultid="8401" />
                    <RANKING order="8" place="-1" resultid="8685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6741" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9941" />
                    <RANKING order="2" place="2" resultid="8369" />
                    <RANKING order="3" place="3" resultid="11352" />
                    <RANKING order="4" place="4" resultid="9708" />
                    <RANKING order="5" place="5" resultid="8584" />
                    <RANKING order="6" place="6" resultid="9744" />
                    <RANKING order="7" place="7" resultid="6931" />
                    <RANKING order="8" place="-1" resultid="7241" />
                    <RANKING order="9" place="-1" resultid="7262" />
                    <RANKING order="10" place="-1" resultid="8691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6742" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7695" />
                    <RANKING order="2" place="2" resultid="7434" />
                    <RANKING order="3" place="3" resultid="9120" />
                    <RANKING order="4" place="4" resultid="9088" />
                    <RANKING order="5" place="5" resultid="7482" />
                    <RANKING order="6" place="6" resultid="8381" />
                    <RANKING order="7" place="7" resultid="8222" />
                    <RANKING order="8" place="-1" resultid="8388" />
                    <RANKING order="9" place="-1" resultid="9517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6743" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7574" />
                    <RANKING order="2" place="2" resultid="8755" />
                    <RANKING order="3" place="3" resultid="6958" />
                    <RANKING order="4" place="4" resultid="7019" />
                    <RANKING order="5" place="5" resultid="7868" />
                    <RANKING order="6" place="6" resultid="9072" />
                    <RANKING order="7" place="7" resultid="8905" />
                    <RANKING order="8" place="8" resultid="8635" />
                    <RANKING order="9" place="-1" resultid="7495" />
                    <RANKING order="10" place="-1" resultid="7717" />
                    <RANKING order="11" place="-1" resultid="7972" />
                    <RANKING order="12" place="-1" resultid="8645" />
                    <RANKING order="13" place="-1" resultid="9303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6744" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8714" />
                    <RANKING order="2" place="2" resultid="7046" />
                    <RANKING order="3" place="3" resultid="9850" />
                    <RANKING order="4" place="4" resultid="8776" />
                    <RANKING order="5" place="5" resultid="9646" />
                    <RANKING order="6" place="6" resultid="9603" />
                    <RANKING order="7" place="7" resultid="8706" />
                    <RANKING order="8" place="8" resultid="7329" />
                    <RANKING order="9" place="9" resultid="9294" />
                    <RANKING order="10" place="10" resultid="9384" />
                    <RANKING order="11" place="11" resultid="6941" />
                    <RANKING order="12" place="12" resultid="8720" />
                    <RANKING order="13" place="-1" resultid="7225" />
                    <RANKING order="14" place="-1" resultid="7754" />
                    <RANKING order="15" place="-1" resultid="9079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6745" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9107" />
                    <RANKING order="2" place="2" resultid="8874" />
                    <RANKING order="3" place="3" resultid="7858" />
                    <RANKING order="4" place="4" resultid="9529" />
                    <RANKING order="5" place="5" resultid="8768" />
                    <RANKING order="6" place="6" resultid="8890" />
                    <RANKING order="7" place="7" resultid="8833" />
                    <RANKING order="8" place="8" resultid="8737" />
                    <RANKING order="9" place="9" resultid="7787" />
                    <RANKING order="10" place="-1" resultid="9190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6746" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8653" />
                    <RANKING order="2" place="2" resultid="9019" />
                    <RANKING order="3" place="3" resultid="7690" />
                    <RANKING order="4" place="4" resultid="9845" />
                    <RANKING order="5" place="5" resultid="6852" />
                    <RANKING order="6" place="-1" resultid="7186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6747" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7039" />
                    <RANKING order="2" place="2" resultid="9376" />
                    <RANKING order="3" place="3" resultid="7747" />
                    <RANKING order="4" place="4" resultid="6860" />
                    <RANKING order="5" place="5" resultid="8262" />
                    <RANKING order="6" place="-1" resultid="7220" />
                    <RANKING order="7" place="-1" resultid="8576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6748" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7529" />
                    <RANKING order="2" place="2" resultid="9428" />
                    <RANKING order="3" place="3" resultid="8916" />
                    <RANKING order="4" place="4" resultid="6842" />
                    <RANKING order="5" place="-1" resultid="9329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6749" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7644" />
                    <RANKING order="2" place="2" resultid="9285" />
                    <RANKING order="3" place="3" resultid="9055" />
                    <RANKING order="4" place="4" resultid="7417" />
                    <RANKING order="5" place="5" resultid="7029" />
                    <RANKING order="6" place="-1" resultid="9505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6750" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6751" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7520" />
                    <RANKING order="2" place="2" resultid="8076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6752" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="6753" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="6754" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11629" daytime="11:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11630" daytime="11:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11631" daytime="11:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11632" daytime="11:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11633" daytime="11:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11634" daytime="11:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="11635" daytime="12:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="11636" daytime="12:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="11637" daytime="12:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="11638" daytime="12:20" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6755" daytime="12:26" gender="F" number="41" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6772" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6773" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6774" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9897" />
                    <RANKING order="2" place="2" resultid="9673" />
                    <RANKING order="3" place="3" resultid="8229" />
                    <RANKING order="4" place="-1" resultid="9860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6775" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6776" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9415" />
                    <RANKING order="2" place="2" resultid="8239" />
                    <RANKING order="3" place="-1" resultid="9862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6777" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="6778" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11639" daytime="12:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6779" daytime="12:30" gender="M" number="42" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6780" agemax="-1" agemin="-1" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6781" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="6782" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11375" />
                    <RANKING order="2" place="2" resultid="9097" />
                    <RANKING order="3" place="3" resultid="9895" />
                    <RANKING order="4" place="4" resultid="8846" />
                    <RANKING order="5" place="5" resultid="9129" />
                    <RANKING order="6" place="-1" resultid="11376" />
                    <RANKING order="7" place="-1" resultid="9858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6783" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8919" />
                    <RANKING order="2" place="2" resultid="8782" />
                    <RANKING order="3" place="3" resultid="8241" />
                    <RANKING order="4" place="-1" resultid="9418" />
                    <RANKING order="5" place="-1" resultid="9836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6784" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9910" />
                    <RANKING order="2" place="2" resultid="9674" />
                    <RANKING order="3" place="3" resultid="9838" />
                    <RANKING order="4" place="4" resultid="9911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6785" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="6786" agemax="-1" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9416" />
                    <RANKING order="2" place="2" resultid="9913" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12331" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12332" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="8362" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-01-01" gender="M" nation="POL" athleteid="9840">
              <RESULTS>
                <RESULT eventid="6077" points="739" swimtime="00:00:28.78" resultid="9841" heatid="11412" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="6306" points="672" reactiontime="+86" swimtime="00:01:06.23" resultid="9842" heatid="11474" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="636" reactiontime="+89" swimtime="00:00:32.61" resultid="9843" heatid="11536" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="6535" points="548" reactiontime="+79" swimtime="00:02:34.81" resultid="9844" heatid="11567" lane="0" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="532" swimtime="00:05:32.79" resultid="9845" heatid="11634" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:01:59.72" />
                    <SPLIT distance="200" swimtime="00:02:42.72" />
                    <SPLIT distance="250" swimtime="00:03:25.88" />
                    <SPLIT distance="300" swimtime="00:04:09.20" />
                    <SPLIT distance="350" swimtime="00:04:52.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8465" name="MKP Myślibórz">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Dąbrowski" birthdate="1998-01-01" gender="M" nation="POL" swrid="4352138" athleteid="8464">
              <RESULTS>
                <RESULT eventid="6077" points="811" reactiontime="+69" swimtime="00:00:24.59" resultid="8466" heatid="11418" lane="8" entrytime="00:00:24.71" />
                <RESULT eventid="6340" points="838" reactiontime="+66" swimtime="00:00:59.63" resultid="8467" heatid="11497" lane="1" entrytime="00:01:01.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="748" reactiontime="+72" swimtime="00:01:07.99" resultid="8468" heatid="11520" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="681" reactiontime="+65" swimtime="00:01:02.30" resultid="8469" heatid="11552" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="752" reactiontime="+66" swimtime="00:00:31.07" resultid="8470" heatid="11622" lane="1" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8499" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Bojanowicz" birthdate="1997-01-01" gender="M" nation="POL" athleteid="8498">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="8500" heatid="11414" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="8501" heatid="11432" lane="1" entrytime="00:02:34.00" />
                <RESULT eventid="6306" points="499" reactiontime="+89" swimtime="00:01:01.21" resultid="8502" heatid="11475" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="477" reactiontime="+79" swimtime="00:01:10.61" resultid="8503" heatid="11494" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8472" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Korzuchowski" birthdate="1999-01-01" gender="M" nation="POL" swrid="4598470" athleteid="8471">
              <RESULTS>
                <RESULT eventid="6077" points="609" reactiontime="+68" swimtime="00:00:27.05" resultid="8473" heatid="11415" lane="9" entrytime="00:00:27.10" />
                <RESULT eventid="6111" points="485" reactiontime="+77" swimtime="00:02:41.61" resultid="8474" heatid="11431" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:02:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="549" reactiontime="+65" swimtime="00:00:31.05" resultid="8475" heatid="11449" lane="8" entrytime="00:00:30.60" />
                <RESULT eventid="6340" points="523" swimtime="00:01:09.77" resultid="8476" heatid="11495" lane="9" entrytime="00:01:09.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="506" reactiontime="+60" swimtime="00:01:08.76" resultid="8477" heatid="11552" lane="3" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="365" reactiontime="+81" swimtime="00:06:15.44" resultid="8478" heatid="11579" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:05.83" />
                    <SPLIT distance="200" swimtime="00:02:53.61" />
                    <SPLIT distance="250" swimtime="00:03:49.81" />
                    <SPLIT distance="300" swimtime="00:04:46.56" />
                    <SPLIT distance="350" swimtime="00:05:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="470" reactiontime="+82" swimtime="00:01:09.85" resultid="8479" heatid="11594" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="506" reactiontime="+66" swimtime="00:02:35.45" resultid="8480" heatid="11605" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:56.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8510" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Kapczyński" birthdate="1966-01-01" gender="M" nation="POL" athleteid="8509">
              <RESULTS>
                <RESULT eventid="6272" points="525" reactiontime="+90" swimtime="00:03:20.81" resultid="8511" heatid="11456" lane="5" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:33.33" />
                    <SPLIT distance="150" swimtime="00:02:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="456" reactiontime="+86" swimtime="00:01:28.50" resultid="8512" heatid="11516" lane="4" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7873" name="Swim2Tri">
          <ATHLETES>
            <ATHLETE firstname="Marta" lastname="Mazur" birthdate="1984-10-05" gender="F" nation="POL" athleteid="7874">
              <RESULTS>
                <RESULT eventid="6255" points="437" reactiontime="+92" swimtime="00:03:24.45" resultid="7875" heatid="11453" lane="3" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:34.80" />
                    <SPLIT distance="150" swimtime="00:02:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="449" reactiontime="+91" swimtime="00:01:26.41" resultid="7876" heatid="11484" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="412" reactiontime="+94" swimtime="00:01:32.82" resultid="7877" heatid="11511" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="422" reactiontime="+92" swimtime="00:00:37.90" resultid="7878" heatid="11525" lane="2" entrytime="00:00:37.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8518" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Figarski" birthdate="1985-01-01" gender="M" nation="POL" swrid="4754698" athleteid="8517">
              <RESULTS>
                <RESULT eventid="6169" points="736" reactiontime="+91" swimtime="00:09:28.25" resultid="8519" heatid="11645" lane="2" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:38.97" />
                    <SPLIT distance="200" swimtime="00:02:14.26" />
                    <SPLIT distance="250" swimtime="00:02:50.01" />
                    <SPLIT distance="300" swimtime="00:03:25.90" />
                    <SPLIT distance="350" swimtime="00:04:01.27" />
                    <SPLIT distance="400" swimtime="00:04:36.95" />
                    <SPLIT distance="450" swimtime="00:05:12.60" />
                    <SPLIT distance="500" swimtime="00:05:48.34" />
                    <SPLIT distance="550" swimtime="00:06:24.54" />
                    <SPLIT distance="600" swimtime="00:07:00.79" />
                    <SPLIT distance="650" swimtime="00:07:37.64" />
                    <SPLIT distance="700" swimtime="00:08:14.54" />
                    <SPLIT distance="750" swimtime="00:08:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="580" reactiontime="+67" swimtime="00:00:29.34" resultid="8520" heatid="11449" lane="6" entrytime="00:00:29.80" />
                <RESULT eventid="6340" points="683" reactiontime="+89" swimtime="00:01:04.47" resultid="8521" heatid="11496" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="701" reactiontime="+68" swimtime="00:01:02.96" resultid="8522" heatid="11553" lane="8" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="668" reactiontime="+74" swimtime="00:02:19.04" resultid="8523" heatid="11606" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:43.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" clubid="7320" name="Uks Delfin Masters Tarnobrzeg">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Janus" birthdate="1987-10-02" gender="F" nation="POL" athleteid="7339">
              <RESULTS>
                <RESULT eventid="6059" points="710" reactiontime="+77" swimtime="00:00:29.34" resultid="7340" heatid="11400" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="6094" points="650" reactiontime="+89" swimtime="00:02:47.67" resultid="7341" heatid="11423" lane="2" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:09.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="678" reactiontime="+78" swimtime="00:01:05.77" resultid="7342" heatid="11465" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="708" reactiontime="+86" swimtime="00:01:14.23" resultid="7343" heatid="11485" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="497" reactiontime="+85" swimtime="00:01:27.18" resultid="7344" heatid="11511" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="583" reactiontime="+87" swimtime="00:02:33.36" resultid="7345" heatid="11558" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="524" reactiontime="+72" swimtime="00:02:57.12" resultid="7346" heatid="11600" lane="0" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:23.09" />
                    <SPLIT distance="150" swimtime="00:02:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="508" reactiontime="+85" swimtime="00:00:39.66" resultid="7347" heatid="11611" lane="2" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ślęczka" birthdate="1974-10-23" gender="M" nation="POL" license="500408700205" swrid="4992942" athleteid="7330">
              <RESULTS>
                <RESULT eventid="6077" points="730" reactiontime="+86" swimtime="00:00:26.50" resultid="7331" heatid="11411" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="6111" points="667" reactiontime="+82" swimtime="00:02:31.50" resultid="7332" heatid="11431" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="707" reactiontime="+70" swimtime="00:00:59.39" resultid="7333" heatid="11474" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="692" reactiontime="+80" swimtime="00:01:07.79" resultid="7334" heatid="11493" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="717" reactiontime="+80" swimtime="00:01:13.79" resultid="7335" heatid="11519" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="679" reactiontime="+80" swimtime="00:02:10.48" resultid="7336" heatid="11568" lane="5" entrytime="00:02:16.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:03.86" />
                    <SPLIT distance="150" swimtime="00:01:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="7337" heatid="11594" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="6704" points="753" reactiontime="+76" swimtime="00:00:33.28" resultid="7338" heatid="11620" lane="7" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Płaneta" birthdate="1974-09-12" gender="M" nation="POL" license="500408700210" swrid="4992944" athleteid="7321">
              <RESULTS>
                <RESULT eventid="6077" points="485" reactiontime="+82" swimtime="00:00:30.37" resultid="7322" heatid="11411" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="6169" points="398" reactiontime="+43" swimtime="00:11:46.24" resultid="7323" heatid="11646" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:03.18" />
                    <SPLIT distance="200" swimtime="00:02:46.89" />
                    <SPLIT distance="250" swimtime="00:03:31.30" />
                    <SPLIT distance="300" swimtime="00:04:15.80" />
                    <SPLIT distance="350" swimtime="00:05:00.42" />
                    <SPLIT distance="400" swimtime="00:05:44.67" />
                    <SPLIT distance="450" swimtime="00:06:29.05" />
                    <SPLIT distance="500" swimtime="00:07:13.93" />
                    <SPLIT distance="550" swimtime="00:07:59.14" />
                    <SPLIT distance="600" swimtime="00:08:44.70" />
                    <SPLIT distance="650" swimtime="00:09:30.18" />
                    <SPLIT distance="700" swimtime="00:10:16.43" />
                    <SPLIT distance="750" swimtime="00:11:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="395" reactiontime="+87" swimtime="00:00:37.96" resultid="7324" heatid="11447" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="6374" points="335" reactiontime="+83" swimtime="00:03:09.42" resultid="7325" heatid="11502" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                    <SPLIT distance="150" swimtime="00:02:19.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="360" reactiontime="+74" swimtime="00:01:23.51" resultid="7326" heatid="11551" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="376" reactiontime="+79" swimtime="00:02:38.90" resultid="7327" heatid="11566" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:17.83" />
                    <SPLIT distance="150" swimtime="00:01:59.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="364" reactiontime="+78" swimtime="00:03:04.19" resultid="7328" heatid="11603" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:02:18.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="398" reactiontime="+77" swimtime="00:05:34.24" resultid="7329" heatid="11634" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                    <SPLIT distance="200" swimtime="00:02:43.62" />
                    <SPLIT distance="250" swimtime="00:03:26.83" />
                    <SPLIT distance="300" swimtime="00:04:10.44" />
                    <SPLIT distance="350" swimtime="00:04:53.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" nation="POL" region="05" clubid="9532" name="UKS Nawa Skierniewice">
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Sarna" birthdate="1998-12-02" gender="F" nation="POL" license="100305600120" swrid="4476652" athleteid="9533">
              <RESULTS>
                <RESULT eventid="6220" points="587" reactiontime="+74" swimtime="00:00:34.63" resultid="9534" heatid="11438" lane="7" />
                <RESULT eventid="6323" points="483" reactiontime="+88" swimtime="00:01:20.50" resultid="9535" heatid="11481" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="529" reactiontime="+78" swimtime="00:00:34.44" resultid="9536" heatid="11523" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Dębski" birthdate="1998-08-01" gender="M" nation="POL" license="100305700340" swrid="4476651" athleteid="9537">
              <RESULTS>
                <RESULT eventid="6238" points="525" reactiontime="+71" swimtime="00:00:31.51" resultid="9538" heatid="11443" lane="3" />
                <RESULT eventid="6340" points="471" reactiontime="+74" swimtime="00:01:12.27" resultid="9539" heatid="11487" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="649" reactiontime="+80" swimtime="00:00:28.39" resultid="9540" heatid="11531" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Zyga" birthdate="1996-09-14" gender="F" nation="POL" license="100305600116" swrid="4287931" athleteid="9541">
              <RESULTS>
                <RESULT eventid="6255" points="629" reactiontime="+86" swimtime="00:02:59.26" resultid="9542" heatid="11451" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="632" reactiontime="+82" swimtime="00:01:22.32" resultid="9543" heatid="11508" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pamela" lastname="Broniarek" birthdate="1995-11-21" gender="F" nation="POL" license="100305600178" athleteid="9544">
              <RESULTS>
                <RESULT eventid="6289" points="542" reactiontime="+89" swimtime="00:01:08.80" resultid="9545" heatid="11462" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="402" reactiontime="+82" swimtime="00:03:06.78" resultid="9546" heatid="11498" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="150" swimtime="00:02:15.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="573" reactiontime="+91" swimtime="00:02:30.51" resultid="9547" heatid="11554" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8514" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Poloch" birthdate="1983-01-01" gender="M" nation="POL" athleteid="8513">
              <RESULTS>
                <RESULT eventid="6077" points="316" reactiontime="+93" swimtime="00:00:32.33" resultid="8515" heatid="11407" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="6306" points="267" swimtime="00:01:16.65" resultid="8516" heatid="11469" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6827" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Płonka" birthdate="1948-01-01" gender="M" nation="POL" swrid="4754750" athleteid="6826">
              <RESULTS>
                <RESULT eventid="6111" points="186" reactiontime="+108" swimtime="00:05:11.16" resultid="6828" heatid="11427" lane="8" entrytime="00:05:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.66" />
                    <SPLIT distance="100" swimtime="00:02:37.22" />
                    <SPLIT distance="150" swimtime="00:04:04.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="143" reactiontime="+124" swimtime="00:05:54.29" resultid="6829" heatid="11456" lane="9" entrytime="00:06:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.84" />
                    <SPLIT distance="100" swimtime="00:02:53.41" />
                    <SPLIT distance="150" swimtime="00:04:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="102" reactiontime="+107" swimtime="00:06:20.38" resultid="6830" heatid="11501" lane="0" entrytime="00:06:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.00" />
                    <SPLIT distance="100" swimtime="00:03:08.32" />
                    <SPLIT distance="150" swimtime="00:04:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="158" reactiontime="+121" swimtime="00:00:59.13" resultid="6831" heatid="11531" lane="3" entrytime="00:01:11.00" />
                <RESULT eventid="6569" points="168" reactiontime="+116" swimtime="00:11:57.12" resultid="6832" heatid="11576" lane="1" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.63" />
                    <SPLIT distance="100" swimtime="00:02:50.51" />
                    <SPLIT distance="150" swimtime="00:04:32.09" />
                    <SPLIT distance="250" swimtime="00:07:43.53" />
                    <SPLIT distance="300" swimtime="00:09:18.22" />
                    <SPLIT distance="350" swimtime="00:10:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="112" reactiontime="+125" swimtime="00:02:36.68" resultid="6833" heatid="11590" lane="8" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="130" reactiontime="+116" swimtime="00:01:10.11" resultid="6834" heatid="11615" lane="3" entrytime="00:01:01.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7116" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Kamiński" birthdate="1965-01-01" gender="M" nation="POL" athleteid="7115">
              <RESULTS>
                <RESULT eventid="6077" points="500" reactiontime="+58" swimtime="00:00:32.79" resultid="7117" heatid="11406" lane="9" entrytime="00:00:36.95" />
                <RESULT eventid="6238" points="432" reactiontime="+80" swimtime="00:00:38.80" resultid="7118" heatid="11445" lane="5" entrytime="00:00:43.45" />
                <RESULT eventid="6306" points="521" reactiontime="+84" swimtime="00:01:12.10" resultid="7119" heatid="11471" lane="8" entrytime="00:01:17.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="440" reactiontime="+84" swimtime="00:01:25.14" resultid="7120" heatid="11550" lane="1" entrytime="00:01:33.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="482" reactiontime="+82" swimtime="00:03:02.69" resultid="7121" heatid="11603" lane="4" entrytime="00:03:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:16.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7248" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Orczyk" birthdate="1995-01-01" gender="M" nation="POL" swrid="4195155" athleteid="7247">
              <RESULTS>
                <RESULT eventid="6077" points="384" reactiontime="+76" swimtime="00:00:31.41" resultid="7249" heatid="11410" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="6340" points="670" swimtime="00:01:03.07" resultid="7250" heatid="11496" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="745" reactiontime="+81" swimtime="00:01:08.42" resultid="7251" heatid="11521" lane="7" entrytime="00:01:07.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="733" swimtime="00:00:31.34" resultid="7252" heatid="11622" lane="4" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7937" name="Masters Łódź">
          <ATHLETES>
            <ATHLETE firstname="Artur" lastname="Frąckowiak" birthdate="1978-06-28" gender="M" nation="POL" license="503605700020" swrid="5279744" athleteid="7966">
              <RESULTS>
                <RESULT eventid="6077" points="619" reactiontime="+75" swimtime="00:00:27.22" resultid="7967" heatid="11413" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="6111" points="614" reactiontime="+83" swimtime="00:02:30.45" resultid="7968" heatid="11431" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:56.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7969" heatid="11476" lane="1" entrytime="00:01:01.00" />
                <RESULT eventid="6340" points="698" reactiontime="+79" swimtime="00:01:07.41" resultid="7970" heatid="11494" lane="0" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="630" reactiontime="+75" swimtime="00:00:29.31" resultid="7971" heatid="11539" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7972" heatid="11635" lane="7" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olejarczyk" birthdate="1979-06-12" gender="M" nation="POL" license="503605700007" swrid="4992959" athleteid="7938">
              <RESULTS>
                <RESULT eventid="6077" points="661" reactiontime="+74" swimtime="00:00:26.64" resultid="7939" heatid="11415" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="6306" points="636" reactiontime="+82" swimtime="00:00:59.61" resultid="7940" heatid="11476" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="507" reactiontime="+86" swimtime="00:02:38.08" resultid="7941" heatid="11503" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="667" swimtime="00:00:28.75" resultid="7942" heatid="11538" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="6535" points="526" reactiontime="+77" swimtime="00:02:20.01" resultid="7943" heatid="11567" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="635" reactiontime="+76" swimtime="00:01:05.87" resultid="7944" heatid="11594" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Michniewski" birthdate="1983-04-11" gender="M" nation="POL" license="503605700012" swrid="5537479" athleteid="7973">
              <RESULTS>
                <RESULT eventid="6077" points="573" reactiontime="+85" swimtime="00:00:26.52" resultid="7974" heatid="11415" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="6111" points="600" reactiontime="+89" swimtime="00:02:30.90" resultid="7975" heatid="11429" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:54.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="630" reactiontime="+86" swimtime="00:02:43.97" resultid="7976" heatid="11458" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="639" reactiontime="+77" swimtime="00:01:05.92" resultid="7977" heatid="11495" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="656" reactiontime="+84" swimtime="00:01:13.07" resultid="7978" heatid="11520" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="509" reactiontime="+73" swimtime="00:00:29.59" resultid="7979" heatid="11538" lane="5" entrytime="00:00:29.20" />
                <RESULT eventid="6704" points="627" reactiontime="+74" swimtime="00:00:33.71" resultid="7980" heatid="11621" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Grzeszczuk" birthdate="1991-02-25" gender="F" nation="POL" license="503605600035" swrid="4806334" athleteid="7961">
              <RESULTS>
                <RESULT eventid="6323" points="680" reactiontime="+68" swimtime="00:01:13.69" resultid="7962" heatid="11485" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="746" reactiontime="+71" swimtime="00:01:16.35" resultid="7963" heatid="11512" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="731" reactiontime="+68" swimtime="00:00:31.29" resultid="7964" heatid="11527" lane="5" entrytime="00:00:32.20" />
                <RESULT eventid="6687" points="777" swimtime="00:00:34.10" resultid="7965" heatid="11612" lane="4" entrytime="00:00:34.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Woźniak" birthdate="1981-08-25" gender="M" nation="POL" license="503605700034" swrid="5484423" athleteid="7945">
              <RESULTS>
                <RESULT eventid="6238" points="739" reactiontime="+61" swimtime="00:00:30.02" resultid="7946" heatid="11449" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="6340" points="644" reactiontime="+79" swimtime="00:01:09.26" resultid="7947" heatid="11494" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="611" reactiontime="+92" swimtime="00:00:29.61" resultid="7948" heatid="11531" lane="7" />
                <RESULT eventid="6501" points="711" reactiontime="+68" swimtime="00:01:06.17" resultid="7949" heatid="11553" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="747" reactiontime="+69" swimtime="00:02:23.74" resultid="7950" heatid="11606" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Kruszyna-Kotulski" birthdate="1979-05-25" gender="M" nation="POL" license="503605700044" swrid="4417017" athleteid="7957">
              <RESULTS>
                <RESULT eventid="6238" points="373" reactiontime="+78" swimtime="00:00:37.71" resultid="7958" heatid="11446" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="6340" points="510" reactiontime="+74" swimtime="00:01:14.83" resultid="7959" heatid="11491" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="574" reactiontime="+44" swimtime="00:00:30.23" resultid="7960" heatid="11538" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+78" swimtime="00:01:47.93" resultid="9835" heatid="11584" lane="2" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="100" swimtime="00:00:53.86" />
                    <SPLIT distance="150" swimtime="00:01:21.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7966" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="7973" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="7945" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="7938" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="6779" status="DNS" swimtime="00:00:00.00" resultid="9836" heatid="12331" lane="4" entrytime="00:01:59.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7945" number="1" />
                    <RELAYPOSITION athleteid="7973" number="2" />
                    <RELAYPOSITION athleteid="7938" number="3" />
                    <RELAYPOSITION athleteid="7957" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7188" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Chmielowiec" birthdate="2000-01-01" gender="M" nation="POL" swrid="4750258" athleteid="7187">
              <RESULTS>
                <RESULT eventid="6077" points="754" reactiontime="+68" swimtime="00:00:25.20" resultid="7189" heatid="11417" lane="0" entrytime="00:00:25.44" />
                <RESULT eventid="6467" points="852" reactiontime="+67" swimtime="00:00:25.92" resultid="7190" heatid="11542" lane="8" entrytime="00:00:25.04" />
                <RESULT eventid="6636" points="703" reactiontime="+69" swimtime="00:01:01.09" resultid="7191" heatid="11597" lane="0" entrytime="00:00:57.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8403" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Angelika" lastname="Wróbel" birthdate="1997-01-01" gender="F" nation="POL" swrid="4373387" athleteid="8402">
              <RESULTS>
                <RESULT eventid="6059" points="717" reactiontime="+88" swimtime="00:00:28.25" resultid="8404" heatid="11400" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="6289" points="731" reactiontime="+85" swimtime="00:01:02.28" resultid="8405" heatid="11466" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="8406" heatid="11528" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="6518" points="735" reactiontime="+87" swimtime="00:02:18.54" resultid="8407" heatid="11559" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" status="DNS" swimtime="00:00:00.00" resultid="8408" heatid="11588" lane="7" entrytime="00:01:13.00" />
                <RESULT eventid="6721" points="675" reactiontime="+88" swimtime="00:05:05.28" resultid="8409" heatid="11628" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="150" swimtime="00:01:52.27" />
                    <SPLIT distance="200" swimtime="00:02:32.04" />
                    <SPLIT distance="250" swimtime="00:03:11.56" />
                    <SPLIT distance="300" swimtime="00:03:50.76" />
                    <SPLIT distance="350" swimtime="00:04:28.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8416" name="3Waters">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="Borkowska" birthdate="1975-01-01" gender="F" nation="POL" athleteid="8415">
              <RESULTS>
                <RESULT eventid="6059" points="612" reactiontime="+75" swimtime="00:00:31.68" resultid="8417" heatid="11398" lane="2" entrytime="00:00:33.30" />
                <RESULT eventid="6289" points="558" reactiontime="+76" swimtime="00:01:12.40" resultid="8418" heatid="11464" lane="2" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="523" reactiontime="+78" swimtime="00:01:25.78" resultid="8419" heatid="11484" lane="9" entrytime="00:01:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="498" reactiontime="+71" swimtime="00:00:37.87" resultid="8420" heatid="11525" lane="1" entrytime="00:00:39.10" />
                <RESULT eventid="6687" points="547" reactiontime="+80" swimtime="00:00:42.50" resultid="8421" heatid="11611" lane="8" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7193" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Angelika" lastname="Wojtaszek" birthdate="1997-01-01" gender="F" nation="POL" athleteid="7192">
              <RESULTS>
                <RESULT eventid="6289" status="DNS" swimtime="00:00:00.00" resultid="7194" heatid="11465" lane="0" entrytime="00:01:12.10" />
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="7195" heatid="11526" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="6618" status="DNS" swimtime="00:00:00.00" resultid="7196" heatid="11587" lane="6" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8624" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Szewczyk" birthdate="1996-01-01" gender="M" nation="POL" swrid="4115546" athleteid="8623">
              <RESULTS>
                <RESULT eventid="6467" points="599" reactiontime="+62" swimtime="00:00:28.11" resultid="8625" heatid="11540" lane="9" entrytime="00:00:28.20" />
                <RESULT eventid="6704" points="662" reactiontime="+65" swimtime="00:00:32.41" resultid="8626" heatid="11622" lane="7" entrytime="00:00:32.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6906" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Szklarzewski" birthdate="1985-01-01" gender="M" nation="POL" athleteid="6905">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="6907" heatid="11416" lane="6" entrytime="00:00:25.90" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="6908" heatid="11538" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="6909" heatid="11477" lane="3" entrytime="00:00:58.00" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="6910" heatid="11569" lane="7" entrytime="00:02:15.00" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="6911" heatid="11593" lane="3" entrytime="00:01:12.00" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="6912" heatid="11619" lane="5" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="9177" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Wawrzyniec" lastname="Manczak" birthdate="1948-06-03" gender="M" nation="POL" license="102202700108" swrid="4186189" athleteid="9183">
              <RESULTS>
                <RESULT eventid="6238" points="510" reactiontime="+78" swimtime="00:00:43.38" resultid="9184" heatid="11442" lane="5" />
                <RESULT eventid="6501" points="422" reactiontime="+89" swimtime="00:01:40.02" resultid="9185" heatid="11547" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="546" reactiontime="+94" swimtime="00:03:42.60" resultid="9186" heatid="11601" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.43" />
                    <SPLIT distance="100" swimtime="00:01:49.61" />
                    <SPLIT distance="150" swimtime="00:02:48.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ciężki" birthdate="1994-09-30" gender="M" nation="POL" license="102202700137" swrid="4289450" athleteid="9178">
              <RESULTS>
                <RESULT eventid="6238" points="591" reactiontime="+70" swimtime="00:00:29.85" resultid="9179" heatid="11449" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="6306" points="639" reactiontime="+80" swimtime="00:00:56.40" resultid="9180" heatid="11478" lane="6" entrytime="00:00:55.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="609" reactiontime="+73" swimtime="00:01:04.92" resultid="9181" heatid="11552" lane="4" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="545" reactiontime="+66" swimtime="00:02:22.24" resultid="9182" heatid="11606" lane="1" entrytime="00:02:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:08.48" />
                    <SPLIT distance="150" swimtime="00:01:45.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="9187">
              <RESULTS>
                <RESULT eventid="6501" points="130" reactiontime="+95" swimtime="00:01:59.19" resultid="9188" heatid="11549" lane="8" entrytime="00:01:55.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="150" reactiontime="+106" swimtime="00:04:21.57" resultid="9189" heatid="11602" lane="6" entrytime="00:04:12.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.78" />
                    <SPLIT distance="100" swimtime="00:02:07.08" />
                    <SPLIT distance="150" swimtime="00:03:13.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9190" heatid="11630" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" clubid="7422" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Grzeszewski" birthdate="1953-09-25" gender="M" nation="POL" swrid="4754656" athleteid="7423">
              <RESULTS>
                <RESULT eventid="6111" points="447" reactiontime="+69" swimtime="00:03:27.38" resultid="7424" heatid="11428" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:01:40.56" />
                    <SPLIT distance="150" swimtime="00:02:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="590" reactiontime="+81" swimtime="00:03:36.62" resultid="7425" heatid="11457" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:45.39" />
                    <SPLIT distance="150" swimtime="00:02:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="497" reactiontime="+78" swimtime="00:01:37.09" resultid="7426" heatid="11516" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="450" reactiontime="+80" swimtime="00:00:39.86" resultid="7427" heatid="11534" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="6704" points="550" swimtime="00:00:41.23" resultid="7428" heatid="11618" lane="8" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Szozda" birthdate="1960-01-12" gender="M" nation="POL" swrid="4461547" athleteid="7440">
              <RESULTS>
                <RESULT eventid="6111" points="551" reactiontime="+98" swimtime="00:03:06.49" resultid="7441" heatid="11428" lane="4" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                    <SPLIT distance="150" swimtime="00:02:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="579" reactiontime="+96" swimtime="00:01:21.89" resultid="7442" heatid="11491" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="546" reactiontime="+98" swimtime="00:01:30.36" resultid="7443" heatid="11517" lane="5" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="466" reactiontime="+96" swimtime="00:01:27.15" resultid="7444" heatid="11550" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="443" swimtime="00:01:28.41" resultid="7445" heatid="11592" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="540" reactiontime="+96" swimtime="00:00:40.19" resultid="7446" heatid="11617" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Serbin" birthdate="1966-08-10" gender="F" nation="POL" swrid="4302596" athleteid="7447">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6186" points="848" reactiontime="+82" swimtime="00:20:52.11" resultid="7448" heatid="11650" lane="5" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                    <SPLIT distance="200" swimtime="00:02:40.59" />
                    <SPLIT distance="250" swimtime="00:03:22.34" />
                    <SPLIT distance="300" swimtime="00:04:04.42" />
                    <SPLIT distance="350" swimtime="00:04:46.19" />
                    <SPLIT distance="400" swimtime="00:05:27.91" />
                    <SPLIT distance="450" swimtime="00:06:09.36" />
                    <SPLIT distance="500" swimtime="00:06:50.86" />
                    <SPLIT distance="550" swimtime="00:07:32.26" />
                    <SPLIT distance="600" swimtime="00:08:13.60" />
                    <SPLIT distance="650" swimtime="00:08:55.21" />
                    <SPLIT distance="700" swimtime="00:09:36.79" />
                    <SPLIT distance="750" swimtime="00:10:18.47" />
                    <SPLIT distance="800" swimtime="00:11:00.28" />
                    <SPLIT distance="850" swimtime="00:11:42.29" />
                    <SPLIT distance="900" swimtime="00:12:24.23" />
                    <SPLIT distance="950" swimtime="00:13:06.27" />
                    <SPLIT distance="1000" swimtime="00:13:48.32" />
                    <SPLIT distance="1050" swimtime="00:14:30.48" />
                    <SPLIT distance="1100" swimtime="00:15:12.82" />
                    <SPLIT distance="1150" swimtime="00:15:55.38" />
                    <SPLIT distance="1200" swimtime="00:16:37.88" />
                    <SPLIT distance="1250" swimtime="00:17:20.77" />
                    <SPLIT distance="1300" swimtime="00:18:03.49" />
                    <SPLIT distance="1350" swimtime="00:18:46.23" />
                    <SPLIT distance="1400" swimtime="00:19:28.96" />
                    <SPLIT distance="1450" swimtime="00:20:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="687" reactiontime="+83" swimtime="00:01:11.06" resultid="7449" heatid="11465" lane="2" entrytime="00:01:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="744" reactiontime="+78" swimtime="00:02:32.03" resultid="7450" heatid="11559" lane="1" entrytime="00:02:28.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:01:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="768" reactiontime="+82" swimtime="00:05:18.17" resultid="7451" heatid="11628" lane="2" entrytime="00:05:08.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:56.33" />
                    <SPLIT distance="200" swimtime="00:02:36.64" />
                    <SPLIT distance="250" swimtime="00:03:16.99" />
                    <SPLIT distance="300" swimtime="00:03:57.67" />
                    <SPLIT distance="350" swimtime="00:04:38.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Chmurski" birthdate="1987-09-23" gender="M" nation="POL" swrid="4060941" athleteid="7429">
              <RESULTS>
                <RESULT eventid="6077" points="677" reactiontime="+77" swimtime="00:00:25.08" resultid="7430" heatid="11417" lane="8" entrytime="00:00:25.40" />
                <RESULT eventid="6238" points="606" reactiontime="+82" swimtime="00:00:28.92" resultid="7431" heatid="11449" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="6340" points="674" reactiontime="+78" swimtime="00:01:04.77" resultid="7432" heatid="11496" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="688" reactiontime="+77" swimtime="00:02:06.25" resultid="7433" heatid="11570" lane="0" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:01:00.65" />
                    <SPLIT distance="150" swimtime="00:01:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="751" reactiontime="+76" swimtime="00:04:26.55" resultid="7434" heatid="11637" lane="7" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                    <SPLIT distance="150" swimtime="00:01:38.76" />
                    <SPLIT distance="200" swimtime="00:02:13.54" />
                    <SPLIT distance="250" swimtime="00:02:48.03" />
                    <SPLIT distance="300" swimtime="00:03:22.21" />
                    <SPLIT distance="350" swimtime="00:03:55.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11342" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" athleteid="9846">
              <RESULTS>
                <RESULT eventid="6077" points="694" reactiontime="+71" swimtime="00:00:26.95" resultid="9847" heatid="11415" lane="5" entrytime="00:00:26.44" />
                <RESULT eventid="6306" points="729" reactiontime="+76" swimtime="00:00:58.79" resultid="9848" heatid="11477" lane="9" entrytime="00:00:59.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="680" reactiontime="+74" swimtime="00:02:10.42" resultid="9849" heatid="11569" lane="5" entrytime="00:02:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:01.51" />
                    <SPLIT distance="150" swimtime="00:01:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="649" reactiontime="+78" swimtime="00:04:43.96" resultid="9850" heatid="11637" lane="1" entrytime="00:04:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="150" swimtime="00:01:42.98" />
                    <SPLIT distance="200" swimtime="00:02:20.12" />
                    <SPLIT distance="250" swimtime="00:02:57.11" />
                    <SPLIT distance="300" swimtime="00:03:34.55" />
                    <SPLIT distance="350" swimtime="00:04:10.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" clubid="7886" name="UKS Wodnik 29 Katowice">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Koenig" birthdate="1987-01-01" gender="F" nation="POL" swrid="5464149" athleteid="7901">
              <RESULTS>
                <RESULT eventid="6059" status="DNS" swimtime="00:00:00.00" resultid="7902" heatid="11395" lane="4" entrytime="00:00:59.00" />
                <RESULT eventid="6255" points="147" swimtime="00:04:53.60" resultid="7903" heatid="11452" lane="4" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.57" />
                    <SPLIT distance="100" swimtime="00:02:15.88" />
                    <SPLIT distance="150" swimtime="00:03:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="143" swimtime="00:02:11.84" resultid="7904" heatid="11510" lane="2" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="143" swimtime="00:01:00.47" resultid="7905" heatid="11609" lane="3" entrytime="00:00:59.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ilnicki" birthdate="1956-01-01" gender="M" nation="POL" swrid="5484406" athleteid="7906">
              <RESULTS>
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7907" heatid="11428" lane="1" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:04:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7908" heatid="11468" lane="1" entrytime="00:01:45.00" />
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="7909" heatid="11516" lane="9" entrytime="00:01:46.70" entrycourse="SCM" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7910" heatid="11616" lane="2" entrytime="00:00:46.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Dąbrowski" birthdate="1988-02-20" gender="M" nation="POL" swrid="4092977" athleteid="9676">
              <RESULTS>
                <RESULT eventid="6077" points="766" reactiontime="+80" swimtime="00:00:24.18" resultid="9677" heatid="11418" lane="7" entrytime="00:00:24.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Mroziński" birthdate="1959-01-01" gender="M" nation="POL" athleteid="9866">
              <RESULTS>
                <RESULT eventid="6077" points="618" reactiontime="+79" swimtime="00:00:31.51" resultid="9867" heatid="11409" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="6272" points="733" reactiontime="+85" swimtime="00:03:04.02" resultid="9868" heatid="11458" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:26.64" />
                    <SPLIT distance="150" swimtime="00:02:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="668" reactiontime="+80" swimtime="00:01:18.09" resultid="9869" heatid="11492" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="720" reactiontime="+81" swimtime="00:01:22.39" resultid="9870" heatid="11519" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="727" reactiontime="+78" swimtime="00:00:36.41" resultid="9871" heatid="11620" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Władyka" birthdate="2002-01-01" gender="M" nation="POL" swrid="4780552" athleteid="9819">
              <RESULTS>
                <RESULT eventid="6704" points="926" reactiontime="+64" swimtime="00:00:28.99" resultid="9820" heatid="11623" lane="5" entrytime="00:00:28.05" entrycourse="SCM" />
                <RESULT eventid="6433" points="907" reactiontime="+64" swimtime="00:01:03.76" resultid="9821" heatid="11521" lane="5" entrytime="00:01:01.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Mróz" birthdate="1979-01-01" gender="F" nation="POL" athleteid="9872">
              <RESULTS>
                <RESULT eventid="6059" points="503" swimtime="00:00:33.03" resultid="9873" heatid="11399" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="6094" points="550" reactiontime="+86" swimtime="00:02:59.13" resultid="9874" heatid="11422" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:02:19.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="514" reactiontime="+86" swimtime="00:01:13.00" resultid="9875" heatid="11465" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="540" reactiontime="+74" swimtime="00:01:23.64" resultid="9876" heatid="11484" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="482" reactiontime="+83" swimtime="00:00:37.36" resultid="9877" heatid="11526" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="6518" points="548" reactiontime="+92" swimtime="00:02:38.02" resultid="9878" heatid="11557" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="589" swimtime="00:05:30.27" resultid="9879" heatid="11627" lane="1" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:01.22" />
                    <SPLIT distance="200" swimtime="00:02:43.67" />
                    <SPLIT distance="250" swimtime="00:03:25.73" />
                    <SPLIT distance="300" swimtime="00:04:07.66" />
                    <SPLIT distance="350" swimtime="00:04:49.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7650" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" swrid="5471789" athleteid="7736">
              <RESULTS>
                <RESULT eventid="6636" points="679" reactiontime="+84" swimtime="00:01:06.59" resultid="7737" heatid="11594" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="571" reactiontime="+67" swimtime="00:02:38.53" resultid="7738" heatid="11605" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" swrid="4258728" athleteid="7788">
              <RESULTS>
                <RESULT eventid="6059" points="836" reactiontime="+63" swimtime="00:00:26.84" resultid="7789" heatid="11401" lane="5" entrytime="00:00:26.94" />
                <RESULT eventid="6289" points="882" swimtime="00:00:58.51" resultid="7790" heatid="11466" lane="4" entrytime="00:00:58.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="780" reactiontime="+66" swimtime="00:01:09.28" resultid="7791" heatid="11486" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="773" reactiontime="+65" swimtime="00:00:30.06" resultid="7792" heatid="11528" lane="3" entrytime="00:00:29.35" />
                <RESULT eventid="6518" points="874" reactiontime="+67" swimtime="00:02:10.75" resultid="7793" heatid="11559" lane="5" entrytime="00:02:13.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:01:03.44" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="638" reactiontime="+70" swimtime="00:00:36.68" resultid="7794" heatid="11608" lane="6" />
                <RESULT eventid="6721" points="884" reactiontime="+67" swimtime="00:04:39.08" resultid="7795" heatid="11624" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                    <SPLIT distance="150" swimtime="00:01:41.40" />
                    <SPLIT distance="200" swimtime="00:02:17.45" />
                    <SPLIT distance="250" swimtime="00:02:53.90" />
                    <SPLIT distance="300" swimtime="00:03:30.65" />
                    <SPLIT distance="350" swimtime="00:04:06.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Żemier" birthdate="1982-11-09" gender="M" nation="POL" swrid="4228280" athleteid="7701">
              <RESULTS>
                <RESULT eventid="6077" points="834" swimtime="00:00:24.65" resultid="7702" heatid="11403" lane="9" />
                <RESULT eventid="6111" points="814" reactiontime="+72" swimtime="00:02:16.92" resultid="7703" heatid="11425" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="909" reactiontime="+66" swimtime="00:00:28.02" resultid="7704" heatid="11449" lane="4" entrytime="00:00:27.99" />
                <RESULT eventid="6340" points="917" reactiontime="+76" swimtime="00:01:01.56" resultid="7705" heatid="11497" lane="8" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="783" reactiontime="+74" swimtime="00:00:27.26" resultid="7706" heatid="11530" lane="2" />
                <RESULT eventid="6501" points="908" reactiontime="+63" swimtime="00:01:00.98" resultid="7707" heatid="11553" lane="7" entrytime="00:01:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="809" swimtime="00:01:00.76" resultid="7708" heatid="11589" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="871" reactiontime="+68" swimtime="00:02:16.61" resultid="7709" heatid="11606" lane="4" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="150" swimtime="00:01:41.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Mikicin" birthdate="1993-10-18" gender="M" nation="POL" swrid="4801125" athleteid="7734">
              <RESULTS>
                <RESULT eventid="6238" points="849" reactiontime="+56" swimtime="00:00:26.45" resultid="7735" heatid="11450" lane="4" entrytime="00:00:24.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" swrid="4806379" athleteid="7696">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6203" points="905" reactiontime="+76" swimtime="00:16:41.10" resultid="7697" heatid="11652" lane="5" entrytime="00:17:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:01.48" />
                    <SPLIT distance="150" swimtime="00:01:34.84" />
                    <SPLIT distance="200" swimtime="00:02:08.42" />
                    <SPLIT distance="250" swimtime="00:02:41.68" />
                    <SPLIT distance="300" swimtime="00:03:15.15" />
                    <SPLIT distance="350" swimtime="00:03:48.78" />
                    <SPLIT distance="400" swimtime="00:04:22.36" />
                    <SPLIT distance="450" swimtime="00:04:55.64" />
                    <SPLIT distance="500" swimtime="00:05:28.97" />
                    <SPLIT distance="550" swimtime="00:06:02.17" />
                    <SPLIT distance="600" swimtime="00:06:35.78" />
                    <SPLIT distance="650" swimtime="00:07:09.41" />
                    <SPLIT distance="700" swimtime="00:07:43.12" />
                    <SPLIT distance="750" swimtime="00:08:16.83" />
                    <SPLIT distance="800" swimtime="00:08:50.43" />
                    <SPLIT distance="850" swimtime="00:09:24.09" />
                    <SPLIT distance="900" swimtime="00:09:58.07" />
                    <SPLIT distance="950" swimtime="00:10:31.75" />
                    <SPLIT distance="1000" swimtime="00:11:05.75" />
                    <SPLIT distance="1050" swimtime="00:11:39.69" />
                    <SPLIT distance="1100" swimtime="00:12:13.56" />
                    <SPLIT distance="1150" swimtime="00:12:47.72" />
                    <SPLIT distance="1200" swimtime="00:13:21.93" />
                    <SPLIT distance="1250" swimtime="00:13:55.41" />
                    <SPLIT distance="1300" swimtime="00:14:29.10" />
                    <SPLIT distance="1350" swimtime="00:15:02.64" />
                    <SPLIT distance="1400" swimtime="00:15:36.62" />
                    <SPLIT distance="1450" swimtime="00:16:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="945" reactiontime="+73" swimtime="00:02:21.01" resultid="7698" heatid="11460" lane="5" entrytime="00:02:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:07.53" />
                    <SPLIT distance="150" swimtime="00:01:43.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="911" reactiontime="+71" swimtime="00:04:38.07" resultid="7699" heatid="11579" lane="4" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="100" swimtime="00:01:02.79" />
                    <SPLIT distance="150" swimtime="00:01:41.76" />
                    <SPLIT distance="200" swimtime="00:02:19.25" />
                    <SPLIT distance="250" swimtime="00:02:56.69" />
                    <SPLIT distance="300" swimtime="00:03:34.78" />
                    <SPLIT distance="350" swimtime="00:04:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="937" swimtime="00:04:07.53" resultid="7700" heatid="11638" lane="4" entrytime="00:04:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:00:59.54" />
                    <SPLIT distance="150" swimtime="00:01:31.09" />
                    <SPLIT distance="200" swimtime="00:02:03.14" />
                    <SPLIT distance="250" swimtime="00:02:35.02" />
                    <SPLIT distance="300" swimtime="00:03:07.23" />
                    <SPLIT distance="350" swimtime="00:03:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" swrid="5416809" athleteid="7748">
              <RESULTS>
                <RESULT eventid="6077" points="547" swimtime="00:00:29.18" resultid="7749" heatid="11409" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="6306" points="551" swimtime="00:01:04.55" resultid="7750" heatid="11472" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="530" reactiontime="+88" swimtime="00:00:31.73" resultid="7751" heatid="11534" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="6535" points="482" reactiontime="+87" swimtime="00:02:26.25" resultid="7752" heatid="11567" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="432" reactiontime="+82" swimtime="00:01:17.41" resultid="7753" heatid="11590" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7754" heatid="11634" lane="9" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" swrid="4251116" athleteid="7755">
              <RESULTS>
                <RESULT eventid="6059" points="530" reactiontime="+83" swimtime="00:00:31.99" resultid="7756" heatid="11399" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="6289" points="506" swimtime="00:01:12.10" resultid="7757" heatid="11465" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="423" swimtime="00:01:26.33" resultid="7758" heatid="11483" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="367" reactiontime="+89" swimtime="00:01:29.79" resultid="7759" heatid="11545" lane="1" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="475" reactiontime="+89" swimtime="00:02:41.06" resultid="7760" heatid="11558" lane="9" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="446" reactiontime="+103" swimtime="00:05:52.64" resultid="7761" heatid="11624" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:06.76" />
                    <SPLIT distance="200" swimtime="00:02:53.20" />
                    <SPLIT distance="250" swimtime="00:03:39.21" />
                    <SPLIT distance="300" swimtime="00:04:25.51" />
                    <SPLIT distance="350" swimtime="00:05:11.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Fluder" birthdate="1986-03-01" gender="M" nation="POL" swrid="4073249" athleteid="7691">
              <RESULTS>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7692" heatid="11540" lane="3" entrytime="00:00:27.70" />
                <RESULT eventid="6535" points="763" reactiontime="+78" swimtime="00:02:01.95" resultid="7693" heatid="11571" lane="8" entrytime="00:02:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="100" swimtime="00:01:00.04" />
                    <SPLIT distance="150" swimtime="00:01:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="683" swimtime="00:01:02.67" resultid="7694" heatid="11595" lane="6" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="797" reactiontime="+83" swimtime="00:04:21.34" resultid="7695" heatid="11638" lane="2" entrytime="00:04:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:02.76" />
                    <SPLIT distance="150" swimtime="00:01:35.79" />
                    <SPLIT distance="200" swimtime="00:02:09.78" />
                    <SPLIT distance="250" swimtime="00:02:43.68" />
                    <SPLIT distance="300" swimtime="00:03:17.40" />
                    <SPLIT distance="350" swimtime="00:03:50.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" swrid="5425564" athleteid="7681">
              <RESULTS>
                <RESULT eventid="6077" points="808" reactiontime="+72" swimtime="00:00:27.94" resultid="7682" heatid="11413" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="6272" points="851" reactiontime="+76" swimtime="00:02:50.96" resultid="7683" heatid="11459" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="877" reactiontime="+72" swimtime="00:01:08.67" resultid="7684" heatid="11495" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6433" points="761" reactiontime="+79" swimtime="00:01:14.60" resultid="7685" heatid="11520" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6704" points="767" reactiontime="+76" swimtime="00:00:33.31" resultid="7686" heatid="11621" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" swrid="5240601" athleteid="7718">
              <RESULTS>
                <RESULT eventid="6094" points="589" swimtime="00:03:02.95" resultid="7719" heatid="11423" lane="9" entrytime="00:03:02.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:30.12" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="540" swimtime="00:11:58.28" resultid="7720" heatid="11643" lane="1" entrytime="00:11:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:07.31" />
                    <SPLIT distance="200" swimtime="00:02:52.52" />
                    <SPLIT distance="250" swimtime="00:03:38.39" />
                    <SPLIT distance="300" swimtime="00:04:23.84" />
                    <SPLIT distance="350" swimtime="00:05:09.45" />
                    <SPLIT distance="400" swimtime="00:05:54.93" />
                    <SPLIT distance="450" swimtime="00:06:40.46" />
                    <SPLIT distance="500" swimtime="00:07:25.83" />
                    <SPLIT distance="550" swimtime="00:08:11.71" />
                    <SPLIT distance="600" swimtime="00:08:57.96" />
                    <SPLIT distance="650" swimtime="00:09:44.20" />
                    <SPLIT distance="700" swimtime="00:10:30.06" />
                    <SPLIT distance="750" swimtime="00:11:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="716" reactiontime="+86" swimtime="00:03:07.94" resultid="7721" heatid="11454" lane="2" entrytime="00:03:04.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:29.38" />
                    <SPLIT distance="150" swimtime="00:02:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="593" reactiontime="+86" swimtime="00:01:22.19" resultid="7722" heatid="11484" lane="5" entrytime="00:01:23.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="681" reactiontime="+83" swimtime="00:01:27.62" resultid="7723" heatid="11512" lane="8" entrytime="00:01:23.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="578" reactiontime="+86" swimtime="00:02:40.79" resultid="7724" heatid="11558" lane="2" entrytime="00:02:41.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:00.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="833" reactiontime="+75" swimtime="00:00:38.05" resultid="7725" heatid="11612" lane="8" entrytime="00:00:38.11" />
                <RESULT eventid="6721" points="604" reactiontime="+84" swimtime="00:05:38.59" resultid="7726" heatid="11627" lane="3" entrytime="00:05:38.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                    <SPLIT distance="200" swimtime="00:02:47.97" />
                    <SPLIT distance="250" swimtime="00:03:30.46" />
                    <SPLIT distance="300" swimtime="00:04:13.44" />
                    <SPLIT distance="350" swimtime="00:04:56.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Matyszewski" birthdate="1971-10-11" gender="M" nation="POL" athleteid="7779">
              <RESULTS>
                <RESULT eventid="6077" points="374" swimtime="00:00:33.99" resultid="7780" heatid="11408" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="6111" points="286" reactiontime="+80" swimtime="00:03:20.27" resultid="7781" heatid="11426" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:37.83" />
                    <SPLIT distance="150" swimtime="00:02:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="455" reactiontime="+71" swimtime="00:03:21.06" resultid="7782" heatid="11457" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.40" />
                    <SPLIT distance="100" swimtime="00:01:35.93" />
                    <SPLIT distance="150" swimtime="00:02:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="318" reactiontime="+73" swimtime="00:01:26.89" resultid="7783" heatid="11491" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="405" reactiontime="+75" swimtime="00:01:30.76" resultid="7784" heatid="11518" lane="1" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="247" reactiontime="+80" swimtime="00:03:08.14" resultid="7785" heatid="11564" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:19.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="493" reactiontime="+44" swimtime="00:00:38.92" resultid="7786" heatid="11618" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="6738" points="258" reactiontime="+82" swimtime="00:06:48.79" resultid="7787" heatid="11631" lane="6" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:31.83" />
                    <SPLIT distance="150" swimtime="00:02:23.35" />
                    <SPLIT distance="200" swimtime="00:03:15.38" />
                    <SPLIT distance="250" swimtime="00:04:07.93" />
                    <SPLIT distance="300" swimtime="00:05:02.82" />
                    <SPLIT distance="350" swimtime="00:05:57.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Hebel" birthdate="1987-06-22" gender="F" nation="POL" swrid="4754694" athleteid="7767">
              <RESULTS>
                <RESULT eventid="6059" points="463" reactiontime="+98" swimtime="00:00:33.82" resultid="7768" heatid="11398" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="6289" points="469" swimtime="00:01:14.37" resultid="7769" heatid="11464" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" status="DNS" swimtime="00:00:00.00" resultid="7770" heatid="11511" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="6518" points="453" swimtime="00:02:46.80" resultid="7771" heatid="11557" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:19.10" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" status="DNS" swimtime="00:00:00.00" resultid="7772" heatid="11599" lane="5" entrytime="00:03:20.00" />
                <RESULT eventid="6721" points="439" swimtime="00:05:59.20" resultid="7773" heatid="11624" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:02:07.08" />
                    <SPLIT distance="200" swimtime="00:02:53.34" />
                    <SPLIT distance="250" swimtime="00:03:40.06" />
                    <SPLIT distance="300" swimtime="00:04:27.49" />
                    <SPLIT distance="350" swimtime="00:05:13.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dąbrowska" birthdate="1987-05-20" gender="F" nation="POL" swrid="4655165" athleteid="7672">
              <RESULTS>
                <RESULT eventid="6059" points="311" swimtime="00:00:38.61" resultid="7673" heatid="11397" lane="1" entrytime="00:00:39.84" />
                <RESULT eventid="6094" points="256" reactiontime="+115" swimtime="00:03:48.65" resultid="7674" heatid="11421" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                    <SPLIT distance="100" swimtime="00:01:53.02" />
                    <SPLIT distance="150" swimtime="00:02:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="284" swimtime="00:01:27.82" resultid="7675" heatid="11463" lane="9" entrytime="00:01:29.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="233" reactiontime="+102" swimtime="00:01:47.50" resultid="7676" heatid="11480" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="216" reactiontime="+95" swimtime="00:00:47.35" resultid="7677" heatid="11524" lane="5" entrytime="00:00:46.84" />
                <RESULT eventid="6518" points="269" reactiontime="+104" swimtime="00:03:18.36" resultid="7678" heatid="11556" lane="6" entrytime="00:03:22.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="178" reactiontime="+118" swimtime="00:01:53.29" resultid="7679" heatid="11586" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="270" reactiontime="+118" swimtime="00:07:02.31" resultid="7680" heatid="11624" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                    <SPLIT distance="100" swimtime="00:01:39.97" />
                    <SPLIT distance="150" swimtime="00:02:33.89" />
                    <SPLIT distance="200" swimtime="00:03:28.06" />
                    <SPLIT distance="250" swimtime="00:04:23.01" />
                    <SPLIT distance="300" swimtime="00:05:17.27" />
                    <SPLIT distance="350" swimtime="00:06:11.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" swrid="4282341" athleteid="7666">
              <RESULTS>
                <RESULT eventid="6059" points="751" swimtime="00:00:27.82" resultid="7667" heatid="11401" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="6255" points="882" reactiontime="+85" swimtime="00:02:40.21" resultid="7668" heatid="11454" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:01:59.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="767" reactiontime="+82" swimtime="00:01:09.68" resultid="7669" heatid="11486" lane="2" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="824" reactiontime="+80" swimtime="00:01:15.35" resultid="7670" heatid="11512" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="766" reactiontime="+78" swimtime="00:00:34.52" resultid="7671" heatid="11612" lane="5" entrytime="00:00:34.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" swrid="4043251" athleteid="7660">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6077" points="935" reactiontime="+72" swimtime="00:00:24.41" resultid="7661" heatid="11418" lane="9" entrytime="00:00:24.82" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek., Czas lepszy od Rekordu Świata danej kat. wiek." eventid="6238" points="1270" reactiontime="+67" swimtime="00:00:25.73" resultid="7662" heatid="11450" lane="1" entrytime="00:00:26.88" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6467" points="1064" reactiontime="+72" swimtime="00:00:25.15" resultid="7663" heatid="11542" lane="0" entrytime="00:00:25.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6501" points="1088" reactiontime="+66" swimtime="00:00:57.76" resultid="7664" heatid="11553" lane="3" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6636" points="1069" reactiontime="+74" swimtime="00:00:57.26" resultid="7665" heatid="11597" lane="1" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bożena" lastname="Ayomo" birthdate="1966-02-08" gender="F" nation="POL" athleteid="7762">
              <RESULTS>
                <RESULT eventid="6059" points="376" reactiontime="+95" swimtime="00:00:39.79" resultid="7763" heatid="11396" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="6220" points="438" swimtime="00:00:44.56" resultid="7764" heatid="11439" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="6323" points="381" reactiontime="+88" swimtime="00:01:40.53" resultid="7765" heatid="11481" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="412" reactiontime="+96" swimtime="00:00:50.46" resultid="7766" heatid="11608" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" swrid="4992964" athleteid="7687">
              <RESULTS>
                <RESULT eventid="6272" points="742" reactiontime="+70" swimtime="00:02:58.94" resultid="7688" heatid="11458" lane="2" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="150" swimtime="00:02:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="630" reactiontime="+77" swimtime="00:05:54.57" resultid="7689" heatid="11578" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:12.04" />
                    <SPLIT distance="200" swimtime="00:02:56.80" />
                    <SPLIT distance="250" swimtime="00:03:45.31" />
                    <SPLIT distance="300" swimtime="00:04:35.28" />
                    <SPLIT distance="350" swimtime="00:05:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="663" reactiontime="+76" swimtime="00:05:09.25" resultid="7690" heatid="11635" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:01:53.81" />
                    <SPLIT distance="200" swimtime="00:02:33.45" />
                    <SPLIT distance="250" swimtime="00:03:12.48" />
                    <SPLIT distance="300" swimtime="00:03:51.49" />
                    <SPLIT distance="350" swimtime="00:04:30.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" swrid="5312396" athleteid="7710">
              <RESULTS>
                <RESULT eventid="6111" points="513" reactiontime="+82" swimtime="00:02:39.67" resultid="7711" heatid="11431" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="489" reactiontime="+71" swimtime="00:00:34.45" resultid="7712" heatid="11448" lane="5" entrytime="00:00:32.45" />
                <RESULT eventid="6340" points="560" reactiontime="+84" swimtime="00:01:12.55" resultid="7713" heatid="11493" lane="6" entrytime="00:01:12.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="552" reactiontime="+74" swimtime="00:01:11.98" resultid="7714" heatid="11552" lane="1" entrytime="00:01:10.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="443" reactiontime="+89" swimtime="00:05:55.41" resultid="7715" heatid="11578" lane="6" entrytime="00:05:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:05.88" />
                    <SPLIT distance="200" swimtime="00:02:49.47" />
                    <SPLIT distance="250" swimtime="00:03:43.00" />
                    <SPLIT distance="300" swimtime="00:04:35.97" />
                    <SPLIT distance="350" swimtime="00:05:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="588" reactiontime="+71" swimtime="00:02:35.71" resultid="7716" heatid="11605" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7717" heatid="11634" lane="4" entrytime="00:05:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" swrid="4754654" athleteid="7739">
              <RESULTS>
                <RESULT eventid="6077" points="463" reactiontime="+108" swimtime="00:00:34.69" resultid="7740" heatid="11407" lane="4" entrytime="00:00:34.46" />
                <RESULT eventid="6169" points="493" reactiontime="+127" swimtime="00:13:04.43" resultid="7741" heatid="11647" lane="7" entrytime="00:13:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:02:19.40" />
                    <SPLIT distance="200" swimtime="00:03:11.10" />
                    <SPLIT distance="250" swimtime="00:04:02.25" />
                    <SPLIT distance="300" swimtime="00:04:54.36" />
                    <SPLIT distance="350" swimtime="00:05:45.69" />
                    <SPLIT distance="400" swimtime="00:06:37.01" />
                    <SPLIT distance="450" swimtime="00:07:27.81" />
                    <SPLIT distance="500" swimtime="00:08:19.74" />
                    <SPLIT distance="550" swimtime="00:09:08.99" />
                    <SPLIT distance="600" swimtime="00:09:58.16" />
                    <SPLIT distance="650" swimtime="00:10:47.47" />
                    <SPLIT distance="700" swimtime="00:11:35.30" />
                    <SPLIT distance="750" swimtime="00:12:22.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="419" reactiontime="+68" swimtime="00:00:41.95" resultid="7742" heatid="11446" lane="0" entrytime="00:00:42.18" />
                <RESULT eventid="6306" points="474" reactiontime="+114" swimtime="00:01:16.76" resultid="7743" heatid="11471" lane="2" entrytime="00:01:15.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="405" reactiontime="+73" swimtime="00:01:31.31" resultid="7744" heatid="11550" lane="7" entrytime="00:01:33.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="498" reactiontime="+105" swimtime="00:02:52.14" resultid="7745" heatid="11565" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:09.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="517" reactiontime="+67" swimtime="00:03:15.65" resultid="7746" heatid="11603" lane="6" entrytime="00:03:20.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="100" swimtime="00:01:35.95" />
                    <SPLIT distance="150" swimtime="00:02:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="487" reactiontime="+118" swimtime="00:06:09.94" resultid="7747" heatid="11633" lane="9" entrytime="00:06:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="150" swimtime="00:02:16.58" />
                    <SPLIT distance="200" swimtime="00:03:05.41" />
                    <SPLIT distance="250" swimtime="00:03:53.76" />
                    <SPLIT distance="300" swimtime="00:04:41.77" />
                    <SPLIT distance="350" swimtime="00:05:28.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" swrid="5240932" athleteid="7651">
              <RESULTS>
                <RESULT eventid="6059" points="692" reactiontime="+79" swimtime="00:00:29.59" resultid="7652" heatid="11400" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="6094" points="770" reactiontime="+85" swimtime="00:02:38.42" resultid="7653" heatid="11424" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:02:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="845" reactiontime="+71" swimtime="00:00:32.67" resultid="7654" heatid="11441" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="6323" points="761" reactiontime="+81" swimtime="00:01:12.47" resultid="7655" heatid="11486" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="698" reactiontime="+79" swimtime="00:00:32.05" resultid="7656" heatid="11522" lane="4" />
                <RESULT eventid="6484" points="838" reactiontime="+72" swimtime="00:01:09.92" resultid="7657" heatid="11546" lane="3" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6653" points="790" reactiontime="+74" swimtime="00:02:34.42" resultid="7658" heatid="11600" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:01:53.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="576" reactiontime="+80" swimtime="00:00:38.05" resultid="7659" heatid="11612" lane="9" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" swrid="4655152" athleteid="7727">
              <RESULTS>
                <RESULT eventid="6077" points="347" reactiontime="+75" swimtime="00:00:37.03" resultid="7728" heatid="11405" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="6306" points="281" reactiontime="+87" swimtime="00:01:28.57" resultid="7729" heatid="11468" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="286" reactiontime="+90" swimtime="00:01:39.72" resultid="7730" heatid="11489" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="331" reactiontime="+78" swimtime="00:01:38.41" resultid="7731" heatid="11516" lane="6" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="210" swimtime="00:03:32.90" resultid="7732" heatid="11563" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="370" swimtime="00:00:42.48" resultid="7733" heatid="11618" lane="9" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+68" swimtime="00:01:54.98" resultid="9895" heatid="12332" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:02.73" />
                    <SPLIT distance="150" swimtime="00:01:29.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7710" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7696" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="7701" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="7691" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek., Czas lepszy od Rekordu Polski na 1 zmianie," eventid="6610" reactiontime="+74" swimtime="00:01:40.66" resultid="9907" heatid="11584" lane="5" entrytime="00:01:41.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                    <SPLIT distance="100" swimtime="00:00:48.48" />
                    <SPLIT distance="150" swimtime="00:01:16.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7660" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7701" number="2" reactiontime="+115" />
                    <RELAYPOSITION athleteid="7681" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="7696" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+78" swimtime="00:01:59.40" resultid="9908" heatid="11584" lane="0" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:33.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7748" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="7739" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7687" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="7691" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="6">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6779" reactiontime="+64" swimtime="00:01:58.39" resultid="9910" heatid="12331" lane="5" entrytime="00:02:01.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.23" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:29.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7660" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="7681" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="7736" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="7687" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+68" swimtime="00:02:30.92" resultid="9911" heatid="12331" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:01:58.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7739" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7727" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="7748" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="7779" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+98" swimtime="00:02:08.40" resultid="9896" heatid="11581" lane="5" entrytime="00:02:01.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:41.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7762" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="7718" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="7651" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="7788" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6755" reactiontime="+75" swimtime="00:02:08.99" resultid="9897" heatid="11639" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="150" swimtime="00:01:36.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7651" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="7666" number="2" reactiontime="+180" />
                    <RELAYPOSITION athleteid="7788" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="7755" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="6755" reactiontime="+93" swimtime="00:02:46.55" resultid="9906" heatid="11639" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7762" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="7718" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="7672" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7767" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6391" reactiontime="+55" swimtime="00:01:53.08" resultid="9898" heatid="11507" lane="4" entrytime="00:01:55.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.44" />
                    <SPLIT distance="100" swimtime="00:01:01.26" />
                    <SPLIT distance="150" swimtime="00:01:26.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7734" number="1" reactiontime="+55" />
                    <RELAYPOSITION athleteid="7666" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="7660" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="7788" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6128" reactiontime="+79" swimtime="00:01:42.20" resultid="9899" heatid="11436" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:00:51.76" />
                    <SPLIT distance="150" swimtime="00:01:18.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7666" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="7701" number="2" reactiontime="+181" />
                    <RELAYPOSITION athleteid="7788" number="3" reactiontime="+122" />
                    <RELAYPOSITION athleteid="7696" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+82" swimtime="00:02:14.11" resultid="9900" heatid="11507" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:39.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7762" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="7696" number="2" reactiontime="+9" />
                    <RELAYPOSITION athleteid="7701" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="7767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6128" swimtime="00:02:08.80" resultid="9901" heatid="11436" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:39.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7779" number="1" />
                    <RELAYPOSITION athleteid="7767" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="7755" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="7748" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+77" swimtime="00:01:58.65" resultid="9902" heatid="11436" lane="2" entrytime="00:01:58.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:30.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7718" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="7687" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="7651" number="3" reactiontime="+183" />
                    <RELAYPOSITION athleteid="7681" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6391" reactiontime="+74" swimtime="00:02:09.72" resultid="9903" heatid="11507" lane="7" entrytime="00:02:13.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:10.41" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7651" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7718" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="7681" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="7687" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+92" swimtime="00:02:30.05" resultid="9904" heatid="11435" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:55.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7762" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="7727" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="7672" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="7739" number="4" reactiontime="+79" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+67" swimtime="00:02:30.07" resultid="9905" heatid="11507" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:57.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7710" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7779" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="7672" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7755" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01813" nation="POL" region="13" clubid="9448" name="SWIMLAND Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Wójtowicz" birthdate="1995-02-20" gender="F" nation="POL" license="101813600026" swrid="4265548" athleteid="9449">
              <RESULTS>
                <RESULT eventid="6059" points="865" reactiontime="+61" swimtime="00:00:26.54" resultid="9450" heatid="11401" lane="4" entrytime="00:00:26.30" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6220" points="1119" reactiontime="+63" swimtime="00:00:28.45" resultid="9451" heatid="11441" lane="4" entrytime="00:00:28.72" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6484" points="1129" reactiontime="+66" swimtime="00:01:01.23" resultid="9452" heatid="11546" lane="4" entrytime="00:01:00.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" status="DNS" swimtime="00:00:00.00" resultid="9453" heatid="11600" lane="4" entrytime="00:02:19.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7202" name="Kościańskie Towarzystwo Pływackie">
          <ATHLETES>
            <ATHLETE firstname="Mariusz" lastname="Wesołowski" birthdate="1981-01-01" gender="M" nation="POL" athleteid="7226">
              <RESULTS>
                <RESULT eventid="6340" points="232" reactiontime="+88" swimtime="00:01:37.24" resultid="7227" heatid="11489" lane="1" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="187" reactiontime="+96" swimtime="00:00:43.94" resultid="7228" heatid="11532" lane="7" entrytime="00:00:46.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Naglik" birthdate="1968-01-01" gender="M" nation="POL" athleteid="7214">
              <RESULTS>
                <RESULT eventid="6374" points="203" reactiontime="+97" swimtime="00:03:56.07" resultid="7215" heatid="11501" lane="5" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.37" />
                    <SPLIT distance="100" swimtime="00:01:48.36" />
                    <SPLIT distance="150" swimtime="00:02:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="7216" heatid="11576" lane="3" entrytime="00:08:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Pelec" birthdate="1987-01-01" gender="M" nation="POL" athleteid="7229">
              <RESULTS>
                <RESULT eventid="6306" points="236" swimtime="00:01:19.85" resultid="7230" heatid="11468" lane="7" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="195" swimtime="00:01:49.49" resultid="7231" heatid="11515" lane="6" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="167" swimtime="00:00:42.90" resultid="7232" heatid="11533" lane="3" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Szmyt" birthdate="1962-01-01" gender="M" nation="POL" athleteid="7217">
              <RESULTS>
                <RESULT eventid="6203" points="322" swimtime="00:28:34.60" resultid="7218" heatid="11653" lane="7" entrytime="00:26:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:40.70" />
                    <SPLIT distance="150" swimtime="00:02:34.38" />
                    <SPLIT distance="200" swimtime="00:03:30.67" />
                    <SPLIT distance="250" swimtime="00:04:29.94" />
                    <SPLIT distance="300" swimtime="00:05:29.58" />
                    <SPLIT distance="350" swimtime="00:06:28.35" />
                    <SPLIT distance="400" swimtime="00:07:27.70" />
                    <SPLIT distance="450" swimtime="00:08:26.24" />
                    <SPLIT distance="500" swimtime="00:09:25.84" />
                    <SPLIT distance="550" swimtime="00:10:24.22" />
                    <SPLIT distance="600" swimtime="00:11:22.47" />
                    <SPLIT distance="650" swimtime="00:12:21.53" />
                    <SPLIT distance="700" swimtime="00:13:19.61" />
                    <SPLIT distance="750" swimtime="00:14:17.73" />
                    <SPLIT distance="800" swimtime="00:15:15.78" />
                    <SPLIT distance="850" swimtime="00:16:12.23" />
                    <SPLIT distance="900" swimtime="00:17:08.94" />
                    <SPLIT distance="950" swimtime="00:18:05.62" />
                    <SPLIT distance="1000" swimtime="00:19:02.34" />
                    <SPLIT distance="1050" swimtime="00:19:58.64" />
                    <SPLIT distance="1100" swimtime="00:20:55.50" />
                    <SPLIT distance="1150" swimtime="00:21:51.99" />
                    <SPLIT distance="1200" swimtime="00:22:49.24" />
                    <SPLIT distance="1250" swimtime="00:23:46.94" />
                    <SPLIT distance="1300" swimtime="00:24:45.15" />
                    <SPLIT distance="1350" swimtime="00:25:43.11" />
                    <SPLIT distance="1400" swimtime="00:26:41.47" />
                    <SPLIT distance="1450" swimtime="00:27:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="7219" heatid="11602" lane="2" entrytime="00:04:15.00" entrycourse="SCM" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7220" heatid="11631" lane="4" entrytime="00:06:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Brygier" birthdate="1979-01-01" gender="F" nation="POL" athleteid="7203">
              <RESULTS>
                <RESULT eventid="6357" status="DNF" swimtime="00:00:00.00" resultid="7204" heatid="11499" lane="9" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" status="DNS" swimtime="00:00:00.00" resultid="7205" heatid="11573" lane="1" entrytime="00:08:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Skrzypczak" birthdate="1966-01-01" gender="M" nation="POL" swrid="4992721" athleteid="7209">
              <RESULTS>
                <RESULT eventid="6077" points="473" reactiontime="+81" swimtime="00:00:33.39" resultid="7210" heatid="11408" lane="0" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="6111" points="322" reactiontime="+90" swimtime="00:03:26.90" resultid="7211" heatid="11427" lane="4" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:01:34.88" />
                    <SPLIT distance="150" swimtime="00:02:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="313" reactiontime="+81" swimtime="00:03:24.74" resultid="7212" heatid="11502" lane="0" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="7213" heatid="11577" lane="8" entrytime="00:07:35.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Morawski" birthdate="1991-02-22" gender="M" nation="POL" athleteid="7233">
              <RESULTS>
                <RESULT eventid="6077" points="339" reactiontime="+87" swimtime="00:00:31.73" resultid="7234" heatid="11407" lane="6" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="6169" reactiontime="+92" status="OTL" swimtime="00:00:00.00" resultid="7235" heatid="11646" lane="5" entrytime="00:10:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:01:27.90" />
                    <SPLIT distance="150" swimtime="00:02:20.28" />
                    <SPLIT distance="200" swimtime="00:03:16.33" />
                    <SPLIT distance="250" swimtime="00:04:13.09" />
                    <SPLIT distance="300" swimtime="00:05:11.77" />
                    <SPLIT distance="350" swimtime="00:06:11.48" />
                    <SPLIT distance="400" swimtime="00:08:10.43" />
                    <SPLIT distance="450" swimtime="00:09:10.58" />
                    <SPLIT distance="500" swimtime="00:10:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="283" reactiontime="+93" swimtime="00:03:33.91" resultid="7236" heatid="11456" lane="1" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                    <SPLIT distance="100" swimtime="00:01:42.27" />
                    <SPLIT distance="150" swimtime="00:02:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="231" reactiontime="+97" swimtime="00:01:29.58" resultid="7237" heatid="11489" lane="0" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="267" reactiontime="+93" swimtime="00:01:35.23" resultid="7238" heatid="11515" lane="3" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="172" reactiontime="+98" swimtime="00:03:11.25" resultid="7239" heatid="11564" lane="7" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:19.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7240" heatid="11618" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7241" heatid="11636" lane="0" entrytime="00:05:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewelina" lastname="Braun" birthdate="1976-01-01" gender="F" nation="POL" athleteid="7206">
              <RESULTS>
                <RESULT eventid="6255" points="287" reactiontime="+119" swimtime="00:04:16.35" resultid="7207" heatid="11452" lane="7" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.36" />
                    <SPLIT distance="100" swimtime="00:02:04.89" />
                    <SPLIT distance="150" swimtime="00:03:11.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="291" reactiontime="+94" swimtime="00:01:56.94" resultid="7208" heatid="11510" lane="5" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Kunc" birthdate="1961-01-01" gender="M" nation="POL" athleteid="7242">
              <RESULTS>
                <RESULT eventid="6306" points="175" reactiontime="+157" swimtime="00:01:46.90" resultid="7243" heatid="11468" lane="0" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="150" reactiontime="+153" swimtime="00:00:54.85" resultid="7244" heatid="11532" lane="9" entrytime="00:00:54.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Mulczyński" birthdate="1976-01-01" gender="M" nation="POL" athleteid="7221">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7222" heatid="11409" lane="9" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="6203" points="251" reactiontime="+87" swimtime="00:26:06.60" resultid="7223" heatid="11653" lane="3" entrytime="00:24:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:24.48" />
                    <SPLIT distance="150" swimtime="00:02:12.30" />
                    <SPLIT distance="200" swimtime="00:03:01.67" />
                    <SPLIT distance="250" swimtime="00:03:52.40" />
                    <SPLIT distance="300" swimtime="00:04:43.70" />
                    <SPLIT distance="350" swimtime="00:05:35.82" />
                    <SPLIT distance="400" swimtime="00:06:28.26" />
                    <SPLIT distance="450" swimtime="00:07:20.68" />
                    <SPLIT distance="500" swimtime="00:08:13.88" />
                    <SPLIT distance="550" swimtime="00:09:06.65" />
                    <SPLIT distance="600" swimtime="00:09:59.98" />
                    <SPLIT distance="650" swimtime="00:10:53.17" />
                    <SPLIT distance="700" swimtime="00:11:46.59" />
                    <SPLIT distance="750" swimtime="00:12:39.93" />
                    <SPLIT distance="800" swimtime="00:13:33.58" />
                    <SPLIT distance="850" swimtime="00:14:27.19" />
                    <SPLIT distance="900" swimtime="00:15:19.88" />
                    <SPLIT distance="950" swimtime="00:16:12.69" />
                    <SPLIT distance="1000" swimtime="00:17:06.82" />
                    <SPLIT distance="1050" swimtime="00:18:01.72" />
                    <SPLIT distance="1100" swimtime="00:18:55.41" />
                    <SPLIT distance="1150" swimtime="00:19:49.94" />
                    <SPLIT distance="1200" swimtime="00:20:43.97" />
                    <SPLIT distance="1250" swimtime="00:21:38.73" />
                    <SPLIT distance="1300" swimtime="00:22:33.53" />
                    <SPLIT distance="1350" swimtime="00:23:27.82" />
                    <SPLIT distance="1400" swimtime="00:24:21.03" />
                    <SPLIT distance="1450" swimtime="00:25:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="297" reactiontime="+68" swimtime="00:00:38.45" resultid="7224" heatid="11532" lane="3" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7225" heatid="11633" lane="2" entrytime="00:05:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" status="DNS" swimtime="00:00:00.00" resultid="7245" heatid="11583" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7229" number="1" />
                    <RELAYPOSITION athleteid="7233" number="2" />
                    <RELAYPOSITION athleteid="7214" number="3" />
                    <RELAYPOSITION athleteid="7226" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+86" swimtime="00:03:05.39" resultid="7246" heatid="11505" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                    <SPLIT distance="100" swimtime="00:01:38.15" />
                    <SPLIT distance="150" swimtime="00:02:06.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7209" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="7206" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="7214" number="3" />
                    <RELAYPOSITION athleteid="7203" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA 191" nation="POL" clubid="8007" name="Korona 1919 Kraków">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Mleczko" birthdate="1947-08-26" gender="M" nation="POL" swrid="4992812" athleteid="8029">
              <RESULTS>
                <RESULT eventid="6077" points="557" reactiontime="+117" swimtime="00:00:38.04" resultid="8030" heatid="11405" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="6169" points="402" reactiontime="+139" swimtime="00:16:27.40" resultid="8031" heatid="11648" lane="4" entrytime="00:14:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                    <SPLIT distance="100" swimtime="00:01:54.16" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                    <SPLIT distance="200" swimtime="00:03:56.70" />
                    <SPLIT distance="250" swimtime="00:04:58.31" />
                    <SPLIT distance="300" swimtime="00:06:00.25" />
                    <SPLIT distance="350" swimtime="00:07:02.49" />
                    <SPLIT distance="400" swimtime="00:08:04.12" />
                    <SPLIT distance="450" swimtime="00:09:06.58" />
                    <SPLIT distance="500" swimtime="00:10:09.01" />
                    <SPLIT distance="550" swimtime="00:11:12.00" />
                    <SPLIT distance="600" swimtime="00:12:14.56" />
                    <SPLIT distance="650" swimtime="00:13:18.82" />
                    <SPLIT distance="700" swimtime="00:14:23.27" />
                    <SPLIT distance="750" swimtime="00:15:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="522" reactiontime="+123" swimtime="00:01:28.33" resultid="8032" heatid="11469" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="344" reactiontime="+130" swimtime="00:01:59.10" resultid="8033" heatid="11489" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="324" reactiontime="+127" swimtime="00:03:51.22" resultid="8034" heatid="11563" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.75" />
                    <SPLIT distance="100" swimtime="00:01:51.72" />
                    <SPLIT distance="150" swimtime="00:02:51.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="288" reactiontime="+140" swimtime="00:10:24.66" resultid="8035" heatid="11576" lane="2" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.20" />
                    <SPLIT distance="100" swimtime="00:02:37.13" />
                    <SPLIT distance="150" swimtime="00:04:01.95" />
                    <SPLIT distance="200" swimtime="00:05:25.10" />
                    <SPLIT distance="250" swimtime="00:06:51.61" />
                    <SPLIT distance="300" swimtime="00:08:17.49" />
                    <SPLIT distance="350" swimtime="00:09:22.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="234" reactiontime="+134" swimtime="00:02:17.91" resultid="8036" heatid="11590" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="362" reactiontime="+141" swimtime="00:08:11.74" resultid="8037" heatid="11631" lane="7" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.02" />
                    <SPLIT distance="100" swimtime="00:01:58.12" />
                    <SPLIT distance="150" swimtime="00:03:01.91" />
                    <SPLIT distance="200" swimtime="00:04:05.68" />
                    <SPLIT distance="250" swimtime="00:05:09.32" />
                    <SPLIT distance="300" swimtime="00:06:12.17" />
                    <SPLIT distance="350" swimtime="00:07:14.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" swrid="4218717" athleteid="8056">
              <RESULTS>
                <RESULT eventid="6323" points="354" swimtime="00:01:37.58" resultid="8057" heatid="11482" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="622" reactiontime="+95" swimtime="00:00:36.49" resultid="8058" heatid="11524" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="6484" points="312" reactiontime="+95" swimtime="00:01:38.92" resultid="8059" heatid="11545" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="258" swimtime="00:01:46.20" resultid="8060" heatid="11586" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="363" reactiontime="+107" swimtime="00:03:25.81" resultid="8061" heatid="11599" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:43.89" />
                    <SPLIT distance="150" swimtime="00:02:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Łysiak" birthdate="1973-03-30" gender="M" nation="POL" swrid="5468085" athleteid="8016">
              <RESULTS>
                <RESULT eventid="6111" points="461" reactiontime="+94" swimtime="00:02:51.35" resultid="8017" heatid="11430" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:22.10" />
                    <SPLIT distance="150" swimtime="00:02:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="538" reactiontime="+97" swimtime="00:03:01.49" resultid="8018" heatid="11459" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:27.23" />
                    <SPLIT distance="150" swimtime="00:02:13.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="500" reactiontime="+86" swimtime="00:01:23.18" resultid="8019" heatid="11519" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8020" heatid="11604" lane="2" entrytime="00:02:55.00" />
                <RESULT eventid="6704" points="443" reactiontime="+88" swimtime="00:00:39.73" resultid="8021" heatid="11620" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Jawień" birthdate="1971-06-11" gender="M" nation="POL" swrid="5468083" athleteid="8101">
              <RESULTS>
                <RESULT eventid="6111" points="524" reactiontime="+77" swimtime="00:02:43.60" resultid="8102" heatid="11430" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:17.04" />
                    <SPLIT distance="150" swimtime="00:02:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="519" reactiontime="+79" swimtime="00:00:35.29" resultid="8103" heatid="11444" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="6272" points="644" swimtime="00:02:59.18" resultid="8104" heatid="11459" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="585" reactiontime="+79" swimtime="00:01:20.27" resultid="8105" heatid="11515" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="514" reactiontime="+77" swimtime="00:01:15.47" resultid="8106" heatid="11551" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="521" reactiontime="+81" swimtime="00:01:14.15" resultid="8107" heatid="11590" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="575" reactiontime="+81" swimtime="00:02:47.31" resultid="8108" heatid="11604" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="150" swimtime="00:02:06.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" swrid="4992907" athleteid="8083">
              <RESULTS>
                <RESULT eventid="6059" status="DNS" swimtime="00:00:00.00" resultid="8084" heatid="11400" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="6094" status="DNS" swimtime="00:00:00.00" resultid="8085" heatid="11423" lane="6" entrytime="00:02:53.00" />
                <RESULT eventid="6220" points="604" reactiontime="+73" swimtime="00:00:36.13" resultid="8086" heatid="11441" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="6323" points="686" reactiontime="+86" swimtime="00:01:17.25" resultid="8087" heatid="11485" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="672" reactiontime="+81" swimtime="00:00:33.45" resultid="8088" heatid="11526" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="6484" points="611" reactiontime="+71" swimtime="00:01:20.08" resultid="8089" heatid="11545" lane="4" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="647" reactiontime="+69" swimtime="00:02:52.73" resultid="8090" heatid="11600" lane="1" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                    <SPLIT distance="150" swimtime="00:02:09.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="585" reactiontime="+84" swimtime="00:00:41.05" resultid="8091" heatid="11611" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska" birthdate="1984-04-20" gender="F" nation="POL" swrid="5468078" athleteid="8077">
              <RESULTS>
                <RESULT eventid="6059" status="DNS" swimtime="00:00:00.00" resultid="8078" heatid="11396" lane="7" entrytime="00:00:49.00" />
                <RESULT eventid="6220" status="DNS" swimtime="00:00:00.00" resultid="8079" heatid="11439" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="6255" status="DNS" swimtime="00:00:00.00" resultid="8080" heatid="11452" lane="2" entrytime="00:04:15.00" />
                <RESULT eventid="6415" status="DNS" swimtime="00:00:00.00" resultid="8081" heatid="11510" lane="6" entrytime="00:01:58.00" />
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="8082" heatid="11610" lane="0" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" swrid="4992740" athleteid="8062">
              <RESULTS>
                <RESULT eventid="6077" points="815" reactiontime="+75" swimtime="00:00:26.21" resultid="8063" heatid="11415" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="6306" points="707" swimtime="00:00:59.59" resultid="8064" heatid="11475" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="593" reactiontime="+75" swimtime="00:01:10.60" resultid="8065" heatid="11495" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="799" reactiontime="+79" swimtime="00:00:28.89" resultid="8066" heatid="11539" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="6636" points="598" reactiontime="+77" swimtime="00:01:10.82" resultid="8067" heatid="11594" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="749" reactiontime="+78" swimtime="00:00:33.86" resultid="8068" heatid="11621" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Orlewicz-Musiał" birthdate="1960-05-29" gender="F" nation="POL" swrid="5352178" athleteid="8092">
              <RESULTS>
                <RESULT eventid="6094" points="248" swimtime="00:04:37.35" resultid="8093" heatid="11420" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.04" />
                    <SPLIT distance="100" swimtime="00:02:11.43" />
                    <SPLIT distance="150" swimtime="00:03:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="268" reactiontime="+107" swimtime="00:33:25.79" resultid="8094" heatid="11651" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:57.46" />
                    <SPLIT distance="150" swimtime="00:03:04.92" />
                    <SPLIT distance="200" swimtime="00:04:11.45" />
                    <SPLIT distance="250" swimtime="00:05:17.85" />
                    <SPLIT distance="300" swimtime="00:06:24.54" />
                    <SPLIT distance="350" swimtime="00:07:31.55" />
                    <SPLIT distance="400" swimtime="00:08:40.11" />
                    <SPLIT distance="450" swimtime="00:09:46.61" />
                    <SPLIT distance="500" swimtime="00:10:54.86" />
                    <SPLIT distance="550" swimtime="00:12:01.67" />
                    <SPLIT distance="600" swimtime="00:13:09.23" />
                    <SPLIT distance="650" swimtime="00:14:15.99" />
                    <SPLIT distance="700" swimtime="00:15:23.75" />
                    <SPLIT distance="750" swimtime="00:16:29.80" />
                    <SPLIT distance="800" swimtime="00:17:35.97" />
                    <SPLIT distance="850" swimtime="00:18:43.40" />
                    <SPLIT distance="900" swimtime="00:19:51.25" />
                    <SPLIT distance="950" swimtime="00:20:58.05" />
                    <SPLIT distance="1000" swimtime="00:22:05.67" />
                    <SPLIT distance="1050" swimtime="00:23:13.82" />
                    <SPLIT distance="1100" swimtime="00:24:20.36" />
                    <SPLIT distance="1150" swimtime="00:25:29.25" />
                    <SPLIT distance="1200" swimtime="00:26:36.93" />
                    <SPLIT distance="1250" swimtime="00:27:45.56" />
                    <SPLIT distance="1300" swimtime="00:28:52.42" />
                    <SPLIT distance="1350" swimtime="00:30:01.51" />
                    <SPLIT distance="1400" swimtime="00:31:09.36" />
                    <SPLIT distance="1450" swimtime="00:32:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="191" reactiontime="+47" swimtime="00:01:03.05" resultid="8095" heatid="11437" lane="3" />
                <RESULT eventid="6357" points="230" reactiontime="+105" swimtime="00:05:31.50" resultid="8096" heatid="11498" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.99" />
                    <SPLIT distance="100" swimtime="00:02:29.36" />
                    <SPLIT distance="150" swimtime="00:04:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" status="DNS" swimtime="00:00:00.00" resultid="8097" heatid="11544" lane="1" />
                <RESULT eventid="6552" points="261" reactiontime="+95" swimtime="00:09:56.65" resultid="8098" heatid="11572" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.37" />
                    <SPLIT distance="100" swimtime="00:02:27.12" />
                    <SPLIT distance="150" swimtime="00:03:44.36" />
                    <SPLIT distance="200" swimtime="00:05:00.49" />
                    <SPLIT distance="250" swimtime="00:06:24.24" />
                    <SPLIT distance="300" swimtime="00:07:48.21" />
                    <SPLIT distance="350" swimtime="00:08:52.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="172" reactiontime="+92" swimtime="00:02:26.22" resultid="8099" heatid="11585" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="200" reactiontime="+102" swimtime="00:08:58.97" resultid="8100" heatid="11624" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.84" />
                    <SPLIT distance="100" swimtime="00:02:03.03" />
                    <SPLIT distance="150" swimtime="00:03:11.48" />
                    <SPLIT distance="200" swimtime="00:04:21.38" />
                    <SPLIT distance="250" swimtime="00:05:30.97" />
                    <SPLIT distance="300" swimtime="00:06:38.73" />
                    <SPLIT distance="350" swimtime="00:07:47.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-03-21" gender="M" nation="POL" swrid="4992712" athleteid="8038">
              <RESULTS>
                <RESULT eventid="6077" points="594" reactiontime="+93" swimtime="00:00:30.96" resultid="8039" heatid="11410" lane="5" entrytime="00:00:30.76" />
                <RESULT eventid="6111" points="482" reactiontime="+86" swimtime="00:03:00.98" resultid="8040" heatid="11429" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="150" swimtime="00:02:20.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="552" reactiontime="+99" swimtime="00:03:17.51" resultid="8041" heatid="11457" lane="5" entrytime="00:03:17.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:32.13" />
                    <SPLIT distance="150" swimtime="00:02:24.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="505" reactiontime="+98" swimtime="00:01:22.51" resultid="8042" heatid="11491" lane="6" entrytime="00:01:21.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="457" reactiontime="+98" swimtime="00:01:28.42" resultid="8043" heatid="11514" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="434" swimtime="00:00:37.04" resultid="8044" heatid="11533" lane="4" entrytime="00:00:38.42" />
                <RESULT eventid="6670" points="437" reactiontime="+92" swimtime="00:03:08.66" resultid="8045" heatid="11601" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:34.11" />
                    <SPLIT distance="150" swimtime="00:02:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="470" reactiontime="+93" swimtime="00:00:39.22" resultid="8046" heatid="11618" lane="2" entrytime="00:00:39.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mucha" birthdate="1967-04-24" gender="M" nation="POL" swrid="4218718" athleteid="8113">
              <RESULTS>
                <RESULT eventid="6433" points="461" reactiontime="+89" swimtime="00:01:28.18" resultid="8114" heatid="11518" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="501" reactiontime="+84" swimtime="00:00:38.39" resultid="8115" heatid="11619" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" swrid="5484421" athleteid="8022">
              <RESULTS>
                <RESULT eventid="6272" points="432" reactiontime="+101" swimtime="00:03:39.38" resultid="8023" heatid="11456" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:47.09" />
                    <SPLIT distance="150" swimtime="00:02:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="276" reactiontime="+94" swimtime="00:04:05.10" resultid="8024" heatid="11501" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                    <SPLIT distance="100" swimtime="00:01:56.37" />
                    <SPLIT distance="150" swimtime="00:03:01.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="338" reactiontime="+81" swimtime="00:01:46.02" resultid="8025" heatid="11515" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="228" swimtime="00:00:47.66" resultid="8026" heatid="11531" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="6636" points="231" reactiontime="+87" swimtime="00:01:49.75" resultid="8027" heatid="11590" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="329" reactiontime="+99" swimtime="00:00:47.40" resultid="8028" heatid="11615" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" swrid="4992827" athleteid="8047">
              <RESULTS>
                <RESULT eventid="6059" points="704" swimtime="00:00:34.85" resultid="8048" heatid="11398" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="6145" points="739" swimtime="00:12:45.36" resultid="8049" heatid="11643" lane="8" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:02:12.72" />
                    <SPLIT distance="200" swimtime="00:03:01.01" />
                    <SPLIT distance="250" swimtime="00:03:49.60" />
                    <SPLIT distance="300" swimtime="00:04:37.97" />
                    <SPLIT distance="350" swimtime="00:05:26.69" />
                    <SPLIT distance="400" swimtime="00:06:15.54" />
                    <SPLIT distance="450" swimtime="00:07:04.50" />
                    <SPLIT distance="500" swimtime="00:07:54.00" />
                    <SPLIT distance="550" swimtime="00:08:42.99" />
                    <SPLIT distance="600" swimtime="00:09:32.15" />
                    <SPLIT distance="650" swimtime="00:10:21.02" />
                    <SPLIT distance="700" swimtime="00:11:09.99" />
                    <SPLIT distance="750" swimtime="00:11:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="644" swimtime="00:01:18.89" resultid="8050" heatid="11464" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="915" swimtime="00:03:29.30" resultid="8051" heatid="11499" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                    <SPLIT distance="100" swimtime="00:01:37.24" />
                    <SPLIT distance="150" swimtime="00:02:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="8052" heatid="11525" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="6518" points="624" swimtime="00:02:51.66" resultid="8053" heatid="11557" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                    <SPLIT distance="150" swimtime="00:02:07.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="663" swimtime="00:01:33.39" resultid="8054" heatid="11587" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="615" swimtime="00:06:10.99" resultid="8055" heatid="11627" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:26.11" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                    <SPLIT distance="200" swimtime="00:03:00.38" />
                    <SPLIT distance="250" swimtime="00:03:48.30" />
                    <SPLIT distance="300" swimtime="00:04:36.51" />
                    <SPLIT distance="350" swimtime="00:05:24.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisłąw" lastname="Waga" birthdate="1940-07-04" gender="M" nation="POL" swrid="4992823" athleteid="8069">
              <RESULTS>
                <RESULT eventid="6077" points="267" reactiontime="+110" swimtime="00:00:49.78" resultid="8070" heatid="11404" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="6169" points="315" reactiontime="+105" swimtime="00:18:52.34" resultid="8071" heatid="11648" lane="8" entrytime="00:17:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.81" />
                    <SPLIT distance="100" swimtime="00:02:17.94" />
                    <SPLIT distance="150" swimtime="00:03:31.61" />
                    <SPLIT distance="200" swimtime="00:04:44.11" />
                    <SPLIT distance="250" swimtime="00:05:54.68" />
                    <SPLIT distance="300" swimtime="00:07:06.46" />
                    <SPLIT distance="350" swimtime="00:08:18.73" />
                    <SPLIT distance="400" swimtime="00:09:30.55" />
                    <SPLIT distance="450" swimtime="00:10:42.35" />
                    <SPLIT distance="500" swimtime="00:11:53.50" />
                    <SPLIT distance="550" swimtime="00:13:05.40" />
                    <SPLIT distance="600" swimtime="00:14:16.51" />
                    <SPLIT distance="650" swimtime="00:15:26.38" />
                    <SPLIT distance="700" swimtime="00:16:38.13" />
                    <SPLIT distance="750" swimtime="00:17:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="270" swimtime="00:01:53.97" resultid="8072" heatid="11467" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="169" reactiontime="+108" swimtime="00:02:55.21" resultid="8073" heatid="11514" lane="4" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="244" reactiontime="+116" swimtime="00:04:26.48" resultid="8074" heatid="11562" lane="5" entrytime="00:04:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.35" />
                    <SPLIT distance="100" swimtime="00:02:11.68" />
                    <SPLIT distance="150" swimtime="00:03:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="205" reactiontime="+105" swimtime="00:01:12.89" resultid="8075" heatid="11615" lane="2" entrytime="00:01:13.00" />
                <RESULT eventid="6738" points="268" reactiontime="+116" swimtime="00:09:18.27" resultid="8076" heatid="11630" lane="6" entrytime="00:09:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.17" />
                    <SPLIT distance="100" swimtime="00:02:18.28" />
                    <SPLIT distance="150" swimtime="00:03:31.08" />
                    <SPLIT distance="200" swimtime="00:04:43.15" />
                    <SPLIT distance="250" swimtime="00:05:53.77" />
                    <SPLIT distance="300" swimtime="00:07:04.36" />
                    <SPLIT distance="350" swimtime="00:08:14.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Pyczek" birthdate="1991-07-20" gender="F" nation="POL" athleteid="8109">
              <RESULTS>
                <RESULT eventid="6450" points="509" reactiontime="+69" swimtime="00:00:35.30" resultid="8110" heatid="11526" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="6518" points="498" reactiontime="+74" swimtime="00:02:38.49" resultid="8111" heatid="11558" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="449" swimtime="00:05:51.85" resultid="8112" heatid="11627" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                    <SPLIT distance="200" swimtime="00:02:48.06" />
                    <SPLIT distance="250" swimtime="00:03:33.28" />
                    <SPLIT distance="300" swimtime="00:04:19.53" />
                    <SPLIT distance="350" swimtime="00:05:06.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" swrid="4992797" athleteid="8008">
              <RESULTS>
                <RESULT eventid="6059" points="814" reactiontime="+75" swimtime="00:00:30.77" resultid="8009" heatid="11399" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="6220" points="786" reactiontime="+69" swimtime="00:00:36.67" resultid="8010" heatid="11440" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="6323" points="803" reactiontime="+80" swimtime="00:01:18.45" resultid="8011" heatid="11485" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6415" points="842" reactiontime="+81" swimtime="00:01:28.13" resultid="8012" heatid="11511" lane="4" entrytime="00:01:29.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="744" reactiontime="+72" swimtime="00:01:22.10" resultid="8013" heatid="11546" lane="9" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" status="DNS" swimtime="00:00:00.00" resultid="8014" heatid="11600" lane="9" entrytime="00:03:02.00" />
                <RESULT eventid="6687" points="930" swimtime="00:00:38.48" resultid="8015" heatid="11611" lane="4" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona 1919 Kroaków" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+91" swimtime="00:02:17.09" resultid="9829" heatid="11583" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:00:57.39" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8016" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="8062" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="8022" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="8029" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona 1919 Kroaków" number="1">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+80" swimtime="00:02:13.00" resultid="9830" heatid="11581" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:41.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8008" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="8056" number="2" />
                    <RELAYPOSITION athleteid="8047" number="3" />
                    <RELAYPOSITION athleteid="8083" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona 1919 Kroaków" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6128" reactiontime="+74" swimtime="00:01:58.04" resultid="9826" heatid="11436" lane="6" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:31.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8008" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="8101" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="8083" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="8062" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+70" swimtime="00:02:12.72" resultid="9827" heatid="11507" lane="1" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:01:46.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8083" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="8101" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="8008" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="8062" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona 1919 Kroaków 2" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+89" swimtime="00:02:36.63" resultid="9828" heatid="11506" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8047" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="8113" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="8056" number="3" reactiontime="+83" />
                    <RELAYPOSITION athleteid="8029" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6918" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Zdzisława" lastname="Wiese" birthdate="1952-01-01" gender="F" nation="POL" athleteid="6917">
              <RESULTS>
                <RESULT eventid="6255" points="298" reactiontime="+158" swimtime="00:05:19.19" resultid="6919" heatid="11452" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.53" />
                    <SPLIT distance="100" swimtime="00:02:31.21" />
                    <SPLIT distance="150" swimtime="00:03:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="271" reactiontime="+101" swimtime="00:02:30.04" resultid="6920" heatid="11509" lane="5" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="286" reactiontime="+101" swimtime="00:01:05.48" resultid="6921" heatid="11609" lane="0" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" clubid="7565" name="Landsberg Crew Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Kaczmarek" birthdate="1992-08-23" gender="F" nation="POL" license="501304600002" athleteid="7575">
              <RESULTS>
                <RESULT eventid="6059" points="708" swimtime="00:00:29.05" resultid="7576" heatid="11401" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="6094" points="796" reactiontime="+74" swimtime="00:02:34.19" resultid="7577" heatid="11424" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:13.63" />
                    <SPLIT distance="150" swimtime="00:01:58.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="763" reactiontime="+75" swimtime="00:01:02.87" resultid="7578" heatid="11466" lane="2" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="756" reactiontime="+77" swimtime="00:01:11.15" resultid="7579" heatid="11486" lane="7" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="651" reactiontime="+75" swimtime="00:01:19.90" resultid="7580" heatid="11512" lane="5" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6552" points="763" reactiontime="+81" swimtime="00:05:26.76" resultid="7581" heatid="11574" lane="5" entrytime="00:05:32.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:57.14" />
                    <SPLIT distance="200" swimtime="00:02:39.32" />
                    <SPLIT distance="250" swimtime="00:03:24.73" />
                    <SPLIT distance="300" swimtime="00:04:12.07" />
                    <SPLIT distance="350" swimtime="00:04:49.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="662" reactiontime="+75" swimtime="00:00:35.96" resultid="7582" heatid="11612" lane="7" entrytime="00:00:36.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6721" points="762" reactiontime="+82" swimtime="00:04:54.97" resultid="7583" heatid="11628" lane="3" entrytime="00:04:56.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:49.38" />
                    <SPLIT distance="200" swimtime="00:02:26.94" />
                    <SPLIT distance="250" swimtime="00:03:04.60" />
                    <SPLIT distance="300" swimtime="00:03:42.13" />
                    <SPLIT distance="350" swimtime="00:04:19.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" license="501304700001" swrid="4432188" athleteid="7566">
              <RESULTS>
                <RESULT eventid="6111" points="691" reactiontime="+77" swimtime="00:02:24.60" resultid="7567" heatid="11433" lane="6" entrytime="00:02:19.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" points="707" reactiontime="+74" swimtime="00:09:34.32" resultid="7568" heatid="11645" lane="4" entrytime="00:09:10.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:44.76" />
                    <SPLIT distance="200" swimtime="00:02:20.81" />
                    <SPLIT distance="250" swimtime="00:02:57.11" />
                    <SPLIT distance="300" swimtime="00:03:33.35" />
                    <SPLIT distance="350" swimtime="00:04:09.61" />
                    <SPLIT distance="400" swimtime="00:04:46.20" />
                    <SPLIT distance="450" swimtime="00:05:22.68" />
                    <SPLIT distance="500" swimtime="00:05:59.35" />
                    <SPLIT distance="550" swimtime="00:06:35.98" />
                    <SPLIT distance="600" swimtime="00:07:12.70" />
                    <SPLIT distance="650" swimtime="00:07:48.97" />
                    <SPLIT distance="700" swimtime="00:08:24.91" />
                    <SPLIT distance="750" swimtime="00:09:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="702" swimtime="00:02:40.77" resultid="7569" heatid="11459" lane="4" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:58.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="657" reactiontime="+77" swimtime="00:02:24.99" resultid="7570" heatid="11504" lane="3" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="706" swimtime="00:02:06.90" resultid="7571" heatid="11569" lane="4" entrytime="00:02:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="664" reactiontime="+78" swimtime="00:05:10.65" resultid="7572" heatid="11579" lane="3" entrytime="00:05:05.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:50.93" />
                    <SPLIT distance="200" swimtime="00:02:32.95" />
                    <SPLIT distance="250" swimtime="00:03:16.79" />
                    <SPLIT distance="300" swimtime="00:04:01.32" />
                    <SPLIT distance="350" swimtime="00:04:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="707" reactiontime="+82" swimtime="00:01:03.54" resultid="7573" heatid="11596" lane="8" entrytime="00:01:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="668" reactiontime="+78" swimtime="00:04:35.23" resultid="7574" heatid="11638" lane="7" entrytime="00:04:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:42.15" />
                    <SPLIT distance="200" swimtime="00:02:17.11" />
                    <SPLIT distance="250" swimtime="00:02:51.90" />
                    <SPLIT distance="300" swimtime="00:03:26.36" />
                    <SPLIT distance="350" swimtime="00:04:01.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03401" nation="POL" clubid="7584" name="UKS PATOMSWIM Bogatynia">
          <ATHLETES>
            <ATHLETE firstname="Tadeusz" lastname="Okorski" birthdate="1950-05-17" gender="M" nation="POL" license="103401700042" athleteid="7585">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7586" heatid="11404" lane="9" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="7587" heatid="11443" lane="5" />
                <RESULT eventid="6272" status="DNS" swimtime="00:00:00.00" resultid="7588" heatid="11455" lane="5" />
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="7589" heatid="11514" lane="8" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="7590" heatid="11548" lane="7" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="7591" heatid="11601" lane="4" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7592" heatid="11613" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8371" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Paszkiewicz" birthdate="1975-01-01" gender="M" nation="POL" athleteid="8370">
              <RESULTS>
                <RESULT eventid="6077" points="389" reactiontime="+68" swimtime="00:00:32.69" resultid="8372" heatid="11407" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="6306" points="292" reactiontime="+49" swimtime="00:01:19.71" resultid="8373" heatid="11470" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="285" swimtime="00:00:38.99" resultid="8374" heatid="11534" lane="9" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8396" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Szymaniak" birthdate="1993-01-01" gender="M" nation="POL" athleteid="8395">
              <RESULTS>
                <RESULT eventid="6077" points="315" reactiontime="+84" swimtime="00:00:33.55" resultid="8397" heatid="11403" lane="5" />
                <RESULT eventid="6306" points="263" reactiontime="+81" swimtime="00:01:15.82" resultid="8398" heatid="11467" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="244" reactiontime="+79" swimtime="00:00:37.89" resultid="8399" heatid="11531" lane="0" />
                <RESULT eventid="6535" points="225" reactiontime="+80" swimtime="00:03:02.72" resultid="8400" heatid="11562" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:01.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="246" reactiontime="+81" swimtime="00:06:26.18" resultid="8401" heatid="11629" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                    <SPLIT distance="200" swimtime="00:03:03.99" />
                    <SPLIT distance="250" swimtime="00:03:53.46" />
                    <SPLIT distance="300" swimtime="00:04:44.85" />
                    <SPLIT distance="350" swimtime="00:05:35.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7489" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Stasiukiewicz" birthdate="1980-01-01" gender="M" nation="POL" athleteid="7488">
              <RESULTS>
                <RESULT eventid="6238" points="139" reactiontime="+103" swimtime="00:00:52.35" resultid="7490" heatid="11445" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="6306" points="181" reactiontime="+107" swimtime="00:01:30.60" resultid="7491" heatid="11470" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="130" reactiontime="+104" swimtime="00:01:56.58" resultid="7492" heatid="11549" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7493" heatid="11564" lane="4" entrytime="00:02:55.00" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="7494" heatid="11603" lane="0" entrytime="00:03:50.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7495" heatid="11632" lane="1" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11341" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-01-01" gender="M" nation="POL" swrid="4062177" athleteid="8361">
              <RESULTS>
                <RESULT eventid="6077" points="864" reactiontime="+71" swimtime="00:00:23.23" resultid="8363" heatid="11419" lane="7" entrytime="00:00:23.34" entrycourse="SCM" />
                <RESULT eventid="6238" points="886" reactiontime="+74" swimtime="00:00:27.59" resultid="8364" heatid="11449" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="6306" points="854" swimtime="00:00:51.68" resultid="8365" heatid="11479" lane="4" entrytime="00:00:51.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="791" reactiontime="+65" swimtime="00:00:24.72" resultid="8366" heatid="11542" lane="6" entrytime="00:00:24.35" entrycourse="SCM" />
                <RESULT eventid="6535" points="724" reactiontime="+70" swimtime="00:01:58.62" resultid="8367" heatid="11570" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                    <SPLIT distance="150" swimtime="00:01:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="729" reactiontime="+67" swimtime="00:00:58.46" resultid="8368" heatid="11596" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="688" reactiontime="+74" swimtime="00:04:32.08" resultid="8369" heatid="11637" lane="2" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="100" swimtime="00:01:01.28" />
                    <SPLIT distance="150" swimtime="00:01:34.80" />
                    <SPLIT distance="200" swimtime="00:02:09.65" />
                    <SPLIT distance="250" swimtime="00:02:44.74" />
                    <SPLIT distance="300" swimtime="00:03:19.77" />
                    <SPLIT distance="350" swimtime="00:03:56.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="8990" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Mendowska" birthdate="1997-07-13" gender="F" nation="POL" license="100115600340" swrid="4229190" athleteid="9080">
              <RESULTS>
                <RESULT eventid="6323" points="548" swimtime="00:01:17.95" resultid="9081" heatid="11481" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="9082" heatid="11523" lane="8" />
                <RESULT eventid="6484" status="DNS" swimtime="00:00:00.00" resultid="9083" heatid="11543" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" swrid="4992782" athleteid="9013">
              <RESULTS>
                <RESULT eventid="6077" points="803" reactiontime="+67" swimtime="00:00:28.00" resultid="9014" heatid="11402" lane="2" />
                <RESULT eventid="6238" points="766" reactiontime="+67" swimtime="00:00:32.07" resultid="9015" heatid="11448" lane="2" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="6501" points="811" reactiontime="+73" swimtime="00:01:09.43" resultid="9016" heatid="11552" lane="8" entrytime="00:01:10.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="767" reactiontime="+81" swimtime="00:02:18.38" resultid="9017" heatid="11568" lane="2" entrytime="00:02:18.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="787" reactiontime="+69" swimtime="00:02:35.12" resultid="9018" heatid="11605" lane="3" entrytime="00:02:37.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="705" reactiontime="+81" swimtime="00:05:03.09" resultid="9019" heatid="11629" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:49.88" />
                    <SPLIT distance="200" swimtime="00:02:28.27" />
                    <SPLIT distance="250" swimtime="00:03:07.26" />
                    <SPLIT distance="300" swimtime="00:03:46.53" />
                    <SPLIT distance="350" swimtime="00:04:26.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Osik" birthdate="1976-01-02" gender="M" nation="POL" license="500115700521" swrid="5506634" athleteid="9073">
              <RESULTS>
                <RESULT eventid="6203" status="DNS" swimtime="00:00:00.00" resultid="9074" heatid="11654" lane="2" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="9075" heatid="11442" lane="4" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="9076" heatid="11548" lane="0" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="9077" heatid="11561" lane="4" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="9078" heatid="11606" lane="9" entrytime="00:02:32.97" entrycourse="SCM" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9079" heatid="11630" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Zajączek" birthdate="1976-07-17" gender="F" nation="POL" license="500115600524" swrid="5455051" athleteid="8991">
              <RESULTS>
                <RESULT eventid="6059" points="139" swimtime="00:00:51.87" resultid="8992" heatid="11395" lane="1" />
                <RESULT eventid="6094" points="155" swimtime="00:04:38.85" resultid="8993" heatid="11420" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.89" />
                    <SPLIT distance="100" swimtime="00:02:27.07" />
                    <SPLIT distance="150" swimtime="00:03:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="276" swimtime="00:04:19.75" resultid="8994" heatid="11451" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.62" />
                    <SPLIT distance="100" swimtime="00:02:05.21" />
                    <SPLIT distance="150" swimtime="00:03:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="90" swimtime="00:05:25.78" resultid="8995" heatid="11498" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.79" />
                    <SPLIT distance="100" swimtime="00:02:33.24" />
                    <SPLIT distance="150" swimtime="00:04:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="227" swimtime="00:02:07.06" resultid="8996" heatid="11509" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="92" swimtime="00:01:06.39" resultid="8997" heatid="11523" lane="7" />
                <RESULT eventid="6618" points="96" swimtime="00:02:23.81" resultid="8998" heatid="11586" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="196" swimtime="00:00:59.81" resultid="8999" heatid="11607" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Majchrzak" birthdate="1983-01-21" gender="M" nation="POL" license="100115700630" swrid="4431795" athleteid="9084">
              <RESULTS>
                <RESULT eventid="6467" points="559" reactiontime="+75" swimtime="00:00:28.68" resultid="9085" heatid="11530" lane="6" />
                <RESULT eventid="6535" points="621" reactiontime="+79" swimtime="00:02:10.65" resultid="9086" heatid="11560" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:03.38" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="564" swimtime="00:01:06.80" resultid="9087" heatid="11590" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="581" reactiontime="+86" swimtime="00:04:50.33" resultid="9088" heatid="11629" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                    <SPLIT distance="200" swimtime="00:02:22.70" />
                    <SPLIT distance="250" swimtime="00:02:59.82" />
                    <SPLIT distance="300" swimtime="00:03:37.71" />
                    <SPLIT distance="350" swimtime="00:04:15.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" swrid="5062813" athleteid="9020">
              <RESULTS>
                <RESULT eventid="6077" points="758" reactiontime="+71" swimtime="00:00:24.27" resultid="9021" heatid="11418" lane="2" entrytime="00:00:24.34" entrycourse="SCM" />
                <RESULT eventid="6306" points="760" reactiontime="+73" swimtime="00:00:53.72" resultid="9022" heatid="11479" lane="7" entrytime="00:00:53.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="653" reactiontime="+70" swimtime="00:00:26.35" resultid="9023" heatid="11541" lane="3" entrytime="00:00:26.52" entrycourse="SCM" />
                <RESULT eventid="6535" points="692" reactiontime="+69" swimtime="00:02:00.40" resultid="9024" heatid="11570" lane="3" entrytime="00:02:04.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="100" swimtime="00:00:57.47" />
                    <SPLIT distance="150" swimtime="00:01:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="662" reactiontime="+70" swimtime="00:01:00.36" resultid="9025" heatid="11595" lane="3" entrytime="00:01:03.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" swrid="4595659" athleteid="9068">
              <RESULTS>
                <RESULT eventid="6169" points="486" reactiontime="+94" swimtime="00:10:50.74" resultid="9069" heatid="11645" lane="8" entrytime="00:10:20.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                    <SPLIT distance="150" swimtime="00:01:57.08" />
                    <SPLIT distance="200" swimtime="00:02:37.72" />
                    <SPLIT distance="250" swimtime="00:03:18.88" />
                    <SPLIT distance="300" swimtime="00:04:00.24" />
                    <SPLIT distance="350" swimtime="00:04:41.70" />
                    <SPLIT distance="400" swimtime="00:05:23.10" />
                    <SPLIT distance="450" swimtime="00:06:04.59" />
                    <SPLIT distance="500" swimtime="00:06:45.77" />
                    <SPLIT distance="550" swimtime="00:07:27.44" />
                    <SPLIT distance="600" swimtime="00:08:09.05" />
                    <SPLIT distance="650" swimtime="00:08:50.20" />
                    <SPLIT distance="700" swimtime="00:09:31.53" />
                    <SPLIT distance="750" swimtime="00:10:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="441" reactiontime="+83" swimtime="00:02:45.52" resultid="9070" heatid="11504" lane="1" entrytime="00:02:38.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="9071" heatid="11568" lane="3" entrytime="00:02:16.80" entrycourse="SCM" />
                <RESULT eventid="6738" points="481" reactiontime="+85" swimtime="00:05:06.96" resultid="9072" heatid="11636" lane="7" entrytime="00:04:57.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:52.69" />
                    <SPLIT distance="200" swimtime="00:02:31.69" />
                    <SPLIT distance="250" swimtime="00:03:10.94" />
                    <SPLIT distance="300" swimtime="00:03:50.30" />
                    <SPLIT distance="350" swimtime="00:04:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Bartkowiak" birthdate="1949-03-13" gender="M" nation="POL" license="100115700738" athleteid="9047">
              <RESULTS>
                <RESULT eventid="6111" points="340" reactiontime="+103" swimtime="00:04:14.62" resultid="9048" heatid="11426" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.86" />
                    <SPLIT distance="100" swimtime="00:02:10.02" />
                    <SPLIT distance="150" swimtime="00:03:20.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="531" swimtime="00:28:30.14" resultid="9049" heatid="11654" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                    <SPLIT distance="100" swimtime="00:01:43.88" />
                    <SPLIT distance="150" swimtime="00:02:40.60" />
                    <SPLIT distance="200" swimtime="00:03:37.89" />
                    <SPLIT distance="250" swimtime="00:04:35.46" />
                    <SPLIT distance="300" swimtime="00:05:32.77" />
                    <SPLIT distance="350" swimtime="00:06:30.68" />
                    <SPLIT distance="400" swimtime="00:07:27.99" />
                    <SPLIT distance="450" swimtime="00:08:26.42" />
                    <SPLIT distance="500" swimtime="00:09:24.00" />
                    <SPLIT distance="550" swimtime="00:10:21.41" />
                    <SPLIT distance="600" swimtime="00:11:18.44" />
                    <SPLIT distance="650" swimtime="00:12:16.53" />
                    <SPLIT distance="700" swimtime="00:13:14.40" />
                    <SPLIT distance="750" swimtime="00:14:11.42" />
                    <SPLIT distance="800" swimtime="00:15:09.57" />
                    <SPLIT distance="850" swimtime="00:16:06.59" />
                    <SPLIT distance="900" swimtime="00:17:04.82" />
                    <SPLIT distance="950" swimtime="00:18:02.12" />
                    <SPLIT distance="1000" swimtime="00:18:59.64" />
                    <SPLIT distance="1050" swimtime="00:19:56.83" />
                    <SPLIT distance="1100" swimtime="00:20:54.59" />
                    <SPLIT distance="1150" swimtime="00:21:52.36" />
                    <SPLIT distance="1200" swimtime="00:22:50.20" />
                    <SPLIT distance="1250" swimtime="00:23:48.19" />
                    <SPLIT distance="1300" swimtime="00:24:45.92" />
                    <SPLIT distance="1350" swimtime="00:25:43.45" />
                    <SPLIT distance="1400" swimtime="00:26:40.92" />
                    <SPLIT distance="1450" swimtime="00:27:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="380" reactiontime="+80" swimtime="00:04:15.63" resultid="9050" heatid="11455" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.70" />
                    <SPLIT distance="100" swimtime="00:02:02.53" />
                    <SPLIT distance="150" swimtime="00:03:10.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2 - Pływak pokonał jednym stylem więcej niż 1 dystansu." eventid="6340" reactiontime="+109" status="DSQ" swimtime="00:00:00.00" resultid="9051" heatid="11487" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="335" reactiontime="+94" swimtime="00:01:58.69" resultid="9052" heatid="11514" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="403" reactiontime="+98" swimtime="00:03:20.34" resultid="9053" heatid="11560" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:34.39" />
                    <SPLIT distance="150" swimtime="00:02:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="102" reactiontime="+104" swimtime="00:02:41.67" resultid="9054" heatid="11590" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="443" swimtime="00:07:10.04" resultid="9055" heatid="11630" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                    <SPLIT distance="150" swimtime="00:02:32.85" />
                    <SPLIT distance="200" swimtime="00:03:29.72" />
                    <SPLIT distance="250" swimtime="00:04:25.24" />
                    <SPLIT distance="300" swimtime="00:05:20.62" />
                    <SPLIT distance="350" swimtime="00:06:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" swrid="5312534" athleteid="9031">
              <RESULTS>
                <RESULT eventid="6077" points="724" swimtime="00:00:25.84" resultid="9032" heatid="11416" lane="4" entrytime="00:00:25.64" entrycourse="SCM" />
                <RESULT eventid="6111" points="664" reactiontime="+79" swimtime="00:02:26.55" resultid="9033" heatid="11426" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6272" points="821" reactiontime="+80" swimtime="00:02:32.55" resultid="9034" heatid="11459" lane="5" entrytime="00:02:43.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="881" swimtime="00:01:02.39" resultid="9035" heatid="11495" lane="4" entrytime="00:01:06.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6433" points="854" reactiontime="+72" swimtime="00:01:07.02" resultid="9036" heatid="11521" lane="0" entrytime="00:01:08.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="716" reactiontime="+67" swimtime="00:00:28.09" resultid="9037" heatid="11540" lane="2" entrytime="00:00:27.84" entrycourse="SCM" />
                <RESULT eventid="6704" points="876" reactiontime="+71" swimtime="00:00:30.39" resultid="9038" heatid="11623" lane="9" entrytime="00:00:30.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="9000">
              <RESULTS>
                <RESULT eventid="6059" points="85" swimtime="00:01:01.04" resultid="9001" heatid="11395" lane="6" />
                <RESULT eventid="6255" points="217" swimtime="00:04:41.28" resultid="9002" heatid="11452" lane="1" entrytime="00:04:46.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.92" />
                    <SPLIT distance="100" swimtime="00:02:14.94" />
                    <SPLIT distance="150" swimtime="00:03:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="130" reactiontime="+115" swimtime="00:02:16.32" resultid="9003" heatid="11482" lane="7" entrytime="00:02:13.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="190" reactiontime="+102" swimtime="00:02:14.69" resultid="9004" heatid="11510" lane="0" entrytime="00:02:10.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="207" reactiontime="+105" swimtime="00:00:58.72" resultid="9005" heatid="11609" lane="5" entrytime="00:00:57.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Wiśniewska" birthdate="1997-10-01" gender="F" nation="POL" license="500115600544" swrid="4273989" athleteid="9039">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /K1" eventid="6094" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="9040" heatid="11420" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="737" reactiontime="+82" swimtime="00:10:16.13" resultid="9041" heatid="11644" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:48.77" />
                    <SPLIT distance="200" swimtime="00:02:27.61" />
                    <SPLIT distance="250" swimtime="00:03:07.54" />
                    <SPLIT distance="300" swimtime="00:03:46.72" />
                    <SPLIT distance="350" swimtime="00:04:26.27" />
                    <SPLIT distance="400" swimtime="00:05:04.98" />
                    <SPLIT distance="450" swimtime="00:05:44.24" />
                    <SPLIT distance="500" swimtime="00:06:24.00" />
                    <SPLIT distance="550" swimtime="00:07:03.75" />
                    <SPLIT distance="600" swimtime="00:07:43.09" />
                    <SPLIT distance="650" swimtime="00:08:22.46" />
                    <SPLIT distance="700" swimtime="00:09:01.11" />
                    <SPLIT distance="750" swimtime="00:09:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6255" points="892" swimtime="00:02:39.62" resultid="9042" heatid="11454" lane="4" entrytime="00:02:41.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="794" reactiontime="+82" swimtime="00:01:08.88" resultid="9043" heatid="11481" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="830" reactiontime="+83" swimtime="00:01:15.15" resultid="9044" heatid="11508" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="804" reactiontime="+88" swimtime="00:05:22.81" resultid="9045" heatid="11573" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                    <SPLIT distance="200" swimtime="00:02:36.90" />
                    <SPLIT distance="250" swimtime="00:03:21.16" />
                    <SPLIT distance="300" swimtime="00:04:05.66" />
                    <SPLIT distance="350" swimtime="00:04:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="9046" heatid="11608" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" swrid="4992790" athleteid="9006">
              <RESULTS>
                <RESULT eventid="6059" points="260" reactiontime="+114" swimtime="00:00:50.47" resultid="9007" heatid="11393" lane="3" />
                <RESULT eventid="6255" points="457" reactiontime="+109" swimtime="00:04:20.63" resultid="9008" heatid="11452" lane="6" entrytime="00:04:14.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                    <SPLIT distance="100" swimtime="00:02:09.15" />
                    <SPLIT distance="150" swimtime="00:03:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="229" reactiontime="+111" swimtime="00:01:55.93" resultid="9009" heatid="11461" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="409" reactiontime="+108" swimtime="00:01:59.14" resultid="9010" heatid="11509" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="250" reactiontime="+114" swimtime="00:04:20.16" resultid="9011" heatid="11555" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.60" />
                    <SPLIT distance="100" swimtime="00:02:04.98" />
                    <SPLIT distance="150" swimtime="00:03:14.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="389" swimtime="00:00:53.25" resultid="9012" heatid="11610" lane="8" entrytime="00:00:53.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" swrid="4213120" athleteid="9026">
              <RESULTS>
                <RESULT eventid="6077" points="908" reactiontime="+62" swimtime="00:00:23.58" resultid="9027" heatid="11419" lane="0" entrytime="00:00:23.55" entrycourse="SCM" />
                <RESULT eventid="6306" points="798" reactiontime="+64" swimtime="00:00:52.37" resultid="9028" heatid="11479" lane="5" entrytime="00:00:51.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="816" reactiontime="+66" swimtime="00:00:25.36" resultid="9029" heatid="11531" lane="2" />
                <RESULT eventid="6636" points="837" reactiontime="+67" swimtime="00:00:57.21" resultid="9030" heatid="11597" lane="7" entrytime="00:00:56.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="9056">
              <RESULTS>
                <RESULT eventid="6111" points="627" reactiontime="+90" swimtime="00:02:58.57" resultid="9057" heatid="11426" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="150" swimtime="00:02:16.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="669" swimtime="00:03:09.66" resultid="9058" heatid="11455" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.79" />
                    <SPLIT distance="150" swimtime="00:02:18.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="628" reactiontime="+88" swimtime="00:01:26.26" resultid="9059" heatid="11513" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="612" swimtime="00:00:38.55" resultid="9060" heatid="11614" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+72" swimtime="00:01:37.97" resultid="9094" heatid="11584" lane="4" entrytime="00:01:37.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.19" />
                    <SPLIT distance="100" swimtime="00:00:49.24" />
                    <SPLIT distance="150" swimtime="00:01:15.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9020" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9031" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="9084" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="9026" number="4" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" reactiontime="+73" swimtime="00:01:49.84" resultid="9097" heatid="12332" lane="4" entrytime="00:01:49.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:00:58.62" />
                    <SPLIT distance="150" swimtime="00:01:23.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9020" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="9031" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="9026" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="9084" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+69" swimtime="00:01:50.74" resultid="9089" heatid="11436" lane="5" entrytime="00:01:48.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.47" />
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                    <SPLIT distance="150" swimtime="00:01:25.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9020" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="9039" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="9080" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9031" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+78" swimtime="00:02:00.49" resultid="9091" heatid="11507" lane="5" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:31.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9020" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="9031" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="9080" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9039" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+73" swimtime="00:02:54.57" resultid="9090" heatid="11435" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:01:00.68" />
                    <SPLIT distance="150" swimtime="00:01:53.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9013" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="9056" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="9006" number="3" reactiontime="+87" />
                    <RELAYPOSITION athleteid="9000" number="4" reactiontime="+94" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+59" swimtime="00:03:17.44" resultid="9092" heatid="11506" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:02:18.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9013" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="9056" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="8991" number="3" />
                    <RELAYPOSITION athleteid="9000" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" clubid="7452" name="Uks Delfin Legionowo">
          <ATHLETES>
            <ATHLETE firstname="Andzrej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" license="101414700141" athleteid="7453">
              <RESULTS>
                <RESULT eventid="6077" points="476" reactiontime="+83" swimtime="00:00:30.56" resultid="7454" heatid="11410" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="6238" points="369" reactiontime="+88" swimtime="00:00:38.85" resultid="7455" heatid="11446" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="6306" points="407" reactiontime="+71" swimtime="00:01:11.39" resultid="7456" heatid="11473" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="346" reactiontime="+78" swimtime="00:01:24.56" resultid="7457" heatid="11550" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="320" reactiontime="+78" swimtime="00:02:47.61" resultid="7458" heatid="11566" lane="8" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:03.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="343" reactiontime="+84" swimtime="00:03:07.83" resultid="7459" heatid="11604" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michałj" lastname="Perl" birthdate="1996-06-07" gender="M" nation="POL" license="101414700068" swrid="4282344" athleteid="7460">
              <RESULTS>
                <RESULT eventid="6704" points="891" reactiontime="+65" swimtime="00:00:29.36" resultid="7461" heatid="11623" lane="3" entrytime="00:00:28.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Żbikowska" birthdate="1996-01-01" gender="F" nation="POL" license="S01414100028" swrid="4605445" athleteid="7462">
              <RESULTS>
                <RESULT eventid="6059" points="601" reactiontime="+76" swimtime="00:00:29.96" resultid="7463" heatid="11400" lane="0" entrytime="00:00:30.12" />
                <RESULT eventid="6094" points="620" reactiontime="+83" swimtime="00:02:45.28" resultid="7464" heatid="11423" lane="3" entrytime="00:02:50.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:02:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="628" reactiontime="+84" swimtime="00:02:59.43" resultid="7465" heatid="11454" lane="6" entrytime="00:03:02.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="615" reactiontime="+81" swimtime="00:01:15.01" resultid="7466" heatid="11486" lane="9" entrytime="00:01:15.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="676" reactiontime="+82" swimtime="00:01:20.49" resultid="7467" heatid="11512" lane="1" entrytime="00:01:22.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="657" swimtime="00:00:31.73" resultid="7468" heatid="11527" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="6687" points="690" reactiontime="+80" swimtime="00:00:35.74" resultid="7469" heatid="11612" lane="2" entrytime="00:00:36.19" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="9099" name="Masters Avia Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Lis" birthdate="1996-04-03" gender="M" nation="POL" license="104303700011" swrid="4251399" athleteid="9121">
              <RESULTS>
                <RESULT eventid="6169" points="696" reactiontime="+72" swimtime="00:09:36.78" resultid="9122" heatid="11645" lane="5" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="150" swimtime="00:01:40.37" />
                    <SPLIT distance="200" swimtime="00:02:15.71" />
                    <SPLIT distance="250" swimtime="00:02:50.88" />
                    <SPLIT distance="300" swimtime="00:03:25.62" />
                    <SPLIT distance="350" swimtime="00:04:00.73" />
                    <SPLIT distance="400" swimtime="00:04:36.54" />
                    <SPLIT distance="450" swimtime="00:05:12.33" />
                    <SPLIT distance="500" swimtime="00:05:48.84" />
                    <SPLIT distance="550" swimtime="00:06:25.96" />
                    <SPLIT distance="600" swimtime="00:07:03.56" />
                    <SPLIT distance="650" swimtime="00:07:41.77" />
                    <SPLIT distance="700" swimtime="00:08:20.46" />
                    <SPLIT distance="750" swimtime="00:08:58.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="709" reactiontime="+75" swimtime="00:00:54.47" resultid="9123" heatid="11479" lane="9" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="761" reactiontime="+72" swimtime="00:02:01.76" resultid="9124" heatid="11571" lane="6" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:00.25" />
                    <SPLIT distance="150" swimtime="00:01:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="758" reactiontime="+74" swimtime="00:04:25.58" resultid="9125" heatid="11638" lane="6" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:03.86" />
                    <SPLIT distance="150" swimtime="00:01:37.14" />
                    <SPLIT distance="200" swimtime="00:02:10.71" />
                    <SPLIT distance="250" swimtime="00:02:44.20" />
                    <SPLIT distance="300" swimtime="00:03:17.90" />
                    <SPLIT distance="350" swimtime="00:03:52.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" swrid="5439542" athleteid="9108">
              <RESULTS>
                <RESULT eventid="6077" points="680" swimtime="00:00:27.14" resultid="9109" heatid="11414" lane="1" entrytime="00:00:27.51" />
                <RESULT eventid="6238" points="718" reactiontime="+61" swimtime="00:00:31.12" resultid="9110" heatid="11448" lane="4" entrytime="00:00:31.94" />
                <RESULT eventid="6340" points="635" reactiontime="+70" swimtime="00:01:09.78" resultid="9111" heatid="11495" lane="0" entrytime="00:01:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="625" reactiontime="+71" swimtime="00:01:09.47" resultid="9112" heatid="11552" lane="7" entrytime="00:01:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="539" reactiontime="+67" swimtime="00:02:41.68" resultid="9113" heatid="11605" lane="9" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:01:59.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" swrid="4061691" athleteid="9114">
              <RESULTS>
                <RESULT eventid="6077" points="650" swimtime="00:00:25.43" resultid="9115" heatid="11417" lane="1" entrytime="00:00:25.30" />
                <RESULT eventid="6306" points="705" reactiontime="+74" swimtime="00:00:55.47" resultid="9116" heatid="11478" lane="7" entrytime="00:00:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="568" reactiontime="+67" swimtime="00:00:28.53" resultid="9117" heatid="11540" lane="7" entrytime="00:00:27.99" />
                <RESULT eventid="6535" points="698" reactiontime="+78" swimtime="00:02:05.64" resultid="9118" heatid="11571" lane="9" entrytime="00:02:03.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:01.06" />
                    <SPLIT distance="150" swimtime="00:01:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="647" reactiontime="+69" swimtime="00:01:03.80" resultid="9119" heatid="11595" lane="4" entrytime="00:01:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="672" reactiontime="+69" swimtime="00:04:36.55" resultid="9120" heatid="11637" lane="5" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:40.41" />
                    <SPLIT distance="200" swimtime="00:02:16.04" />
                    <SPLIT distance="250" swimtime="00:02:51.70" />
                    <SPLIT distance="300" swimtime="00:03:26.49" />
                    <SPLIT distance="350" swimtime="00:04:01.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Wółkiewicz" birthdate="1987-03-01" gender="M" nation="POL" license="504303700012" swrid="4633330" athleteid="9126">
              <RESULTS>
                <RESULT eventid="6704" points="663" reactiontime="+88" swimtime="00:00:33.09" resultid="9127" heatid="11622" lane="6" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="9100">
              <RESULTS>
                <RESULT eventid="6077" points="650" reactiontime="+72" swimtime="00:00:28.27" resultid="9101" heatid="11411" lane="3" entrytime="00:00:29.94" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6203" points="647" reactiontime="+75" swimtime="00:19:36.03" resultid="9102" heatid="11652" lane="0" entrytime="00:21:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="550" swimtime="00:07:07.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="626" reactiontime="+80" swimtime="00:01:02.06" resultid="9103" heatid="11475" lane="9" entrytime="00:01:03.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="475" reactiontime="+79" swimtime="00:01:15.98" resultid="9104" heatid="11492" lane="5" entrytime="00:01:15.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="545" reactiontime="+69" swimtime="00:00:32.81" resultid="9105" heatid="11535" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="6535" points="596" reactiontime="+79" swimtime="00:02:20.31" resultid="9106" heatid="11567" lane="8" entrytime="00:02:30.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="677" reactiontime="+77" swimtime="00:04:56.55" resultid="9107" heatid="11636" lane="9" entrytime="00:05:00.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                    <SPLIT distance="200" swimtime="00:02:26.62" />
                    <SPLIT distance="250" swimtime="00:03:04.45" />
                    <SPLIT distance="300" swimtime="00:03:42.49" />
                    <SPLIT distance="350" swimtime="00:04:20.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+70" swimtime="00:01:44.77" resultid="9128" heatid="11584" lane="6" entrytime="00:01:45.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                    <SPLIT distance="100" swimtime="00:00:53.13" />
                    <SPLIT distance="150" swimtime="00:01:19.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9121" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="9100" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="9108" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="9114" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+57" swimtime="00:01:57.81" resultid="9129" heatid="12332" lane="3" entrytime="00:01:58.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:33.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9108" number="1" reactiontime="+57" />
                    <RELAYPOSITION athleteid="9126" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="9114" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="9121" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6871" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jarosław" lastname="Guziński" birthdate="1966-01-01" gender="M" nation="POL" swrid="5484405" athleteid="6870">
              <RESULTS>
                <RESULT eventid="6374" status="DNS" swimtime="00:00:00.00" resultid="6872" heatid="11500" lane="4" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="6873" heatid="11532" lane="6" entrytime="00:00:43.17" entrycourse="SCM" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="6874" heatid="11591" lane="8" entrytime="00:01:45.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7349" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Skurczyńska" birthdate="1971-01-01" gender="F" nation="POL" athleteid="7348">
              <RESULTS>
                <RESULT eventid="6059" points="279" reactiontime="+80" swimtime="00:00:43.25" resultid="7350" heatid="11396" lane="3" entrytime="00:00:43.53" />
                <RESULT eventid="6255" points="270" reactiontime="+81" swimtime="00:04:19.97" resultid="7351" heatid="11452" lane="3" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.14" />
                    <SPLIT distance="100" swimtime="00:01:55.81" />
                    <SPLIT distance="150" swimtime="00:03:07.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="364" reactiontime="+83" swimtime="00:01:47.90" resultid="7352" heatid="11510" lane="3" entrytime="00:01:55.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="216" reactiontime="+91" swimtime="00:00:51.91" resultid="7353" heatid="11524" lane="7" entrytime="00:00:55.37" />
                <RESULT eventid="6687" points="401" reactiontime="+79" swimtime="00:00:48.53" resultid="7354" heatid="11610" lane="1" entrytime="00:00:52.01" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06711" nation="POL" clubid="11343" name="UKS DRAGON Będzin">
          <ATHLETES>
            <ATHLETE firstname="Emil" lastname="Strumiński" birthdate="1988-05-18" gender="M" nation="POL" license="306711700032" athleteid="11344">
              <RESULTS>
                <RESULT eventid="6077" points="634" reactiontime="+69" swimtime="00:00:25.76" resultid="11345" heatid="11403" lane="8" />
                <RESULT eventid="6111" points="518" reactiontime="+72" swimtime="00:02:27.04" resultid="11346" heatid="11432" lane="4" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:55.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="672" reactiontime="+71" swimtime="00:00:55.97" resultid="11347" heatid="11478" lane="2" entrytime="00:00:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="532" reactiontime="+77" swimtime="00:02:32.98" resultid="11348" heatid="11504" lane="6" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="11349" heatid="11540" lane="4" entrytime="00:00:27.40" />
                <RESULT eventid="6535" points="613" reactiontime="+72" swimtime="00:02:05.33" resultid="11350" heatid="11570" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:00.80" />
                    <SPLIT distance="150" swimtime="00:01:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="579" reactiontime="+78" swimtime="00:01:03.13" resultid="11351" heatid="11596" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="659" reactiontime="+78" swimtime="00:04:35.97" resultid="11352" heatid="11629" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                    <SPLIT distance="200" swimtime="00:02:18.13" />
                    <SPLIT distance="250" swimtime="00:02:53.99" />
                    <SPLIT distance="300" swimtime="00:03:29.53" />
                    <SPLIT distance="350" swimtime="00:04:04.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7254" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Kamil" lastname="Lubiński" birthdate="1992-01-01" gender="M" nation="POL" swrid="4264463" athleteid="7253">
              <RESULTS>
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7255" heatid="11430" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="6169" status="OTL" swimtime="00:00:00.00" resultid="7256" heatid="11645" lane="9" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:01:55.16" />
                    <SPLIT distance="200" swimtime="00:02:35.23" />
                    <SPLIT distance="250" swimtime="00:03:15.00" />
                    <SPLIT distance="300" swimtime="00:03:54.70" />
                    <SPLIT distance="350" swimtime="00:04:34.69" />
                    <SPLIT distance="400" swimtime="00:05:14.65" />
                    <SPLIT distance="450" swimtime="00:05:55.06" />
                    <SPLIT distance="500" swimtime="00:06:35.58" />
                    <SPLIT distance="550" swimtime="00:07:16.14" />
                    <SPLIT distance="600" swimtime="00:07:57.44" />
                    <SPLIT distance="650" swimtime="00:08:39.13" />
                    <SPLIT distance="700" swimtime="00:09:20.40" />
                    <SPLIT distance="750" swimtime="00:10:01.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="499" reactiontime="+80" swimtime="00:00:33.41" resultid="7257" heatid="11448" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="6340" points="486" reactiontime="+79" swimtime="00:01:09.92" resultid="7258" heatid="11493" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="446" reactiontime="+84" swimtime="00:02:19.32" resultid="7259" heatid="11568" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="7260" heatid="11578" lane="2" entrytime="00:05:50.00" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="7261" heatid="11594" lane="0" entrytime="00:01:10.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7262" heatid="11635" lane="4" entrytime="00:05:05.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00101" nation="POL" region="01" clubid="9216" name="MKS Juvenia Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Makowski" birthdate="1996-01-02" gender="M" nation="POL" license="100101701205" swrid="4283690" athleteid="9217">
              <RESULTS>
                <RESULT eventid="6077" points="1010" reactiontime="+73" swimtime="00:00:22.76" resultid="9218" heatid="11419" lane="2" entrytime="00:00:23.05" entrycourse="SCM" />
                <RESULT eventid="6340" points="829" reactiontime="+76" swimtime="00:00:58.76" resultid="9219" heatid="11497" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="965" reactiontime="+72" swimtime="00:00:23.98" resultid="9220" heatid="11542" lane="3" entrytime="00:00:24.22" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6636" points="966" reactiontime="+75" swimtime="00:00:54.54" resultid="9221" heatid="11597" lane="6" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="9130" name="MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Wójcicka" birthdate="1975-05-28" gender="F" nation="POL" license="103503600002" swrid="5537484" athleteid="9148">
              <RESULTS>
                <RESULT eventid="6145" points="377" reactiontime="+99" swimtime="00:13:16.77" resultid="9149" heatid="11644" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:28.20" />
                    <SPLIT distance="150" swimtime="00:02:17.51" />
                    <SPLIT distance="200" swimtime="00:03:07.44" />
                    <SPLIT distance="250" swimtime="00:03:57.61" />
                    <SPLIT distance="300" swimtime="00:04:48.05" />
                    <SPLIT distance="350" swimtime="00:05:38.21" />
                    <SPLIT distance="400" swimtime="00:06:29.57" />
                    <SPLIT distance="450" swimtime="00:07:19.94" />
                    <SPLIT distance="500" swimtime="00:08:11.25" />
                    <SPLIT distance="550" swimtime="00:09:02.43" />
                    <SPLIT distance="600" swimtime="00:09:55.32" />
                    <SPLIT distance="650" swimtime="00:10:47.00" />
                    <SPLIT distance="700" swimtime="00:11:37.67" />
                    <SPLIT distance="750" swimtime="00:12:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="427" reactiontime="+95" swimtime="00:00:40.49" resultid="9150" heatid="11438" lane="0" />
                <RESULT eventid="6323" points="445" reactiontime="+90" swimtime="00:01:30.54" resultid="9151" heatid="11481" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="444" reactiontime="+93" swimtime="00:01:28.96" resultid="9152" heatid="11545" lane="3" entrytime="00:01:29.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="576" reactiontime="+104" swimtime="00:03:04.70" resultid="9153" heatid="11598" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:29.87" />
                    <SPLIT distance="150" swimtime="00:02:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="439" reactiontime="+102" swimtime="00:00:45.72" resultid="9154" heatid="11608" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-03-13" gender="M" nation="POL" license="103503700029" swrid="5558377" athleteid="9139">
              <RESULTS>
                <RESULT eventid="6077" points="511" reactiontime="+86" swimtime="00:00:27.55" resultid="9140" heatid="11402" lane="7" />
                <RESULT eventid="6111" points="416" reactiontime="+83" swimtime="00:02:50.42" resultid="9141" heatid="11425" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:11.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="504" reactiontime="+85" swimtime="00:01:02.00" resultid="9143" heatid="11475" lane="0" entrytime="00:01:03.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="454" reactiontime="+82" swimtime="00:01:13.86" resultid="9144" heatid="11492" lane="3" entrytime="00:01:16.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="489" reactiontime="+88" swimtime="00:00:29.99" resultid="9145" heatid="11536" lane="3" entrytime="00:00:31.61" entrycourse="SCM" />
                <RESULT eventid="6535" points="425" swimtime="00:02:28.17" resultid="9146" heatid="11560" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="439" reactiontime="+89" swimtime="00:01:12.63" resultid="9147" heatid="11589" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="408" reactiontime="+85" swimtime="00:00:38.89" resultid="11378" heatid="11614" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pietrzak" birthdate="1988-10-21" gender="M" nation="POL" license="103503700011" swrid="5537482" athleteid="9131">
              <RESULTS>
                <RESULT eventid="6077" points="393" reactiontime="+85" swimtime="00:00:30.20" resultid="9132" heatid="11404" lane="8" />
                <RESULT eventid="6238" points="440" reactiontime="+73" swimtime="00:00:34.83" resultid="9133" heatid="11442" lane="3" />
                <RESULT eventid="6340" points="353" reactiontime="+83" swimtime="00:01:17.77" resultid="9134" heatid="11487" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="386" reactiontime="+73" swimtime="00:01:19.04" resultid="9135" heatid="11547" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="270" reactiontime="+83" swimtime="00:02:44.73" resultid="9136" heatid="11560" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:01.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="297" reactiontime="+81" swimtime="00:02:54.67" resultid="9137" heatid="11602" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:02:10.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="363" reactiontime="+82" swimtime="00:00:38.96" resultid="9138" heatid="11615" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wójcicki" birthdate="1975-04-28" gender="M" nation="POL" license="103503700001" swrid="5455050" athleteid="9155">
              <RESULTS>
                <RESULT eventid="6238" points="435" reactiontime="+82" swimtime="00:00:36.76" resultid="9157" heatid="11444" lane="9" />
                <RESULT eventid="6340" points="420" swimtime="00:01:20.07" resultid="9158" heatid="11487" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="398" reactiontime="+83" swimtime="00:01:29.75" resultid="9159" heatid="11518" lane="0" entrytime="00:01:30.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="389" reactiontime="+84" swimtime="00:01:21.36" resultid="9160" heatid="11547" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="429" reactiontime="+84" swimtime="00:00:40.15" resultid="9161" heatid="11614" lane="1" />
                <RESULT eventid="6203" points="376" reactiontime="+85" swimtime="00:22:48.82" resultid="11386" heatid="11654" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                    <SPLIT distance="200" swimtime="00:02:49.91" />
                    <SPLIT distance="250" swimtime="00:03:35.16" />
                    <SPLIT distance="300" swimtime="00:04:20.63" />
                    <SPLIT distance="350" swimtime="00:05:06.48" />
                    <SPLIT distance="400" swimtime="00:06:38.31" />
                    <SPLIT distance="450" swimtime="00:07:23.88" />
                    <SPLIT distance="500" swimtime="00:08:09.33" />
                    <SPLIT distance="550" swimtime="00:08:55.68" />
                    <SPLIT distance="600" swimtime="00:09:41.31" />
                    <SPLIT distance="650" swimtime="00:10:27.59" />
                    <SPLIT distance="700" swimtime="00:11:14.29" />
                    <SPLIT distance="750" swimtime="00:12:00.56" />
                    <SPLIT distance="800" swimtime="00:12:46.73" />
                    <SPLIT distance="850" swimtime="00:13:33.39" />
                    <SPLIT distance="900" swimtime="00:14:19.35" />
                    <SPLIT distance="950" swimtime="00:15:05.43" />
                    <SPLIT distance="1000" swimtime="00:15:51.72" />
                    <SPLIT distance="1050" swimtime="00:16:38.19" />
                    <SPLIT distance="1100" swimtime="00:17:24.38" />
                    <SPLIT distance="1150" swimtime="00:18:10.73" />
                    <SPLIT distance="1200" swimtime="00:18:56.63" />
                    <SPLIT distance="1250" swimtime="00:19:43.29" />
                    <SPLIT distance="1300" swimtime="00:20:29.53" />
                    <SPLIT distance="1350" swimtime="00:21:16.42" />
                    <SPLIT distance="1400" swimtime="00:22:02.95" />
                    <SPLIT distance="1450" swimtime="00:22:48.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" swrid="5537480" athleteid="9162">
              <RESULTS>
                <RESULT eventid="6374" points="286" reactiontime="+100" swimtime="00:03:30.90" resultid="9163" heatid="11500" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.90" />
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                    <SPLIT distance="150" swimtime="00:02:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="377" reactiontime="+88" swimtime="00:00:37.09" resultid="9164" heatid="11533" lane="6" entrytime="00:00:39.04" entrycourse="SCM" />
                <RESULT eventid="6636" points="242" reactiontime="+99" swimtime="00:01:35.66" resultid="9165" heatid="11591" lane="2" entrytime="00:01:38.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="308" reactiontime="+124" swimtime="00:00:45.54" resultid="9166" heatid="11613" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7277" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jarosław" lastname="Tuszyński" birthdate="1975-01-01" gender="M" nation="POL" athleteid="7276">
              <RESULTS>
                <RESULT eventid="6272" points="423" reactiontime="+85" swimtime="00:03:16.55" resultid="7278" heatid="11458" lane="0" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="491" reactiontime="+87" swimtime="00:01:23.73" resultid="7279" heatid="11519" lane="0" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="546" reactiontime="+88" swimtime="00:00:37.04" resultid="7280" heatid="11619" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="100111" nation="POL" clubid="7593" name="UKS TRÓJKA  Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" swrid="4289072" athleteid="7611">
              <RESULTS>
                <RESULT eventid="6059" points="571" swimtime="00:00:30.47" resultid="7612" heatid="11399" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="6145" points="714" reactiontime="+83" swimtime="00:10:22.52" resultid="7613" heatid="11643" lane="6" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:55.94" />
                    <SPLIT distance="200" swimtime="00:02:35.27" />
                    <SPLIT distance="250" swimtime="00:03:14.30" />
                    <SPLIT distance="300" swimtime="00:03:53.29" />
                    <SPLIT distance="350" swimtime="00:04:32.80" />
                    <SPLIT distance="400" swimtime="00:05:11.81" />
                    <SPLIT distance="450" swimtime="00:05:50.99" />
                    <SPLIT distance="500" swimtime="00:06:30.15" />
                    <SPLIT distance="550" swimtime="00:07:09.51" />
                    <SPLIT distance="600" swimtime="00:07:48.85" />
                    <SPLIT distance="650" swimtime="00:08:27.70" />
                    <SPLIT distance="700" swimtime="00:09:06.43" />
                    <SPLIT distance="750" swimtime="00:09:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="641" reactiontime="+80" swimtime="00:01:05.07" resultid="7614" heatid="11466" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="643" reactiontime="+94" swimtime="00:02:39.71" resultid="7615" heatid="11499" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="602" reactiontime="+86" swimtime="00:00:32.67" resultid="7616" heatid="11527" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="6518" points="727" reactiontime="+86" swimtime="00:02:19.02" resultid="7617" heatid="11559" lane="3" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="631" swimtime="00:01:11.11" resultid="7618" heatid="11588" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="725" reactiontime="+93" swimtime="00:04:58.06" resultid="7619" heatid="11628" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                    <SPLIT distance="200" swimtime="00:02:27.34" />
                    <SPLIT distance="250" swimtime="00:03:05.50" />
                    <SPLIT distance="300" swimtime="00:03:43.76" />
                    <SPLIT distance="350" swimtime="00:04:21.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" swrid="4762175" athleteid="7594">
              <RESULTS>
                <RESULT eventid="6077" points="811" swimtime="00:00:24.49" resultid="7595" heatid="11418" lane="1" entrytime="00:00:24.50" />
                <RESULT eventid="6169" points="718" reactiontime="+78" swimtime="00:09:30.74" resultid="7596" heatid="11645" lane="6" entrytime="00:09:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:42.34" />
                    <SPLIT distance="200" swimtime="00:02:18.46" />
                    <SPLIT distance="250" swimtime="00:02:54.72" />
                    <SPLIT distance="300" swimtime="00:03:30.72" />
                    <SPLIT distance="350" swimtime="00:04:07.54" />
                    <SPLIT distance="400" swimtime="00:04:44.64" />
                    <SPLIT distance="450" swimtime="00:05:21.03" />
                    <SPLIT distance="500" swimtime="00:05:57.98" />
                    <SPLIT distance="550" swimtime="00:06:34.18" />
                    <SPLIT distance="600" swimtime="00:07:10.49" />
                    <SPLIT distance="650" swimtime="00:07:46.79" />
                    <SPLIT distance="700" swimtime="00:08:22.31" />
                    <SPLIT distance="750" swimtime="00:08:57.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="705" reactiontime="+69" swimtime="00:00:54.57" resultid="7597" heatid="11479" lane="0" entrytime="00:00:54.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="636" reactiontime="+71" swimtime="00:01:04.18" resultid="7598" heatid="11496" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="720" swimtime="00:00:26.44" resultid="7599" heatid="11542" lane="9" entrytime="00:00:26.02" />
                <RESULT eventid="6535" points="741" reactiontime="+75" swimtime="00:02:02.83" resultid="7600" heatid="11571" lane="0" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="737" swimtime="00:00:59.69" resultid="7601" heatid="11597" lane="9" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="747" reactiontime="+73" swimtime="00:04:26.91" resultid="7602" heatid="11637" lane="8" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:38.86" />
                    <SPLIT distance="200" swimtime="00:02:13.97" />
                    <SPLIT distance="250" swimtime="00:02:48.05" />
                    <SPLIT distance="300" swimtime="00:03:22.30" />
                    <SPLIT distance="350" swimtime="00:03:55.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" swrid="4602697" athleteid="7603">
              <RESULTS>
                <RESULT eventid="6059" points="805" reactiontime="+79" swimtime="00:00:27.18" resultid="7604" heatid="11401" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="6094" points="792" reactiontime="+78" swimtime="00:02:32.37" resultid="7605" heatid="11424" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="814" reactiontime="+79" swimtime="00:01:00.09" resultid="7606" heatid="11466" lane="3" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="777" reactiontime="+78" swimtime="00:01:09.36" resultid="7607" heatid="11486" lane="6" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="761" swimtime="00:00:30.22" resultid="7608" heatid="11528" lane="8" entrytime="00:00:30.80" />
                <RESULT eventid="6618" points="707" reactiontime="+80" swimtime="00:01:08.46" resultid="7609" heatid="11588" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="627" reactiontime="+79" swimtime="00:00:36.89" resultid="7610" heatid="11612" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" swrid="5502059" athleteid="7620">
              <RESULTS>
                <RESULT eventid="6077" points="611" reactiontime="+67" swimtime="00:00:26.91" resultid="7621" heatid="11414" lane="8" entrytime="00:00:27.73" />
                <RESULT eventid="6169" reactiontime="+65" status="OTL" swimtime="00:00:00.00" resultid="7622" heatid="11645" lane="0" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                    <SPLIT distance="200" swimtime="00:02:31.24" />
                    <SPLIT distance="250" swimtime="00:03:10.76" />
                    <SPLIT distance="300" swimtime="00:03:50.84" />
                    <SPLIT distance="350" swimtime="00:04:31.45" />
                    <SPLIT distance="400" swimtime="00:05:12.58" />
                    <SPLIT distance="450" swimtime="00:05:53.70" />
                    <SPLIT distance="500" swimtime="00:06:36.94" />
                    <SPLIT distance="550" swimtime="00:07:20.16" />
                    <SPLIT distance="600" swimtime="00:08:02.68" />
                    <SPLIT distance="650" swimtime="00:08:44.27" />
                    <SPLIT distance="700" swimtime="00:09:26.22" />
                    <SPLIT distance="750" swimtime="00:10:07.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="512" reactiontime="+65" swimtime="00:01:00.69" resultid="7623" heatid="11475" lane="3" entrytime="00:01:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="487" swimtime="00:01:10.14" resultid="7624" heatid="11494" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="443" reactiontime="+63" swimtime="00:00:31.08" resultid="7625" heatid="11536" lane="6" entrytime="00:00:31.90" />
                <RESULT eventid="6535" points="520" reactiontime="+67" swimtime="00:02:18.20" resultid="7626" heatid="11568" lane="9" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="512" reactiontime="+65" swimtime="00:00:35.32" resultid="7627" heatid="11620" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="6738" points="490" reactiontime="+70" swimtime="00:05:07.14" resultid="7628" heatid="11636" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                    <SPLIT distance="200" swimtime="00:02:30.25" />
                    <SPLIT distance="250" swimtime="00:03:10.83" />
                    <SPLIT distance="300" swimtime="00:03:50.77" />
                    <SPLIT distance="350" swimtime="00:04:30.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+82" swimtime="00:01:48.19" resultid="9864" heatid="11436" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                    <SPLIT distance="100" swimtime="00:00:53.97" />
                    <SPLIT distance="150" swimtime="00:01:18.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7603" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="7620" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="7594" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="7611" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+65" swimtime="00:02:04.44" resultid="9865" heatid="11507" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:34.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7603" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="7620" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="7594" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="7611" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8586" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mikołaj" lastname="Konieczny" birthdate="1998-01-01" gender="M" nation="POL" athleteid="8585">
              <RESULTS>
                <RESULT eventid="6340" points="247" reactiontime="+67" swimtime="00:01:29.53" resultid="8587" heatid="11487" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="276" swimtime="00:00:37.75" resultid="8588" heatid="11530" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REKIN" nation="POL" clubid="6797" name="Szkoła pływania REKIN - Koszalin">
          <ATHLETES>
            <ATHLETE firstname="Artem" lastname="Ospishchev" birthdate="1997-09-18" gender="M" nation="POL" athleteid="6798">
              <RESULTS>
                <RESULT eventid="6077" points="667" reactiontime="+74" swimtime="00:00:26.13" resultid="6799" heatid="11415" lane="7" entrytime="00:00:26.90" />
                <RESULT eventid="6306" points="546" reactiontime="+69" swimtime="00:00:59.41" resultid="7318" heatid="11476" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7319" heatid="11538" lane="0" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6950" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kęsik" birthdate="1979-01-01" gender="M" nation="POL" athleteid="6949">
              <RESULTS>
                <RESULT eventid="6077" points="700" swimtime="00:00:26.13" resultid="6951" heatid="11414" lane="4" entrytime="00:00:27.10" />
                <RESULT eventid="6111" points="621" swimtime="00:02:29.87" resultid="6952" heatid="11433" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="669" reactiontime="+75" swimtime="00:00:58.60" resultid="6953" heatid="11477" lane="8" entrytime="00:00:59.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="744" reactiontime="+79" swimtime="00:01:05.99" resultid="6954" heatid="11496" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="722" reactiontime="+75" swimtime="00:00:28.00" resultid="6955" heatid="11539" lane="6" entrytime="00:00:28.90" />
                <RESULT eventid="6535" points="584" reactiontime="+81" swimtime="00:02:15.15" resultid="6956" heatid="11570" lane="8" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="719" reactiontime="+91" swimtime="00:01:03.19" resultid="6957" heatid="11595" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="571" reactiontime="+101" swimtime="00:04:49.96" resultid="6958" heatid="11636" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:44.18" />
                    <SPLIT distance="200" swimtime="00:02:21.37" />
                    <SPLIT distance="250" swimtime="00:02:58.99" />
                    <SPLIT distance="300" swimtime="00:03:36.75" />
                    <SPLIT distance="350" swimtime="00:04:14.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="6980" name="ŠPK Kupele Piešťany">
          <ATHLETES>
            <ATHLETE firstname="Pavel" lastname="Škodný" birthdate="1969-01-01" gender="M" nation="SVK" swrid="4688816" athleteid="6991">
              <RESULTS>
                <RESULT eventid="6111" points="590" reactiontime="+85" swimtime="00:02:37.32" resultid="6992" heatid="11431" lane="2" entrytime="00:02:38.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:15.40" />
                    <SPLIT distance="150" swimtime="00:02:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="560" reactiontime="+81" swimtime="00:00:34.39" resultid="6993" heatid="11447" lane="4" entrytime="00:00:34.33" entrycourse="SCM" />
                <RESULT eventid="6501" points="550" reactiontime="+88" swimtime="00:01:13.81" resultid="6994" heatid="11552" lane="9" entrytime="00:01:13.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="663" reactiontime="+91" swimtime="00:05:43.36" resultid="6995" heatid="11578" lane="3" entrytime="00:05:39.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                    <SPLIT distance="200" swimtime="00:02:45.89" />
                    <SPLIT distance="250" swimtime="00:03:35.28" />
                    <SPLIT distance="300" swimtime="00:04:24.91" />
                    <SPLIT distance="350" swimtime="00:05:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="656" reactiontime="+93" swimtime="00:02:40.09" resultid="6996" heatid="11605" lane="7" entrytime="00:02:39.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juraj" lastname="Horil" birthdate="1972-01-01" gender="M" nation="SVK" swrid="4928173" athleteid="6997">
              <RESULTS>
                <RESULT eventid="6077" points="469" reactiontime="+82" swimtime="00:00:31.50" resultid="6998" heatid="11410" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="6272" points="569" reactiontime="+73" swimtime="00:03:06.70" resultid="6999" heatid="11458" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:26.35" />
                    <SPLIT distance="150" swimtime="00:02:16.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="543" reactiontime="+77" swimtime="00:01:22.28" resultid="7000" heatid="11518" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="382" reactiontime="+90" swimtime="00:02:42.65" resultid="7001" heatid="11566" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:58.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="590" reactiontime="+75" swimtime="00:00:36.67" resultid="7002" heatid="11619" lane="3" entrytime="00:00:37.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzana" lastname="Matúšová" birthdate="1982-01-01" gender="F" nation="SVK" swrid="4270447" athleteid="7003">
              <RESULTS>
                <RESULT eventid="6094" points="720" swimtime="00:02:43.73" resultid="7004" heatid="11424" lane="9" entrytime="00:02:46.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="758" swimtime="00:01:14.72" resultid="7005" heatid="11485" lane="4" entrytime="00:01:15.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="785" reactiontime="+83" swimtime="00:01:22.03" resultid="7006" heatid="11512" lane="7" entrytime="00:01:22.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="707" reactiontime="+80" swimtime="00:00:32.89" resultid="7007" heatid="11527" lane="3" entrytime="00:00:32.50" entrycourse="SCM" />
                <RESULT eventid="6618" points="645" reactiontime="+82" swimtime="00:01:14.75" resultid="7008" heatid="11588" lane="1" entrytime="00:01:13.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="821" reactiontime="+77" swimtime="00:00:36.66" resultid="7009" heatid="11612" lane="1" entrytime="00:00:36.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martin" lastname="Babsky" birthdate="1972-01-01" gender="M" nation="SVK" swrid="5439025" athleteid="6986">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="6987" heatid="11415" lane="6" entrytime="00:00:26.51" entrycourse="SCM" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="6988" heatid="11476" lane="4" entrytime="00:00:59.63" entrycourse="SCM" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="6989" heatid="11568" lane="7" entrytime="00:02:18.36" entrycourse="SCM" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="6990" heatid="11593" lane="2" entrytime="00:01:12.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6933" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-01-01" gender="M" nation="POL" athleteid="6932">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="6077" reactiontime="+69" status="DSQ" swimtime="00:00:00.00" resultid="6934" heatid="11409" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="6169" reactiontime="+108" status="OTL" swimtime="00:00:00.00" resultid="6935" heatid="11647" lane="3" entrytime="00:12:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:13.23" />
                    <SPLIT distance="200" swimtime="00:03:02.62" />
                    <SPLIT distance="250" swimtime="00:03:51.64" />
                    <SPLIT distance="300" swimtime="00:04:41.21" />
                    <SPLIT distance="350" swimtime="00:05:30.43" />
                    <SPLIT distance="400" swimtime="00:06:20.01" />
                    <SPLIT distance="450" swimtime="00:07:08.90" />
                    <SPLIT distance="500" swimtime="00:07:58.81" />
                    <SPLIT distance="550" swimtime="00:08:48.52" />
                    <SPLIT distance="600" swimtime="00:09:38.32" />
                    <SPLIT distance="650" swimtime="00:10:27.37" />
                    <SPLIT distance="700" swimtime="00:11:16.17" />
                    <SPLIT distance="750" swimtime="00:12:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="345" reactiontime="+93" swimtime="00:01:15.41" resultid="6936" heatid="11472" lane="0" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="302" reactiontime="+99" swimtime="00:01:29.38" resultid="6937" heatid="11490" lane="2" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="264" reactiontime="+86" swimtime="00:01:32.58" resultid="6938" heatid="11550" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="311" reactiontime="+86" swimtime="00:02:49.19" resultid="6939" heatid="11565" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:03.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M7 - Pływak wykonał naprzemienne lub nierównoczesne ruchy nóg." eventid="6636" reactiontime="+102" status="DSQ" swimtime="00:00:00.00" resultid="6940" heatid="11591" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="292" swimtime="00:06:10.35" resultid="6941" heatid="11633" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:27.90" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                    <SPLIT distance="200" swimtime="00:03:04.62" />
                    <SPLIT distance="250" swimtime="00:03:53.59" />
                    <SPLIT distance="300" swimtime="00:04:41.51" />
                    <SPLIT distance="350" swimtime="00:05:28.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6962" name="Iks Dss Kraków">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" license="505806600021" swrid="5484417" athleteid="6963">
              <RESULTS>
                <RESULT eventid="6059" points="213" reactiontime="+108" swimtime="00:00:53.97" resultid="6964" heatid="11396" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="6094" points="213" reactiontime="+127" swimtime="00:05:05.66" resultid="6965" heatid="11421" lane="8" entrytime="00:05:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.31" />
                    <SPLIT distance="100" swimtime="00:02:33.42" />
                    <SPLIT distance="150" swimtime="00:03:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="269" reactiontime="+72" swimtime="00:01:02.00" resultid="6966" heatid="11439" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="6289" points="198" swimtime="00:02:01.60" resultid="6967" heatid="11462" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="118" swimtime="00:01:12.12" resultid="6968" heatid="11524" lane="0" entrytime="00:01:16.00" />
                <RESULT eventid="6484" points="264" reactiontime="+79" swimtime="00:02:16.43" resultid="6969" heatid="11544" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="270" reactiontime="+79" swimtime="00:04:51.35" resultid="6970" heatid="11599" lane="8" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.31" />
                    <SPLIT distance="100" swimtime="00:02:24.19" />
                    <SPLIT distance="150" swimtime="00:03:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="276" swimtime="00:09:01.12" resultid="6971" heatid="11625" lane="8" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.56" />
                    <SPLIT distance="100" swimtime="00:02:07.16" />
                    <SPLIT distance="150" swimtime="00:03:15.40" />
                    <SPLIT distance="200" swimtime="00:04:24.63" />
                    <SPLIT distance="250" swimtime="00:05:35.47" />
                    <SPLIT distance="300" swimtime="00:06:45.15" />
                    <SPLIT distance="350" swimtime="00:07:53.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00701" nation="POL" region="01" clubid="9191" name="MKS Dziewiątka Dzierżoniów">
          <ATHLETES>
            <ATHLETE firstname="Edyta" lastname="Bejster" birthdate="1981-05-21" gender="F" nation="POL" license="100701600124" swrid="5464069" athleteid="9200">
              <RESULTS>
                <RESULT eventid="6059" points="324" reactiontime="+102" swimtime="00:00:38.26" resultid="9201" heatid="11395" lane="2" />
                <RESULT eventid="6220" points="197" reactiontime="+81" swimtime="00:00:52.48" resultid="9202" heatid="11438" lane="5" />
                <RESULT eventid="6323" points="298" swimtime="00:01:41.96" resultid="9203" heatid="11482" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="373" swimtime="00:01:45.06" resultid="9204" heatid="11509" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M9 - Pływak wykonał więcej niż jeden ruch nóg do stylu klasycznego w trakcie jednego cyklu ruchowego (dotyczy pływania Masters)." eventid="6450" reactiontime="+102" status="DSQ" swimtime="00:00:00.00" resultid="9205" heatid="11523" lane="1" />
                <RESULT eventid="6687" points="399" reactiontime="+94" swimtime="00:00:46.63" resultid="9206" heatid="11608" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kuszka" birthdate="1977-04-14" gender="M" nation="POL" license="100701700110" athleteid="9207">
              <RESULTS>
                <RESULT eventid="6077" points="311" swimtime="00:00:35.21" resultid="9208" heatid="11403" lane="6" />
                <RESULT eventid="6111" points="242" swimtime="00:03:32.24" resultid="9209" heatid="11426" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:41.59" />
                    <SPLIT distance="150" swimtime="00:02:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="307" reactiontime="+79" swimtime="00:03:38.73" resultid="9210" heatid="11455" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="150" swimtime="00:02:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="274" reactiontime="+78" swimtime="00:01:32.31" resultid="9211" heatid="11488" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="310" reactiontime="+82" swimtime="00:01:37.60" resultid="9212" heatid="11514" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="285" reactiontime="+77" swimtime="00:00:39.01" resultid="9213" heatid="11530" lane="1" />
                <RESULT eventid="6636" points="205" reactiontime="+82" swimtime="00:01:39.21" resultid="9214" heatid="11589" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="393" reactiontime="+78" swimtime="00:00:41.35" resultid="9215" heatid="11615" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Pisarska" birthdate="1981-11-06" gender="F" nation="POL" license="100701600113" swrid="5464072" athleteid="9192">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6059" points="884" reactiontime="+65" swimtime="00:00:27.38" resultid="9193" heatid="11394" lane="6" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6094" points="853" swimtime="00:02:34.74" resultid="9194" heatid="11420" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6220" points="948" reactiontime="+65" swimtime="00:00:31.09" resultid="9195" heatid="11438" lane="9" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6323" points="964" reactiontime="+75" swimtime="00:01:08.96" resultid="9196" heatid="11480" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6450" points="1021" reactiontime="+66" swimtime="00:00:29.09" resultid="9197" heatid="11523" lane="4" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6484" points="993" reactiontime="+68" swimtime="00:01:08.10" resultid="9198" heatid="11544" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6618" points="873" reactiontime="+70" swimtime="00:01:07.59" resultid="9199" heatid="11585" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="9232" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" license="102805600154" athleteid="9399">
              <RESULTS>
                <RESULT eventid="6289" points="382" reactiontime="+100" swimtime="00:01:20.55" resultid="9400" heatid="11463" lane="8" entrytime="00:01:27.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="307" reactiontime="+89" swimtime="00:00:43.42" resultid="9401" heatid="11524" lane="3" entrytime="00:00:48.01" />
                <RESULT eventid="6518" points="401" reactiontime="+97" swimtime="00:02:55.24" resultid="9402" heatid="11557" lane="2" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:24.29" />
                    <SPLIT distance="150" swimtime="00:02:11.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="398" reactiontime="+90" swimtime="00:06:16.30" resultid="9403" heatid="11625" lane="6" entrytime="00:07:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                    <SPLIT distance="150" swimtime="00:02:16.03" />
                    <SPLIT distance="200" swimtime="00:03:05.98" />
                    <SPLIT distance="250" swimtime="00:03:53.65" />
                    <SPLIT distance="300" swimtime="00:04:43.39" />
                    <SPLIT distance="350" swimtime="00:05:31.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Sikorski" birthdate="1951-05-03" gender="M" nation="POL" license="502805700036" athleteid="9385">
              <RESULTS>
                <RESULT eventid="6238" points="217" reactiontime="+91" swimtime="00:00:57.65" resultid="9386" heatid="11444" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="6433" points="293" reactiontime="+92" swimtime="00:02:04.07" resultid="9387" heatid="11515" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="202" reactiontime="+94" swimtime="00:02:07.81" resultid="9388" heatid="11549" lane="9" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="300" reactiontime="+87" swimtime="00:00:53.03" resultid="9389" heatid="11616" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Maciejewski" birthdate="1974-04-11" gender="M" nation="POL" license="502805700028" swrid="5373991" athleteid="9312">
              <RESULTS>
                <RESULT eventid="6077" points="314" reactiontime="+94" swimtime="00:00:35.10" resultid="9313" heatid="11405" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="6169" reactiontime="+95" status="OTL" swimtime="00:00:00.00" resultid="9314" heatid="11648" lane="5" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:27.07" />
                    <SPLIT distance="150" swimtime="00:02:16.47" />
                    <SPLIT distance="200" swimtime="00:03:07.26" />
                    <SPLIT distance="250" swimtime="00:04:00.56" />
                    <SPLIT distance="300" swimtime="00:04:54.63" />
                    <SPLIT distance="350" swimtime="00:05:48.73" />
                    <SPLIT distance="400" swimtime="00:06:46.92" />
                    <SPLIT distance="450" swimtime="00:07:45.91" />
                    <SPLIT distance="500" swimtime="00:08:42.58" />
                    <SPLIT distance="550" swimtime="00:09:38.59" />
                    <SPLIT distance="600" swimtime="00:10:34.73" />
                    <SPLIT distance="650" swimtime="00:11:33.78" />
                    <SPLIT distance="700" swimtime="00:12:28.94" />
                    <SPLIT distance="750" swimtime="00:13:25.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="293" reactiontime="+89" swimtime="00:01:19.64" resultid="9315" heatid="11470" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="276" reactiontime="+98" swimtime="00:01:41.45" resultid="9316" heatid="11517" lane="1" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="326" reactiontime="+92" swimtime="00:00:44.00" resultid="9317" heatid="11616" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Dziarek" birthdate="1959-02-19" gender="M" nation="POL" license="502805700029" swrid="4841500" athleteid="9372">
              <RESULTS>
                <RESULT eventid="6203" points="566" reactiontime="+99" swimtime="00:23:40.65" resultid="9373" heatid="11653" lane="6" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:25.61" />
                    <SPLIT distance="150" swimtime="00:02:11.76" />
                    <SPLIT distance="200" swimtime="00:02:59.25" />
                    <SPLIT distance="250" swimtime="00:03:47.01" />
                    <SPLIT distance="300" swimtime="00:04:34.35" />
                    <SPLIT distance="350" swimtime="00:05:21.91" />
                    <SPLIT distance="400" swimtime="00:06:09.52" />
                    <SPLIT distance="450" swimtime="00:06:56.81" />
                    <SPLIT distance="500" swimtime="00:07:44.40" />
                    <SPLIT distance="550" swimtime="00:08:32.00" />
                    <SPLIT distance="600" swimtime="00:09:19.73" />
                    <SPLIT distance="650" swimtime="00:10:07.18" />
                    <SPLIT distance="700" swimtime="00:10:54.10" />
                    <SPLIT distance="750" swimtime="00:11:40.85" />
                    <SPLIT distance="800" swimtime="00:12:28.56" />
                    <SPLIT distance="850" swimtime="00:13:16.05" />
                    <SPLIT distance="900" swimtime="00:14:04.51" />
                    <SPLIT distance="950" swimtime="00:14:52.08" />
                    <SPLIT distance="1000" swimtime="00:15:40.06" />
                    <SPLIT distance="1050" swimtime="00:16:27.68" />
                    <SPLIT distance="1100" swimtime="00:17:15.20" />
                    <SPLIT distance="1150" swimtime="00:18:03.12" />
                    <SPLIT distance="1200" swimtime="00:18:51.20" />
                    <SPLIT distance="1250" swimtime="00:19:39.36" />
                    <SPLIT distance="1300" swimtime="00:20:27.41" />
                    <SPLIT distance="1350" swimtime="00:21:15.51" />
                    <SPLIT distance="1400" swimtime="00:22:03.87" />
                    <SPLIT distance="1450" swimtime="00:22:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="9374" heatid="11471" lane="9" entrytime="00:01:18.00" />
                <RESULT eventid="6535" points="571" reactiontime="+94" swimtime="00:02:44.45" resultid="9375" heatid="11564" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:02:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="561" reactiontime="+111" swimtime="00:05:53.03" resultid="9376" heatid="11635" lane="9" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                    <SPLIT distance="200" swimtime="00:02:52.11" />
                    <SPLIT distance="250" swimtime="00:03:38.00" />
                    <SPLIT distance="300" swimtime="00:04:23.60" />
                    <SPLIT distance="350" swimtime="00:05:09.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="9233">
              <RESULTS>
                <RESULT eventid="6059" points="310" reactiontime="+69" swimtime="00:00:39.75" resultid="9234" heatid="11397" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="6094" points="318" reactiontime="+71" swimtime="00:03:39.79" resultid="9235" heatid="11421" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.12" />
                    <SPLIT distance="100" swimtime="00:01:48.47" />
                    <SPLIT distance="150" swimtime="00:02:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="459" swimtime="00:03:39.36" resultid="9236" heatid="11453" lane="2" entrytime="00:03:36.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.16" />
                    <SPLIT distance="100" swimtime="00:01:45.52" />
                    <SPLIT distance="150" swimtime="00:02:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="313" swimtime="00:01:41.76" resultid="9237" heatid="11483" lane="0" entrytime="00:01:39.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="437" swimtime="00:01:42.16" resultid="9238" heatid="11511" lane="8" entrytime="00:01:39.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="261" reactiontime="+84" swimtime="00:01:46.10" resultid="9239" heatid="11545" lane="8" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="274" reactiontime="+88" swimtime="00:03:56.72" resultid="9240" heatid="11599" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.66" />
                    <SPLIT distance="100" swimtime="00:01:57.49" />
                    <SPLIT distance="150" swimtime="00:02:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="432" reactiontime="+68" swimtime="00:00:45.98" resultid="9241" heatid="11611" lane="9" entrytime="00:00:45.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="9321">
              <RESULTS>
                <RESULT eventid="6077" points="631" reactiontime="+80" swimtime="00:00:32.15" resultid="9322" heatid="11410" lane="0" entrytime="00:00:31.50" />
                <RESULT eventid="6111" points="657" reactiontime="+88" swimtime="00:03:02.39" resultid="9323" heatid="11429" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                    <SPLIT distance="150" swimtime="00:02:22.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="9324" heatid="11446" lane="3" entrytime="00:00:39.37" entrycourse="SCM" />
                <RESULT eventid="6374" status="DNS" swimtime="00:00:00.00" resultid="9325" heatid="11502" lane="3" entrytime="00:03:12.47" entrycourse="SCM" />
                <RESULT eventid="6467" points="743" reactiontime="+85" swimtime="00:00:33.73" resultid="9326" heatid="11535" lane="6" entrytime="00:00:33.46" entrycourse="SCM" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="9327" heatid="11565" lane="9" entrytime="00:02:52.00" />
                <RESULT eventid="6636" points="553" reactiontime="+90" swimtime="00:01:26.78" resultid="9328" heatid="11592" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9329" heatid="11633" lane="7" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="9248">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6059" points="807" reactiontime="+90" swimtime="00:00:33.30" resultid="9249" heatid="11398" lane="9" entrytime="00:00:34.73" entrycourse="SCM" />
                <RESULT eventid="6220" points="719" reactiontime="+83" swimtime="00:00:40.53" resultid="9250" heatid="11440" lane="9" entrytime="00:00:43.51" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6323" points="815" reactiontime="+87" swimtime="00:01:24.66" resultid="9251" heatid="11484" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6450" points="835" reactiontime="+93" swimtime="00:00:35.50" resultid="9252" heatid="11526" lane="9" entrytime="00:00:36.62" entrycourse="SCM" />
                <RESULT eventid="6484" points="686" reactiontime="+85" swimtime="00:01:31.93" resultid="9253" heatid="11545" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6618" points="860" reactiontime="+89" swimtime="00:01:25.62" resultid="9254" heatid="11587" lane="1" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="642" swimtime="00:00:44.17" resultid="9255" heatid="11610" lane="4" entrytime="00:00:45.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" license="102805700157" swrid="4071609" athleteid="9351">
              <RESULTS>
                <RESULT eventid="6111" points="724" reactiontime="+78" swimtime="00:02:11.54" resultid="9352" heatid="11433" lane="7" entrytime="00:02:22.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                    <SPLIT distance="100" swimtime="00:01:01.23" />
                    <SPLIT distance="150" swimtime="00:01:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="970" reactiontime="+73" swimtime="00:02:21.93" resultid="9353" heatid="11460" lane="3" entrytime="00:02:24.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:08.66" />
                    <SPLIT distance="150" swimtime="00:01:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="721" reactiontime="+73" swimtime="00:01:01.32" resultid="9354" heatid="11497" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="869" reactiontime="+72" swimtime="00:01:04.27" resultid="9355" heatid="11521" lane="2" entrytime="00:01:05.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="784" reactiontime="+73" swimtime="00:04:49.54" resultid="9356" heatid="11579" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                    <SPLIT distance="200" swimtime="00:02:25.04" />
                    <SPLIT distance="250" swimtime="00:03:04.01" />
                    <SPLIT distance="300" swimtime="00:03:43.45" />
                    <SPLIT distance="350" swimtime="00:04:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="815" swimtime="00:00:29.77" resultid="9357" heatid="11623" lane="0" entrytime="00:00:30.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="9390">
              <RESULTS>
                <RESULT eventid="6272" points="334" reactiontime="+95" swimtime="00:03:59.07" resultid="9391" heatid="11456" lane="6" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.59" />
                    <SPLIT distance="100" swimtime="00:01:56.31" />
                    <SPLIT distance="150" swimtime="00:03:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="382" reactiontime="+92" swimtime="00:01:41.78" resultid="9392" heatid="11516" lane="1" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="431" reactiontime="+138" swimtime="00:00:43.34" resultid="9393" heatid="11617" lane="7" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="9272">
              <RESULTS>
                <RESULT eventid="6059" points="801" swimtime="00:00:30.46" resultid="9273" heatid="11399" lane="9" entrytime="00:00:32.88" entrycourse="SCM" />
                <RESULT eventid="6094" points="839" reactiontime="+82" swimtime="00:02:42.54" resultid="9274" heatid="11423" lane="5" entrytime="00:02:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:02:03.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="624" reactiontime="+79" swimtime="00:00:36.62" resultid="9275" heatid="11441" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="6323" points="791" reactiontime="+79" swimtime="00:01:14.67" resultid="9276" heatid="11485" lane="3" entrytime="00:01:16.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="898" reactiontime="+74" swimtime="00:00:32.28" resultid="9277" heatid="11527" lane="6" entrytime="00:00:32.52" entrycourse="SCM" />
                <RESULT eventid="6618" points="750" reactiontime="+85" swimtime="00:01:14.41" resultid="9278" heatid="11588" lane="2" entrytime="00:01:12.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Kaczmarek" birthdate="1976-11-27" gender="F" nation="POL" license="502805600149" athleteid="9242">
              <RESULTS>
                <RESULT eventid="6059" points="152" reactiontime="+65" swimtime="00:00:50.39" resultid="9243" heatid="11396" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="6255" points="211" reactiontime="+85" swimtime="00:04:43.99" resultid="9244" heatid="11452" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.22" />
                    <SPLIT distance="100" swimtime="00:02:14.35" />
                    <SPLIT distance="150" swimtime="00:03:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="114" reactiontime="+79" swimtime="00:02:02.83" resultid="9245" heatid="11462" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="172" swimtime="00:02:19.40" resultid="9246" heatid="11510" lane="1" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="170" reactiontime="+73" swimtime="00:01:02.72" resultid="9247" heatid="11610" lane="2" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="9377">
              <RESULTS>
                <RESULT eventid="6203" points="324" reactiontime="+107" swimtime="00:23:58.86" resultid="9378" heatid="11653" lane="5" entrytime="00:24:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:08.04" />
                    <SPLIT distance="200" swimtime="00:02:54.52" />
                    <SPLIT distance="250" swimtime="00:03:42.51" />
                    <SPLIT distance="300" swimtime="00:04:30.12" />
                    <SPLIT distance="350" swimtime="00:05:19.25" />
                    <SPLIT distance="400" swimtime="00:06:07.32" />
                    <SPLIT distance="450" swimtime="00:06:55.74" />
                    <SPLIT distance="500" swimtime="00:07:44.78" />
                    <SPLIT distance="550" swimtime="00:08:33.14" />
                    <SPLIT distance="600" swimtime="00:09:22.01" />
                    <SPLIT distance="650" swimtime="00:10:10.49" />
                    <SPLIT distance="700" swimtime="00:10:59.27" />
                    <SPLIT distance="750" swimtime="00:11:48.22" />
                    <SPLIT distance="800" swimtime="00:12:37.16" />
                    <SPLIT distance="850" swimtime="00:13:25.98" />
                    <SPLIT distance="900" swimtime="00:14:14.55" />
                    <SPLIT distance="950" swimtime="00:15:03.41" />
                    <SPLIT distance="1000" swimtime="00:15:52.89" />
                    <SPLIT distance="1050" swimtime="00:16:41.64" />
                    <SPLIT distance="1100" swimtime="00:17:31.04" />
                    <SPLIT distance="1150" swimtime="00:18:19.75" />
                    <SPLIT distance="1200" swimtime="00:19:08.28" />
                    <SPLIT distance="1250" swimtime="00:19:57.35" />
                    <SPLIT distance="1300" swimtime="00:20:46.50" />
                    <SPLIT distance="1350" swimtime="00:21:35.60" />
                    <SPLIT distance="1400" swimtime="00:22:23.84" />
                    <SPLIT distance="1450" swimtime="00:23:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="334" reactiontime="+106" swimtime="00:03:32.63" resultid="9379" heatid="11457" lane="7" entrytime="00:03:27.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:39.10" />
                    <SPLIT distance="150" swimtime="00:02:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="310" swimtime="00:01:28.60" resultid="9380" heatid="11490" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="9381" heatid="11549" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="6569" points="275" reactiontime="+107" swimtime="00:07:24.42" resultid="9382" heatid="11577" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:43.07" />
                    <SPLIT distance="150" swimtime="00:02:43.69" />
                    <SPLIT distance="200" swimtime="00:03:44.07" />
                    <SPLIT distance="250" swimtime="00:04:44.21" />
                    <SPLIT distance="300" swimtime="00:05:44.50" />
                    <SPLIT distance="350" swimtime="00:06:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="433" reactiontime="+96" swimtime="00:00:40.01" resultid="9383" heatid="11618" lane="5" entrytime="00:00:39.30" entrycourse="SCM" />
                <RESULT eventid="6738" points="317" reactiontime="+98" swimtime="00:06:00.40" resultid="9384" heatid="11632" lane="3" entrytime="00:06:10.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:20.51" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                    <SPLIT distance="200" swimtime="00:02:54.31" />
                    <SPLIT distance="250" swimtime="00:03:42.72" />
                    <SPLIT distance="300" swimtime="00:04:30.15" />
                    <SPLIT distance="350" swimtime="00:05:16.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" swrid="5464095" athleteid="9265">
              <RESULTS>
                <RESULT eventid="6059" points="285" swimtime="00:00:40.86" resultid="9266" heatid="11397" lane="9" entrytime="00:00:41.10" entrycourse="SCM" />
                <RESULT eventid="6255" points="234" swimtime="00:04:34.67" resultid="9267" heatid="11453" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.31" />
                    <SPLIT distance="100" swimtime="00:02:08.32" />
                    <SPLIT distance="150" swimtime="00:03:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="226" swimtime="00:01:37.77" resultid="9268" heatid="11463" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="256" swimtime="00:02:01.96" resultid="9269" heatid="11511" lane="1" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="194" reactiontime="+92" swimtime="00:03:45.29" resultid="9270" heatid="11556" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.41" />
                    <SPLIT distance="100" swimtime="00:01:46.12" />
                    <SPLIT distance="150" swimtime="00:02:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="285" reactiontime="+91" swimtime="00:00:52.81" resultid="9271" heatid="11610" lane="7" entrytime="00:00:51.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="9358">
              <RESULTS>
                <RESULT eventid="6169" points="424" reactiontime="+100" swimtime="00:15:15.31" resultid="9359" heatid="11648" lane="6" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.28" />
                    <SPLIT distance="100" swimtime="00:01:45.98" />
                    <SPLIT distance="150" swimtime="00:02:45.30" />
                    <SPLIT distance="200" swimtime="00:03:44.52" />
                    <SPLIT distance="250" swimtime="00:04:43.50" />
                    <SPLIT distance="300" swimtime="00:05:42.01" />
                    <SPLIT distance="350" swimtime="00:06:39.90" />
                    <SPLIT distance="400" swimtime="00:07:37.31" />
                    <SPLIT distance="450" swimtime="00:08:35.38" />
                    <SPLIT distance="500" swimtime="00:09:33.21" />
                    <SPLIT distance="550" swimtime="00:10:31.47" />
                    <SPLIT distance="600" swimtime="00:11:29.89" />
                    <SPLIT distance="650" swimtime="00:12:28.75" />
                    <SPLIT distance="700" swimtime="00:13:25.87" />
                    <SPLIT distance="750" swimtime="00:14:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="615" reactiontime="+103" swimtime="00:03:37.80" resultid="9360" heatid="11457" lane="9" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:45.28" />
                    <SPLIT distance="150" swimtime="00:02:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="606" reactiontime="+101" swimtime="00:01:37.40" resultid="9361" heatid="11517" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="587" reactiontime="+81" swimtime="00:03:37.26" resultid="9362" heatid="11603" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:46.92" />
                    <SPLIT distance="150" swimtime="00:02:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="525" reactiontime="+108" swimtime="00:00:44.02" resultid="9363" heatid="11617" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Jagiełło" birthdate="1979-03-01" gender="M" nation="POL" license="502805700042" swrid="4541616" athleteid="9295">
              <RESULTS>
                <RESULT eventid="6077" points="653" reactiontime="+77" swimtime="00:00:26.74" resultid="9296" heatid="11413" lane="0" entrytime="00:00:28.10" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="9297" heatid="11430" lane="3" entrytime="00:02:44.44" />
                <RESULT eventid="6306" points="596" reactiontime="+83" swimtime="00:01:00.92" resultid="9298" heatid="11476" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="667" reactiontime="+86" swimtime="00:01:08.46" resultid="9299" heatid="11495" lane="5" entrytime="00:01:06.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="664" reactiontime="+79" swimtime="00:01:12.88" resultid="9300" heatid="11520" lane="0" entrytime="00:01:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="575" reactiontime="+82" swimtime="00:00:30.22" resultid="9301" heatid="11537" lane="6" entrytime="00:00:30.30" />
                <RESULT eventid="6704" points="700" swimtime="00:00:32.74" resultid="9302" heatid="11621" lane="0" entrytime="00:00:34.80" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9303" heatid="11635" lane="0" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600152" swrid="5464091" athleteid="9342">
              <RESULTS>
                <RESULT eventid="6094" points="304" reactiontime="+104" swimtime="00:03:43.22" resultid="9343" heatid="11421" lane="3" entrytime="00:03:39.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="100" swimtime="00:01:54.06" />
                    <SPLIT distance="150" swimtime="00:02:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="417" reactiontime="+110" swimtime="00:25:58.74" resultid="9344" heatid="11651" lane="3" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:38.56" />
                    <SPLIT distance="150" swimtime="00:02:31.07" />
                    <SPLIT distance="200" swimtime="00:03:23.36" />
                    <SPLIT distance="250" swimtime="00:04:16.22" />
                    <SPLIT distance="300" swimtime="00:05:09.12" />
                    <SPLIT distance="350" swimtime="00:06:02.97" />
                    <SPLIT distance="400" swimtime="00:06:57.04" />
                    <SPLIT distance="450" swimtime="00:07:50.95" />
                    <SPLIT distance="500" swimtime="00:08:44.82" />
                    <SPLIT distance="550" swimtime="00:09:39.09" />
                    <SPLIT distance="600" swimtime="00:10:33.36" />
                    <SPLIT distance="650" swimtime="00:11:27.91" />
                    <SPLIT distance="700" swimtime="00:12:22.91" />
                    <SPLIT distance="750" swimtime="00:13:16.95" />
                    <SPLIT distance="800" swimtime="00:14:11.37" />
                    <SPLIT distance="850" swimtime="00:15:04.74" />
                    <SPLIT distance="900" swimtime="00:15:59.34" />
                    <SPLIT distance="950" swimtime="00:16:55.08" />
                    <SPLIT distance="1000" swimtime="00:17:50.33" />
                    <SPLIT distance="1050" swimtime="00:18:45.19" />
                    <SPLIT distance="1100" swimtime="00:19:39.81" />
                    <SPLIT distance="1150" swimtime="00:20:34.74" />
                    <SPLIT distance="1200" swimtime="00:21:29.64" />
                    <SPLIT distance="1250" swimtime="00:22:24.86" />
                    <SPLIT distance="1300" swimtime="00:23:19.36" />
                    <SPLIT distance="1350" swimtime="00:24:13.75" />
                    <SPLIT distance="1400" swimtime="00:25:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="387" reactiontime="+122" swimtime="00:03:52.17" resultid="9345" heatid="11453" lane="8" entrytime="00:03:50.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                    <SPLIT distance="100" swimtime="00:01:51.49" />
                    <SPLIT distance="150" swimtime="00:02:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="245" reactiontime="+111" swimtime="00:03:53.88" resultid="9346" heatid="11499" lane="0" entrytime="00:03:55.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                    <SPLIT distance="100" swimtime="00:01:51.62" />
                    <SPLIT distance="150" swimtime="00:02:53.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="293" reactiontime="+112" swimtime="00:03:16.42" resultid="9347" heatid="11556" lane="3" entrytime="00:03:13.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                    <SPLIT distance="150" swimtime="00:02:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="328" reactiontime="+117" swimtime="00:07:48.60" resultid="9348" heatid="11573" lane="7" entrytime="00:08:14.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                    <SPLIT distance="100" swimtime="00:01:50.32" />
                    <SPLIT distance="150" swimtime="00:02:56.49" />
                    <SPLIT distance="200" swimtime="00:04:01.53" />
                    <SPLIT distance="250" swimtime="00:05:03.62" />
                    <SPLIT distance="300" swimtime="00:06:04.94" />
                    <SPLIT distance="350" swimtime="00:06:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="227" reactiontime="+143" swimtime="00:04:11.71" resultid="9349" heatid="11599" lane="1" entrytime="00:04:08.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.21" />
                    <SPLIT distance="100" swimtime="00:02:06.14" />
                    <SPLIT distance="150" swimtime="00:03:10.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="336" reactiontime="+105" swimtime="00:06:48.21" resultid="9350" heatid="11625" lane="4" entrytime="00:06:42.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:02:27.76" />
                    <SPLIT distance="200" swimtime="00:03:20.80" />
                    <SPLIT distance="250" swimtime="00:04:13.71" />
                    <SPLIT distance="300" swimtime="00:05:06.65" />
                    <SPLIT distance="350" swimtime="00:05:58.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" swrid="5373999" athleteid="9330">
              <RESULTS>
                <RESULT eventid="6077" points="564" reactiontime="+65" swimtime="00:00:33.38" resultid="9331" heatid="11408" lane="6" entrytime="00:00:33.45" />
                <RESULT eventid="6111" points="458" reactiontime="+63" swimtime="00:03:25.78" resultid="9332" heatid="11428" lane="6" entrytime="00:03:26.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:34.43" />
                    <SPLIT distance="150" swimtime="00:02:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="575" reactiontime="+79" swimtime="00:00:40.07" resultid="9333" heatid="11446" lane="7" entrytime="00:00:40.93" />
                <RESULT eventid="6340" points="532" reactiontime="+73" swimtime="00:01:27.31" resultid="9334" heatid="11491" lane="8" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="494" reactiontime="+76" swimtime="00:01:37.30" resultid="9335" heatid="11516" lane="3" entrytime="00:01:41.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="500" reactiontime="+81" swimtime="00:01:31.15" resultid="9336" heatid="11550" lane="2" entrytime="00:01:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700153" swrid="5558378" athleteid="9286">
              <RESULTS>
                <RESULT eventid="6077" points="446" swimtime="00:00:31.24" resultid="9287" heatid="11410" lane="1" entrytime="00:00:31.05" entrycourse="SCM" />
                <RESULT eventid="6111" points="321" reactiontime="+97" swimtime="00:03:13.27" resultid="9288" heatid="11429" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                    <SPLIT distance="150" swimtime="00:02:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="408" reactiontime="+83" swimtime="00:01:11.34" resultid="9289" heatid="11472" lane="6" entrytime="00:01:11.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="386" swimtime="00:01:22.34" resultid="9290" heatid="11491" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="413" reactiontime="+84" swimtime="00:00:34.46" resultid="9291" heatid="11534" lane="6" entrytime="00:00:35.09" entrycourse="SCM" />
                <RESULT eventid="6535" points="346" swimtime="00:02:43.42" resultid="9292" heatid="11565" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9293" heatid="11591" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="6738" points="320" swimtime="00:05:59.30" resultid="9294" heatid="11632" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:02:07.40" />
                    <SPLIT distance="200" swimtime="00:02:55.81" />
                    <SPLIT distance="250" swimtime="00:03:43.04" />
                    <SPLIT distance="300" swimtime="00:04:31.79" />
                    <SPLIT distance="350" swimtime="00:05:19.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" license="502805700158" swrid="5506643" athleteid="9337">
              <RESULTS>
                <RESULT eventid="6077" points="326" swimtime="00:00:33.72" resultid="9338" heatid="11408" lane="9" entrytime="00:00:34.02" entrycourse="SCM" />
                <RESULT eventid="6306" points="259" reactiontime="+105" swimtime="00:01:20.34" resultid="9339" heatid="11469" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="283" reactiontime="+102" swimtime="00:01:36.84" resultid="9340" heatid="11516" lane="7" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="327" reactiontime="+111" swimtime="00:00:42.18" resultid="9341" heatid="11617" lane="6" entrytime="00:00:43.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Piekarski" birthdate="1986-04-22" gender="M" nation="POL" license="502805700144" swrid="5537481" athleteid="9318">
              <RESULTS>
                <RESULT eventid="6077" points="194" reactiontime="+91" swimtime="00:00:38.02" resultid="9319" heatid="11406" lane="0" entrytime="00:00:36.83" />
                <RESULT eventid="6111" points="128" reactiontime="+104" swimtime="00:04:12.57" resultid="9320" heatid="11428" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.55" />
                    <SPLIT distance="100" swimtime="00:02:14.42" />
                    <SPLIT distance="150" swimtime="00:03:16.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" swrid="5464087" athleteid="9279">
              <RESULTS>
                <RESULT eventid="6077" points="494" reactiontime="+98" swimtime="00:00:35.91" resultid="9280" heatid="11408" lane="3" entrytime="00:00:33.40" />
                <RESULT eventid="6111" points="480" reactiontime="+103" swimtime="00:03:46.89" resultid="9281" heatid="11428" lane="0" entrytime="00:03:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:50.94" />
                    <SPLIT distance="150" swimtime="00:02:59.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="517" reactiontime="+105" swimtime="00:01:20.50" resultid="9282" heatid="11470" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="478" reactiontime="+109" swimtime="00:01:39.21" resultid="9283" heatid="11490" lane="7" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="505" reactiontime="+97" swimtime="00:03:05.79" resultid="9284" heatid="11564" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:17.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="540" reactiontime="+107" swimtime="00:06:42.58" resultid="9285" heatid="11632" lane="2" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:32.46" />
                    <SPLIT distance="150" swimtime="00:02:24.04" />
                    <SPLIT distance="200" swimtime="00:03:15.86" />
                    <SPLIT distance="250" swimtime="00:04:07.28" />
                    <SPLIT distance="300" swimtime="00:04:59.17" />
                    <SPLIT distance="350" swimtime="00:05:51.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="9304">
              <RESULTS>
                <RESULT eventid="6077" points="494" reactiontime="+101" swimtime="00:00:33.95" resultid="9305" heatid="11407" lane="5" entrytime="00:00:34.63" entrycourse="SCM" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="9306" heatid="11429" lane="8" entrytime="00:03:12.00" />
                <RESULT eventid="6238" points="377" reactiontime="+72" swimtime="00:00:43.47" resultid="9307" heatid="11444" lane="3" entrytime="00:00:48.10" entrycourse="SCM" />
                <RESULT eventid="6306" points="455" reactiontime="+77" swimtime="00:01:17.84" resultid="9308" heatid="11470" lane="0" entrytime="00:01:22.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="384" swimtime="00:01:41.55" resultid="9309" heatid="11517" lane="9" entrytime="00:01:40.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="286" reactiontime="+68" swimtime="00:01:42.58" resultid="9310" heatid="11550" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="370" swimtime="00:00:45.58" resultid="9311" heatid="11617" lane="9" entrytime="00:00:44.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska." birthdate="1984-02-23" gender="F" nation="POL" license="102805600050" swrid="5537471" athleteid="9364">
              <RESULTS>
                <RESULT eventid="6186" points="447" reactiontime="+43" swimtime="00:23:59.89" resultid="9365" heatid="11650" lane="9" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                    <SPLIT distance="200" swimtime="00:02:58.68" />
                    <SPLIT distance="250" swimtime="00:03:47.44" />
                    <SPLIT distance="300" swimtime="00:04:37.49" />
                    <SPLIT distance="350" swimtime="00:05:25.90" />
                    <SPLIT distance="400" swimtime="00:06:14.62" />
                    <SPLIT distance="450" swimtime="00:07:02.65" />
                    <SPLIT distance="500" swimtime="00:07:50.48" />
                    <SPLIT distance="550" swimtime="00:08:38.39" />
                    <SPLIT distance="600" swimtime="00:09:27.18" />
                    <SPLIT distance="650" swimtime="00:10:14.87" />
                    <SPLIT distance="700" swimtime="00:11:02.97" />
                    <SPLIT distance="750" swimtime="00:11:51.53" />
                    <SPLIT distance="800" swimtime="00:12:39.63" />
                    <SPLIT distance="850" swimtime="00:13:28.17" />
                    <SPLIT distance="900" swimtime="00:14:17.09" />
                    <SPLIT distance="950" swimtime="00:15:05.67" />
                    <SPLIT distance="1000" swimtime="00:15:54.40" />
                    <SPLIT distance="1050" swimtime="00:16:42.98" />
                    <SPLIT distance="1100" swimtime="00:17:31.75" />
                    <SPLIT distance="1150" swimtime="00:18:20.22" />
                    <SPLIT distance="1200" swimtime="00:19:08.97" />
                    <SPLIT distance="1250" swimtime="00:19:57.90" />
                    <SPLIT distance="1300" swimtime="00:20:46.20" />
                    <SPLIT distance="1350" swimtime="00:21:35.11" />
                    <SPLIT distance="1400" swimtime="00:22:23.75" />
                    <SPLIT distance="1450" swimtime="00:23:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="387" reactiontime="+86" swimtime="00:03:32.90" resultid="9366" heatid="11453" lane="5" entrytime="00:03:28.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="100" swimtime="00:01:39.81" />
                    <SPLIT distance="150" swimtime="00:02:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="408" reactiontime="+82" swimtime="00:01:29.18" resultid="9367" heatid="11483" lane="8" entrytime="00:01:39.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="364" reactiontime="+88" swimtime="00:01:36.70" resultid="9368" heatid="11511" lane="7" entrytime="00:01:36.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" status="DNS" swimtime="00:00:00.00" resultid="9369" heatid="11557" lane="1" entrytime="00:02:56.43" />
                <RESULT eventid="6687" points="381" reactiontime="+81" swimtime="00:00:43.66" resultid="9370" heatid="11611" lane="0" entrytime="00:00:45.01" />
                <RESULT eventid="6721" points="401" reactiontime="+87" swimtime="00:06:10.31" resultid="9371" heatid="11626" lane="4" entrytime="00:06:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                    <SPLIT distance="200" swimtime="00:02:59.28" />
                    <SPLIT distance="250" swimtime="00:03:47.41" />
                    <SPLIT distance="300" swimtime="00:04:36.11" />
                    <SPLIT distance="350" swimtime="00:05:24.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="9256">
              <RESULTS>
                <RESULT eventid="6059" points="184" swimtime="00:00:46.20" resultid="9257" heatid="11396" lane="1" entrytime="00:00:49.01" entrycourse="SCM" />
                <RESULT eventid="6094" status="DNS" swimtime="00:00:00.00" resultid="9258" heatid="11421" lane="1" entrytime="00:04:50.00" />
                <RESULT eventid="6255" points="185" reactiontime="+107" swimtime="00:04:51.23" resultid="9259" heatid="11452" lane="8" entrytime="00:05:02.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.43" />
                    <SPLIT distance="100" swimtime="00:02:21.27" />
                    <SPLIT distance="150" swimtime="00:03:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" status="DNS" swimtime="00:00:00.00" resultid="9260" heatid="11482" lane="0" entrytime="00:02:20.00" />
                <RESULT eventid="6415" points="204" reactiontime="+110" swimtime="00:02:08.44" resultid="9261" heatid="11510" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" status="DNS" swimtime="00:00:00.00" resultid="9262" heatid="11556" lane="9" entrytime="00:04:00.00" />
                <RESULT eventid="6687" points="199" reactiontime="+111" swimtime="00:00:58.74" resultid="9263" heatid="11609" lane="7" entrytime="00:01:00.34" entrycourse="SCM" />
                <RESULT eventid="6721" points="135" swimtime="00:08:59.37" resultid="9264" heatid="11625" lane="0" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.53" />
                    <SPLIT distance="100" swimtime="00:02:08.70" />
                    <SPLIT distance="150" swimtime="00:03:17.12" />
                    <SPLIT distance="200" swimtime="00:04:27.64" />
                    <SPLIT distance="250" swimtime="00:05:38.05" />
                    <SPLIT distance="300" swimtime="00:06:49.01" />
                    <SPLIT distance="350" swimtime="00:07:58.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+94" swimtime="00:02:37.82" resultid="9412" heatid="11583" lane="1" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9385" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="9358" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="9321" number="3" reactiontime="+82" />
                    <RELAYPOSITION athleteid="9279" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" reactiontime="+98" swimtime="00:02:48.19" resultid="9416" heatid="12331" lane="7" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:01:39.35" />
                    <SPLIT distance="150" swimtime="00:02:13.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9385" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="9358" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="9321" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="9279" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+106" status="DNF" swimtime="00:00:00.00" resultid="9413" heatid="11583" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9372" number="1" reactiontime="+106" status="DSQ" />
                    <RELAYPOSITION athleteid="9330" number="2" reactiontime="+10" status="DSQ" />
                    <RELAYPOSITION athleteid="9377" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="9390" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+85" swimtime="00:01:58.69" resultid="9414" heatid="11583" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                    <SPLIT distance="100" swimtime="00:01:02.73" />
                    <SPLIT distance="150" swimtime="00:01:33.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9295" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="9312" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="9286" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9351" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" status="DNS" swimtime="00:00:00.00" resultid="9418" heatid="12331" lane="3" entrytime="00:02:03.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9295" number="1" />
                    <RELAYPOSITION athleteid="9351" number="2" />
                    <RELAYPOSITION athleteid="9286" number="3" />
                    <RELAYPOSITION athleteid="9312" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+91" swimtime="00:02:26.44" resultid="9411" heatid="11581" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9248" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="9233" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="9342" number="3" />
                    <RELAYPOSITION athleteid="9272" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" reactiontime="+79" swimtime="00:02:40.06" resultid="9415" heatid="11639" lane="3" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9248" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="9233" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="9272" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="9342" number="4" reactiontime="+82" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+71" swimtime="00:02:11.43" resultid="9408" heatid="11436" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:39.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9330" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="9248" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9272" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="9321" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+83" swimtime="00:02:29.03" resultid="9410" heatid="11506" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:22.40" />
                    <SPLIT distance="150" swimtime="00:01:55.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9248" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="9358" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="9272" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="9330" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+97" swimtime="00:02:27.84" resultid="9409" heatid="11435" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:55.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9377" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="9265" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="9342" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="9372" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8125" name="SMT Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Bartek" lastname="Lasek" birthdate="1977-02-21" gender="M" nation="POL" athleteid="8223">
              <RESULTS>
                <RESULT eventid="6306" points="232" reactiontime="+98" swimtime="00:01:26.07" resultid="8224" heatid="11468" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="215" swimtime="00:01:39.99" resultid="8225" heatid="11488" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="172" reactiontime="+100" swimtime="00:00:46.13" resultid="8226" heatid="11533" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Sawrymowicz" birthdate="1957-07-26" gender="M" nation="POL" athleteid="8143">
              <RESULTS>
                <RESULT eventid="6340" points="272" swimtime="00:01:49.11" resultid="8144" heatid="11489" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="150" swimtime="00:00:57.41" resultid="8145" heatid="11533" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Kramek" birthdate="1992-02-04" gender="M" nation="POL" swrid="4072220" athleteid="8172">
              <RESULTS>
                <RESULT eventid="6077" points="727" swimtime="00:00:24.61" resultid="8173" heatid="11416" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="6111" points="459" reactiontime="+86" swimtime="00:02:33.04" resultid="8174" heatid="11433" lane="8" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="730" reactiontime="+73" swimtime="00:00:54.45" resultid="8175" heatid="11477" lane="6" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="502" reactiontime="+77" swimtime="00:01:09.18" resultid="8176" heatid="11496" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="597" reactiontime="+74" swimtime="00:00:27.16" resultid="8177" heatid="11537" lane="2" entrytime="00:00:30.48" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Zielińska" birthdate="1980-12-12" gender="F" nation="POL" swrid="5185937" athleteid="8160">
              <RESULTS>
                <RESULT eventid="6094" points="580" swimtime="00:02:56.01" resultid="8161" heatid="11423" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:14.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="552" reactiontime="+81" swimtime="00:00:37.22" resultid="8162" heatid="11440" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="6323" points="599" reactiontime="+76" swimtime="00:01:20.80" resultid="8163" heatid="11484" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="632" reactiontime="+71" swimtime="00:01:19.16" resultid="8164" heatid="11545" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="519" swimtime="00:02:40.88" resultid="8165" heatid="11558" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:01:58.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="647" reactiontime="+74" swimtime="00:02:52.66" resultid="8166" heatid="11600" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:23.73" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" status="DNS" swimtime="00:00:00.00" resultid="8167" heatid="11627" lane="4" entrytime="00:05:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Ryczak" birthdate="1996-04-22" gender="F" nation="POL" swrid="4225999" athleteid="8191">
              <RESULTS>
                <RESULT eventid="6059" points="700" reactiontime="+74" swimtime="00:00:28.48" resultid="8192" heatid="11401" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="6220" points="883" reactiontime="+68" swimtime="00:00:30.79" resultid="8193" heatid="11441" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="6289" status="DNS" swimtime="00:00:00.00" resultid="8194" heatid="11466" lane="7" entrytime="00:01:04.00" />
                <RESULT eventid="6484" points="811" reactiontime="+64" swimtime="00:01:08.36" resultid="8195" heatid="11546" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Wojnowski" birthdate="1966-07-12" gender="M" nation="POL" athleteid="8201">
              <RESULTS>
                <RESULT eventid="6077" points="665" swimtime="00:00:29.82" resultid="8202" heatid="11412" lane="4" entrytime="00:00:28.30" />
                <RESULT eventid="6467" points="709" reactiontime="+82" swimtime="00:00:31.45" resultid="8203" heatid="11538" lane="1" entrytime="00:00:29.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Rożek" birthdate="1984-05-09" gender="M" nation="POL" athleteid="8216">
              <RESULTS>
                <RESULT eventid="6169" reactiontime="+93" status="OTL" swimtime="00:00:00.00" resultid="8217" heatid="11647" lane="2" entrytime="00:12:45.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:14.53" />
                    <SPLIT distance="200" swimtime="00:03:02.59" />
                    <SPLIT distance="250" swimtime="00:03:51.36" />
                    <SPLIT distance="300" swimtime="00:04:40.61" />
                    <SPLIT distance="350" swimtime="00:05:29.13" />
                    <SPLIT distance="400" swimtime="00:06:18.04" />
                    <SPLIT distance="450" swimtime="00:07:07.69" />
                    <SPLIT distance="500" swimtime="00:07:57.25" />
                    <SPLIT distance="550" swimtime="00:08:46.22" />
                    <SPLIT distance="600" swimtime="00:09:35.28" />
                    <SPLIT distance="650" swimtime="00:10:24.66" />
                    <SPLIT distance="700" swimtime="00:11:13.87" />
                    <SPLIT distance="750" swimtime="00:12:02.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="321" reactiontime="+87" swimtime="00:01:12.05" resultid="8218" heatid="11472" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="266" reactiontime="+75" swimtime="00:01:28.30" resultid="8219" heatid="11490" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="241" swimtime="00:00:37.95" resultid="8220" heatid="11534" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="6535" points="297" reactiontime="+83" swimtime="00:02:46.96" resultid="8221" heatid="11565" lane="6" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="298" reactiontime="+82" swimtime="00:06:02.65" resultid="8222" heatid="11632" lane="4" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                    <SPLIT distance="200" swimtime="00:02:55.51" />
                    <SPLIT distance="250" swimtime="00:03:42.93" />
                    <SPLIT distance="300" swimtime="00:04:30.76" />
                    <SPLIT distance="350" swimtime="00:05:18.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Stępień-Gielo" birthdate="1961-05-03" gender="F" nation="POL" athleteid="8151">
              <RESULTS>
                <RESULT eventid="6059" points="551" reactiontime="+89" swimtime="00:00:37.82" resultid="8152" heatid="11397" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="6145" points="474" swimtime="00:14:47.64" resultid="8153" heatid="11644" lane="1" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:43.25" />
                    <SPLIT distance="150" swimtime="00:02:37.37" />
                    <SPLIT distance="200" swimtime="00:04:28.74" />
                    <SPLIT distance="250" swimtime="00:06:22.88" />
                    <SPLIT distance="300" swimtime="00:08:15.57" />
                    <SPLIT distance="450" swimtime="00:10:09.82" />
                    <SPLIT distance="500" swimtime="00:12:02.94" />
                    <SPLIT distance="750" swimtime="00:13:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="622" reactiontime="+90" swimtime="00:03:39.53" resultid="8154" heatid="11453" lane="0" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:44.18" />
                    <SPLIT distance="150" swimtime="00:02:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="530" swimtime="00:01:37.71" resultid="8155" heatid="11482" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="603" reactiontime="+89" swimtime="00:01:40.77" resultid="8156" heatid="11511" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="441" reactiontime="+82" swimtime="00:01:46.51" resultid="8157" heatid="11545" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="649" reactiontime="+90" swimtime="00:00:44.01" resultid="8158" heatid="11610" lane="5" entrytime="00:00:46.50" />
                <RESULT eventid="6721" points="391" reactiontime="+96" swimtime="00:07:11.16" resultid="8159" heatid="11625" lane="2" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                    <SPLIT distance="100" swimtime="00:01:44.38" />
                    <SPLIT distance="150" swimtime="00:02:39.80" />
                    <SPLIT distance="200" swimtime="00:03:34.82" />
                    <SPLIT distance="250" swimtime="00:04:30.04" />
                    <SPLIT distance="300" swimtime="00:05:25.42" />
                    <SPLIT distance="350" swimtime="00:06:20.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Usewicz" birthdate="1994-08-12" gender="F" nation="POL" athleteid="8178">
              <RESULTS>
                <RESULT eventid="6059" points="405" reactiontime="+85" swimtime="00:00:34.17" resultid="8179" heatid="11398" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="6289" points="374" swimtime="00:01:17.83" resultid="8180" heatid="11463" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="354" reactiontime="+87" swimtime="00:02:56.72" resultid="8181" heatid="11558" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="294" reactiontime="+101" swimtime="00:06:42.58" resultid="8182" heatid="11625" lane="3" entrytime="00:06:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:34.84" />
                    <SPLIT distance="150" swimtime="00:02:26.35" />
                    <SPLIT distance="200" swimtime="00:03:19.46" />
                    <SPLIT distance="250" swimtime="00:04:13.00" />
                    <SPLIT distance="300" swimtime="00:05:05.11" />
                    <SPLIT distance="350" swimtime="00:05:56.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tyberiusz" lastname="Frymus" birthdate="1995-01-13" gender="M" nation="POL" swrid="4157782" athleteid="8168">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="8169" heatid="11417" lane="7" entrytime="00:00:25.03" />
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="8170" heatid="11521" lane="1" entrytime="00:01:08.00" />
                <RESULT eventid="6704" points="779" swimtime="00:00:30.71" resultid="8171" heatid="11623" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Adamiak" birthdate="1987-08-03" gender="F" nation="POL" athleteid="8126">
              <RESULTS>
                <RESULT eventid="6094" points="265" reactiontime="+87" swimtime="00:03:46.10" resultid="8127" heatid="11422" lane="9" entrytime="00:03:30.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                    <SPLIT distance="150" swimtime="00:02:54.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" reactiontime="+102" status="OTL" swimtime="00:00:00.00" resultid="8128" heatid="11644" lane="2" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:38.37" />
                    <SPLIT distance="150" swimtime="00:02:32.43" />
                    <SPLIT distance="200" swimtime="00:03:26.91" />
                    <SPLIT distance="250" swimtime="00:04:21.84" />
                    <SPLIT distance="300" swimtime="00:05:17.78" />
                    <SPLIT distance="350" swimtime="00:06:13.97" />
                    <SPLIT distance="400" swimtime="00:07:10.06" />
                    <SPLIT distance="450" swimtime="00:08:05.53" />
                    <SPLIT distance="500" swimtime="00:09:01.69" />
                    <SPLIT distance="550" swimtime="00:09:56.92" />
                    <SPLIT distance="600" swimtime="00:10:52.21" />
                    <SPLIT distance="650" swimtime="00:11:47.69" />
                    <SPLIT distance="700" swimtime="00:12:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="312" reactiontime="+95" swimtime="00:07:44.89" resultid="8129" heatid="11573" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                    <SPLIT distance="100" swimtime="00:01:49.91" />
                    <SPLIT distance="150" swimtime="00:02:54.87" />
                    <SPLIT distance="200" swimtime="00:05:00.81" />
                    <SPLIT distance="250" swimtime="00:06:01.49" />
                    <SPLIT distance="300" swimtime="00:06:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="257" reactiontime="+100" swimtime="00:07:09.34" resultid="8130" heatid="11625" lane="5" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:38.37" />
                    <SPLIT distance="150" swimtime="00:02:33.83" />
                    <SPLIT distance="200" swimtime="00:03:28.63" />
                    <SPLIT distance="250" swimtime="00:04:24.24" />
                    <SPLIT distance="300" swimtime="00:05:20.45" />
                    <SPLIT distance="350" swimtime="00:06:16.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Kowalczyk" birthdate="1976-01-31" gender="F" nation="POL" athleteid="8209">
              <RESULTS>
                <RESULT eventid="6059" points="550" reactiontime="+90" swimtime="00:00:32.84" resultid="8210" heatid="11398" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="6094" points="562" reactiontime="+97" swimtime="00:03:01.87" resultid="8211" heatid="11423" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="150" swimtime="00:02:18.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="574" reactiontime="+98" swimtime="00:01:23.18" resultid="8212" heatid="11485" lane="9" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="579" swimtime="00:00:36.00" resultid="8213" heatid="11526" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="6518" points="481" reactiontime="+93" swimtime="00:02:46.51" resultid="8214" heatid="11558" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" status="DNS" swimtime="00:00:00.00" resultid="8215" heatid="11627" lane="7" entrytime="00:05:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Zieliński" birthdate="1992-09-02" gender="M" nation="POL" swrid="4072211" athleteid="8189">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="8190" heatid="11419" lane="9" entrytime="00:00:23.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Zając" birthdate="1966-06-30" gender="M" nation="POL" athleteid="8196">
              <RESULTS>
                <RESULT eventid="6077" points="629" reactiontime="+93" swimtime="00:00:30.38" resultid="8197" heatid="11410" lane="3" entrytime="00:00:31.00" />
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G2" eventid="6340" reactiontime="+95" status="DSQ" swimtime="00:00:00.00" resultid="8198" heatid="11491" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="584" reactiontime="+88" swimtime="00:00:33.55" resultid="8199" heatid="11535" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="6704" points="397" reactiontime="+92" swimtime="00:00:41.48" resultid="8200" heatid="11619" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Król" birthdate="1977-05-26" gender="M" nation="POL" athleteid="8131">
              <RESULTS>
                <RESULT eventid="6077" points="293" reactiontime="+81" swimtime="00:00:35.92" resultid="8132" heatid="11408" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="6169" reactiontime="+101" status="OTL" swimtime="00:00:00.00" resultid="8133" heatid="11647" lane="8" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:36.51" />
                    <SPLIT distance="150" swimtime="00:02:28.92" />
                    <SPLIT distance="200" swimtime="00:03:21.42" />
                    <SPLIT distance="250" swimtime="00:04:14.65" />
                    <SPLIT distance="300" swimtime="00:05:08.13" />
                    <SPLIT distance="350" swimtime="00:06:03.05" />
                    <SPLIT distance="400" swimtime="00:06:57.35" />
                    <SPLIT distance="450" swimtime="00:07:51.93" />
                    <SPLIT distance="500" swimtime="00:08:46.53" />
                    <SPLIT distance="550" swimtime="00:09:41.60" />
                    <SPLIT distance="600" swimtime="00:10:35.93" />
                    <SPLIT distance="650" swimtime="00:11:29.18" />
                    <SPLIT distance="700" swimtime="00:12:23.24" />
                    <SPLIT distance="750" swimtime="00:13:16.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Kudra" birthdate="1959-11-24" gender="F" nation="POL" athleteid="8146">
              <RESULTS>
                <RESULT eventid="6059" points="247" reactiontime="+158" swimtime="00:00:49.42" resultid="8147" heatid="11396" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="6289" points="168" reactiontime="+135" swimtime="00:02:03.31" resultid="8148" heatid="11462" lane="3" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="364" swimtime="00:01:59.24" resultid="8149" heatid="11510" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="347" swimtime="00:00:54.24" resultid="8150" heatid="11609" lane="4" entrytime="00:00:55.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Moskalenko" birthdate="2000-12-01" gender="F" nation="POL" athleteid="8183">
              <RESULTS>
                <RESULT eventid="6059" points="435" reactiontime="+68" swimtime="00:00:34.34" resultid="8184" heatid="11398" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="6145" points="315" reactiontime="+85" swimtime="00:13:19.24" resultid="8185" heatid="11644" lane="5" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:24.57" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                    <SPLIT distance="200" swimtime="00:03:01.54" />
                    <SPLIT distance="250" swimtime="00:03:51.22" />
                    <SPLIT distance="300" swimtime="00:04:42.01" />
                    <SPLIT distance="350" swimtime="00:06:26.38" />
                    <SPLIT distance="400" swimtime="00:07:20.14" />
                    <SPLIT distance="450" swimtime="00:08:13.43" />
                    <SPLIT distance="500" swimtime="00:09:05.50" />
                    <SPLIT distance="550" swimtime="00:09:56.92" />
                    <SPLIT distance="600" swimtime="00:10:49.57" />
                    <SPLIT distance="650" swimtime="00:11:41.37" />
                    <SPLIT distance="700" swimtime="00:12:31.94" />
                    <SPLIT distance="750" swimtime="00:13:19.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="409" reactiontime="+76" swimtime="00:01:17.85" resultid="8186" heatid="11464" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="388" reactiontime="+75" swimtime="00:02:48.82" resultid="8187" heatid="11557" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="326" swimtime="00:06:12.90" resultid="8188" heatid="11627" lane="0" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:02:14.07" />
                    <SPLIT distance="150" swimtime="00:03:02.37" />
                    <SPLIT distance="200" swimtime="00:03:51.29" />
                    <SPLIT distance="250" swimtime="00:04:39.85" />
                    <SPLIT distance="300" swimtime="00:05:28.24" />
                    <SPLIT distance="350" swimtime="00:06:12.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iwona" lastname="Wacławik" birthdate="1965-04-21" gender="F" nation="POL" athleteid="8134">
              <RESULTS>
                <RESULT eventid="6094" points="438" reactiontime="+68" swimtime="00:03:26.61" resultid="8135" heatid="11421" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:38.26" />
                    <SPLIT distance="150" swimtime="00:02:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="422" swimtime="00:13:28.02" resultid="8136" heatid="11644" lane="6" entrytime="00:14:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="100" swimtime="00:01:32.36" />
                    <SPLIT distance="150" swimtime="00:02:22.96" />
                    <SPLIT distance="200" swimtime="00:03:13.97" />
                    <SPLIT distance="250" swimtime="00:04:05.21" />
                    <SPLIT distance="300" swimtime="00:04:57.76" />
                    <SPLIT distance="350" swimtime="00:05:48.83" />
                    <SPLIT distance="400" swimtime="00:06:40.30" />
                    <SPLIT distance="450" swimtime="00:07:31.83" />
                    <SPLIT distance="500" swimtime="00:08:23.48" />
                    <SPLIT distance="550" swimtime="00:09:15.21" />
                    <SPLIT distance="600" swimtime="00:10:06.71" />
                    <SPLIT distance="650" swimtime="00:10:58.41" />
                    <SPLIT distance="700" swimtime="00:11:49.22" />
                    <SPLIT distance="750" swimtime="00:12:39.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="600" reactiontime="+87" swimtime="00:03:39.65" resultid="8137" heatid="11453" lane="7" entrytime="00:03:45.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:46.97" />
                    <SPLIT distance="150" swimtime="00:02:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="494" reactiontime="+88" swimtime="00:01:32.25" resultid="8138" heatid="11483" lane="2" entrytime="00:01:36.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="563" reactiontime="+75" swimtime="00:01:40.73" resultid="8139" heatid="11510" lane="4" entrytime="00:01:46.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="498" reactiontime="+75" swimtime="00:00:40.29" resultid="8140" heatid="11525" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="6618" points="353" reactiontime="+84" swimtime="00:01:41.94" resultid="8141" heatid="11586" lane="3" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="523" reactiontime="+78" swimtime="00:00:46.61" resultid="8142" heatid="11610" lane="3" entrytime="00:00:46.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Krzyżostaniak" birthdate="1993-01-20" gender="F" nation="POL" swrid="4087097" athleteid="8227">
              <RESULTS>
                <RESULT eventid="6220" points="806" reactiontime="+86" swimtime="00:00:31.73" resultid="8228" heatid="11441" lane="7" entrytime="00:00:32.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Zienkiewicz" birthdate="1974-08-12" gender="M" nation="POL" swrid="5185933" athleteid="8204">
              <RESULTS>
                <RESULT eventid="6077" points="476" reactiontime="+73" swimtime="00:00:30.56" resultid="8205" heatid="11410" lane="8" entrytime="00:00:31.20" />
                <RESULT eventid="6306" points="358" reactiontime="+68" swimtime="00:01:14.48" resultid="8206" heatid="11469" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="418" reactiontime="+74" swimtime="00:00:34.32" resultid="8207" heatid="11535" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="6704" points="479" swimtime="00:00:38.69" resultid="8208" heatid="11619" lane="8" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+75" swimtime="00:02:11.84" resultid="8241" heatid="12332" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                    <SPLIT distance="150" swimtime="00:01:40.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8189" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="8204" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="8196" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="8216" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+70" swimtime="00:02:06.16" resultid="8242" heatid="11582" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:37.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8204" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="8223" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="8196" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="8201" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+80" swimtime="00:02:01.91" resultid="8240" heatid="11582" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.64" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:38.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8172" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="8143" number="2" />
                    <RELAYPOSITION athleteid="8216" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="8189" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6755" reactiontime="+69" swimtime="00:02:24.71" resultid="8229" heatid="11639" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8191" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="8209" number="2" />
                    <RELAYPOSITION athleteid="8160" number="3" />
                    <RELAYPOSITION athleteid="8178" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6586" reactiontime="+73" swimtime="00:02:09.15" resultid="8230" heatid="11580" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:39.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8160" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="8178" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="8209" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="8191" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+68" swimtime="00:02:49.29" resultid="8238" heatid="11580" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:11.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8134" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="8146" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8126" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="8151" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" reactiontime="+86" swimtime="00:03:05.49" resultid="8239" heatid="11639" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:41.60" />
                    <SPLIT distance="150" swimtime="00:02:22.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8151" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="8146" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="8134" number="3" />
                    <RELAYPOSITION athleteid="8126" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+95" swimtime="00:02:26.08" resultid="8233" heatid="11434" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:54.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8151" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="8131" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="8134" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="8216" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+83" swimtime="00:02:54.75" resultid="9851" heatid="11506" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:41.39" />
                    <SPLIT distance="150" swimtime="00:02:13.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8151" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="8146" number="2" reactiontime="+104" />
                    <RELAYPOSITION athleteid="8201" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="8143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+68" swimtime="00:02:02.62" resultid="8232" heatid="11506" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:02.80" />
                    <SPLIT distance="150" swimtime="00:01:28.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8191" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="8172" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="8189" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="8178" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+95" swimtime="00:02:05.92" resultid="8234" heatid="11435" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:33.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8196" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="8209" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="8201" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="8160" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+90" swimtime="00:02:31.23" resultid="8235" heatid="11505" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8209" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="8204" number="2" />
                    <RELAYPOSITION athleteid="8196" number="3" />
                    <RELAYPOSITION athleteid="8134" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+71" swimtime="00:01:50.11" resultid="8236" heatid="11435" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="150" swimtime="00:01:25.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8191" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8227" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="8172" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="8189" number="4" reactiontime="+83" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+76" status="EXH" swimtime="00:02:42.14" resultid="8237" heatid="11505" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:28.41" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8160" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="8183" number="2" reactiontime="+83" />
                    <RELAYPOSITION athleteid="8216" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="8223" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03706" nation="POL" region="06" clubid="9438" name="Stowarzyszenie SIEMACHA">
          <ATHLETES>
            <ATHLETE firstname="Ada" lastname="Malinowska" birthdate="1999-05-27" gender="F" nation="POL" swrid="4780924" athleteid="7500">
              <RESULTS>
                <RESULT eventid="6059" points="681" swimtime="00:00:29.57" resultid="7501" heatid="11400" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="6094" status="DNS" swimtime="00:00:00.00" resultid="7502" heatid="11420" lane="7" />
                <RESULT eventid="6220" points="503" reactiontime="+65" swimtime="00:00:36.46" resultid="7503" heatid="11440" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="6289" points="619" reactiontime="+77" swimtime="00:01:07.81" resultid="7504" heatid="11465" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="666" reactiontime="+78" swimtime="00:00:31.89" resultid="7505" heatid="11527" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="6484" points="490" reactiontime="+76" swimtime="00:01:19.44" resultid="7506" heatid="11543" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="617" reactiontime="+77" swimtime="00:01:12.97" resultid="7507" heatid="11587" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="606" reactiontime="+77" swimtime="00:00:38.41" resultid="7508" heatid="11611" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Palmowska- Latuszek" birthdate="1985-08-01" gender="F" nation="POL" license="503706600141" swrid="4992815" athleteid="9439">
              <RESULTS>
                <RESULT eventid="6059" points="717" swimtime="00:00:29.25" resultid="9440" heatid="11400" lane="9" entrytime="00:00:30.39" entrycourse="SCM" />
                <RESULT eventid="6094" points="704" reactiontime="+67" swimtime="00:02:43.26" resultid="9441" heatid="11424" lane="0" entrytime="00:02:45.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="785" reactiontime="+60" swimtime="00:00:33.48" resultid="9442" heatid="11441" lane="1" entrytime="00:00:33.62" entrycourse="SCM" />
                <RESULT eventid="6289" points="692" reactiontime="+69" swimtime="00:01:05.32" resultid="9443" heatid="11466" lane="9" entrytime="00:01:06.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="766" reactiontime="+64" swimtime="00:01:12.04" resultid="9444" heatid="11546" lane="2" entrytime="00:01:13.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="671" reactiontime="+77" swimtime="00:02:26.31" resultid="9445" heatid="11559" lane="7" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="729" reactiontime="+59" swimtime="00:02:38.66" resultid="9446" heatid="11600" lane="3" entrytime="00:02:39.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:15.38" />
                    <SPLIT distance="150" swimtime="00:01:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="616" swimtime="00:05:20.88" resultid="9447" heatid="11628" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                    <SPLIT distance="200" swimtime="00:02:33.30" />
                    <SPLIT distance="250" swimtime="00:03:15.23" />
                    <SPLIT distance="300" swimtime="00:03:57.06" />
                    <SPLIT distance="350" swimtime="00:04:39.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Kolba" birthdate="1996-10-30" gender="F" nation="POL" athleteid="7497">
              <RESULTS>
                <RESULT eventid="6220" points="721" reactiontime="+64" swimtime="00:00:32.94" resultid="7498" heatid="11441" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="6484" points="697" reactiontime="+71" swimtime="00:01:11.92" resultid="7499" heatid="11546" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8445" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Grzelak" birthdate="1970-01-01" gender="M" nation="POL" swrid="4951293" athleteid="8444">
              <RESULTS>
                <RESULT eventid="6374" points="273" reactiontime="+77" swimtime="00:03:34.10" resultid="8446" heatid="11502" lane="8" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:32.42" />
                    <SPLIT distance="150" swimtime="00:02:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="326" reactiontime="+81" swimtime="00:07:14.80" resultid="8447" heatid="11577" lane="2" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                    <SPLIT distance="150" swimtime="00:02:36.80" />
                    <SPLIT distance="200" swimtime="00:03:39.49" />
                    <SPLIT distance="250" swimtime="00:04:40.64" />
                    <SPLIT distance="300" swimtime="00:05:42.29" />
                    <SPLIT distance="350" swimtime="00:06:29.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="K S PIETRA" nation="POL" clubid="6875" name="Klub  Sportowy PIETRASZYN">
          <ATHLETES>
            <ATHLETE firstname="Adolf" lastname="Piechula" birthdate="1957-04-11" gender="M" nation="POL" swrid="4992724" athleteid="6876">
              <RESULTS>
                <RESULT eventid="6077" points="560" reactiontime="+83" swimtime="00:00:33.46" resultid="6877" heatid="11403" lane="4" />
                <RESULT eventid="6111" points="550" reactiontime="+92" swimtime="00:03:13.52" resultid="6878" heatid="11425" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:31.95" />
                    <SPLIT distance="150" swimtime="00:02:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="636" reactiontime="+93" swimtime="00:03:31.27" resultid="6879" heatid="11455" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:38.38" />
                    <SPLIT distance="150" swimtime="00:02:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="472" reactiontime="+94" swimtime="00:03:34.86" resultid="6880" heatid="11500" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="531" reactiontime="+96" swimtime="00:01:34.96" resultid="6881" heatid="11517" lane="2" entrytime="00:01:36.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="613" swimtime="00:07:13.37" resultid="6882" heatid="11575" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:40.90" />
                    <SPLIT distance="150" swimtime="00:02:37.69" />
                    <SPLIT distance="200" swimtime="00:03:32.81" />
                    <SPLIT distance="250" swimtime="00:04:33.88" />
                    <SPLIT distance="300" swimtime="00:05:34.01" />
                    <SPLIT distance="350" swimtime="00:06:24.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="414" reactiontime="+93" swimtime="00:01:35.53" resultid="6883" heatid="11591" lane="3" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="517" reactiontime="+80" swimtime="00:00:42.09" resultid="6884" heatid="11616" lane="6" entrytime="00:00:46.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7296" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-16" gender="M" nation="POL" license="500309700377" swrid="4186249" athleteid="7297">
              <RESULTS>
                <RESULT eventid="6077" points="792" reactiontime="+74" swimtime="00:00:28.13" resultid="7298" heatid="11412" lane="2" entrytime="00:00:28.75" />
                <RESULT eventid="6111" points="711" reactiontime="+83" swimtime="00:02:38.97" resultid="7299" heatid="11431" lane="7" entrytime="00:02:39.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:02:01.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="804" reactiontime="+77" swimtime="00:01:02.39" resultid="7300" heatid="11475" lane="8" entrytime="00:01:03.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="766" reactiontime="+78" swimtime="00:01:11.84" resultid="7301" heatid="11493" lane="7" entrytime="00:01:12.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="765" reactiontime="+75" swimtime="00:00:30.67" resultid="7302" heatid="11536" lane="5" entrytime="00:00:31.35" />
                <RESULT eventid="6501" points="633" reactiontime="+86" swimtime="00:01:15.40" resultid="7303" heatid="11551" lane="7" entrytime="00:01:16.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="710" reactiontime="+85" swimtime="00:01:10.68" resultid="7304" heatid="11593" lane="7" entrytime="00:01:12.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="588" reactiontime="+77" swimtime="00:00:36.40" resultid="7305" heatid="11619" lane="6" entrytime="00:00:37.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Wasilewicz" birthdate="1959-01-01" gender="F" nation="POL" license="5000309600230" swrid="4876623" athleteid="7306">
              <RESULTS>
                <RESULT eventid="6059" points="570" swimtime="00:00:37.39" resultid="7307" heatid="11397" lane="6" entrytime="00:00:37.93" />
                <RESULT eventid="6289" points="465" swimtime="00:01:27.91" resultid="7308" heatid="11463" lane="0" entrytime="00:01:28.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="361" swimtime="00:03:25.98" resultid="7309" heatid="11556" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="334" swimtime="00:00:54.90" resultid="7310" heatid="11609" lane="8" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Matusik" birthdate="1956-01-01" gender="M" nation="POL" license="5000309700229" swrid="4876624" athleteid="7311">
              <RESULTS>
                <RESULT eventid="6077" points="453" reactiontime="+85" swimtime="00:00:35.89" resultid="7312" heatid="11407" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="6238" points="274" reactiontime="+104" swimtime="00:00:51.28" resultid="7313" heatid="11445" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="6340" points="451" reactiontime="+77" swimtime="00:01:32.19" resultid="7314" heatid="11491" lane="9" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="565" reactiontime="+95" swimtime="00:01:33.02" resultid="7315" heatid="11517" lane="8" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="494" reactiontime="+85" swimtime="00:00:38.65" resultid="7316" heatid="11533" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="6704" points="571" reactiontime="+87" swimtime="00:00:40.73" resultid="7317" heatid="11618" lane="0" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7484" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Zawadka" birthdate="1978-01-10" gender="M" nation="POL" athleteid="7483">
              <RESULTS>
                <RESULT eventid="6238" points="376" reactiontime="+73" swimtime="00:00:37.59" resultid="7485" heatid="11443" lane="2" />
                <RESULT eventid="6340" points="484" reactiontime="+89" swimtime="00:01:16.16" resultid="7486" heatid="11490" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="431" reactiontime="+77" swimtime="00:00:33.26" resultid="7487" heatid="11535" lane="3" entrytime="00:00:33.44" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GER" clubid="6788" name="SG Erkelenz - Hückelhoven">
          <ATHLETES>
            <ATHLETE firstname="Darius" lastname="Andrzejczak" birthdate="1967-01-01" gender="M" nation="GER" swrid="4906823" athleteid="6787">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6077" points="1012" reactiontime="+80" swimtime="00:00:25.92" resultid="6789" heatid="11416" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="6111" points="730" reactiontime="+87" swimtime="00:02:37.59" resultid="6790" heatid="11432" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                    <SPLIT distance="150" swimtime="00:02:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="990" reactiontime="+82" swimtime="00:00:58.22" resultid="6791" heatid="11477" lane="7" entrytime="00:00:58.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="879" reactiontime="+82" swimtime="00:01:08.61" resultid="6792" heatid="11495" lane="3" entrytime="00:01:07.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6467" points="913" reactiontime="+82" swimtime="00:00:28.91" resultid="6793" heatid="11539" lane="3" entrytime="00:00:28.78" entrycourse="SCM" />
                <RESULT eventid="6535" points="819" reactiontime="+86" swimtime="00:02:15.44" resultid="6794" heatid="11569" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="797" reactiontime="+86" swimtime="00:01:08.03" resultid="6795" heatid="11594" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="701" swimtime="00:00:34.33" resultid="6796" heatid="11622" lane="9" entrytime="00:00:33.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11514" nation="POL" region="14" clubid="9432" name="Stowarzyszenie Pływackie Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Diaby - Lipka" birthdate="1980-08-30" gender="F" nation="POL" license="111514600193" athleteid="9436">
              <RESULTS>
                <RESULT eventid="6220" points="670" reactiontime="+91" swimtime="00:00:34.91" resultid="9437" heatid="11437" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" license="511514700195" athleteid="9433">
              <RESULTS>
                <RESULT eventid="6306" points="327" reactiontime="+90" swimtime="00:01:16.79" resultid="9435" heatid="11467" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="287" reactiontime="+84" swimtime="00:02:53.87" resultid="9822" heatid="11561" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:23.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8636" name="START Poznań">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Wróbel" birthdate="1967-02-06" gender="M" nation="POL" athleteid="8654">
              <RESULTS>
                <RESULT eventid="6111" points="712" reactiontime="+84" swimtime="00:02:38.84" resultid="8655" heatid="11431" lane="0" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="760" reactiontime="+84" swimtime="00:01:12.03" resultid="8656" heatid="11494" lane="1" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="807" swimtime="00:00:30.12" resultid="8657" heatid="11537" lane="4" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="6636" points="692" reactiontime="+84" swimtime="00:01:11.29" resultid="8658" heatid="11593" lane="5" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Monczak" birthdate="1967-11-08" gender="M" nation="POL" swrid="4302571" athleteid="8646">
              <RESULTS>
                <RESULT eventid="6077" points="820" reactiontime="+68" swimtime="00:00:27.81" resultid="8647" heatid="11413" lane="2" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="6111" points="806" reactiontime="+74" swimtime="00:02:32.43" resultid="8648" heatid="11431" lane="4" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="905" reactiontime="+72" swimtime="00:00:59.98" resultid="8649" heatid="11477" lane="0" entrytime="00:00:59.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="834" reactiontime="+73" swimtime="00:01:09.84" resultid="8650" heatid="11494" lane="9" entrytime="00:01:11.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="807" reactiontime="+79" swimtime="00:02:16.09" resultid="8651" heatid="11569" lane="3" entrytime="00:02:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:07.31" />
                    <SPLIT distance="150" swimtime="00:01:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="726" reactiontime="+84" swimtime="00:05:38.16" resultid="8652" heatid="11579" lane="9" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:58.86" />
                    <SPLIT distance="200" swimtime="00:02:42.47" />
                    <SPLIT distance="250" swimtime="00:03:32.16" />
                    <SPLIT distance="300" swimtime="00:04:22.72" />
                    <SPLIT distance="350" swimtime="00:05:00.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="802" reactiontime="+77" swimtime="00:04:50.25" resultid="8653" heatid="11637" lane="9" entrytime="00:04:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                    <SPLIT distance="200" swimtime="00:02:22.31" />
                    <SPLIT distance="250" swimtime="00:02:59.77" />
                    <SPLIT distance="300" swimtime="00:03:37.45" />
                    <SPLIT distance="350" swimtime="00:04:14.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Maduzia" birthdate="1984-08-03" gender="F" nation="POL" swrid="4992773" athleteid="8659">
              <RESULTS>
                <RESULT eventid="6059" status="DNS" swimtime="00:00:00.00" resultid="8660" heatid="11398" lane="7" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="6145" reactiontime="+94" status="OTL" swimtime="00:00:00.00" resultid="8661" heatid="11643" lane="0" entrytime="00:12:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="150" swimtime="00:02:14.91" />
                    <SPLIT distance="200" swimtime="00:03:02.34" />
                    <SPLIT distance="250" swimtime="00:03:50.62" />
                    <SPLIT distance="300" swimtime="00:04:38.67" />
                    <SPLIT distance="350" swimtime="00:05:27.32" />
                    <SPLIT distance="400" swimtime="00:06:15.48" />
                    <SPLIT distance="450" swimtime="00:07:04.08" />
                    <SPLIT distance="500" swimtime="00:07:52.19" />
                    <SPLIT distance="550" swimtime="00:08:40.45" />
                    <SPLIT distance="600" swimtime="00:09:28.53" />
                    <SPLIT distance="650" swimtime="00:10:15.51" />
                    <SPLIT distance="700" swimtime="00:11:02.52" />
                    <SPLIT distance="750" swimtime="00:11:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="447" swimtime="00:01:15.54" resultid="8662" heatid="11464" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="408" reactiontime="+88" swimtime="00:03:12.08" resultid="8663" heatid="11499" lane="7" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:22.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="469" reactiontime="+92" swimtime="00:00:36.58" resultid="8664" heatid="11526" lane="0" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="6518" points="445" reactiontime="+91" swimtime="00:02:47.72" resultid="8665" heatid="11557" lane="9" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="424" reactiontime="+93" swimtime="00:01:24.86" resultid="8666" heatid="11587" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="431" reactiontime="+98" swimtime="00:06:01.47" resultid="8667" heatid="11626" lane="5" entrytime="00:06:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:27.06" />
                    <SPLIT distance="150" swimtime="00:02:12.30" />
                    <SPLIT distance="200" swimtime="00:02:58.28" />
                    <SPLIT distance="250" swimtime="00:03:44.21" />
                    <SPLIT distance="300" swimtime="00:04:29.81" />
                    <SPLIT distance="350" swimtime="00:05:16.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kaczmarek" birthdate="1982-10-03" gender="M" nation="POL" swrid="5471723" athleteid="8637">
              <RESULTS>
                <RESULT eventid="6077" points="559" reactiontime="+101" swimtime="00:00:28.16" resultid="8638" heatid="11412" lane="8" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="6111" points="452" reactiontime="+109" swimtime="00:02:46.54" resultid="8639" heatid="11430" lane="8" entrytime="00:02:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="541" reactiontime="+97" swimtime="00:01:02.91" resultid="8640" heatid="11474" lane="9" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" status="DNS" swimtime="00:00:00.00" resultid="8641" heatid="11502" lane="7" entrytime="00:03:20.00" entrycourse="SCM" />
                <RESULT eventid="6467" points="419" reactiontime="+103" swimtime="00:00:33.56" resultid="8642" heatid="11534" lane="5" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="6569" points="378" reactiontime="+110" swimtime="00:06:14.88" resultid="8643" heatid="11577" lane="3" entrytime="00:06:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:19.65" />
                    <SPLIT distance="200" swimtime="00:03:07.11" />
                    <SPLIT distance="250" swimtime="00:03:58.84" />
                    <SPLIT distance="300" swimtime="00:04:50.77" />
                    <SPLIT distance="350" swimtime="00:05:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8644" heatid="11604" lane="0" entrytime="00:03:00.00" entrycourse="SCM" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8645" heatid="11633" lane="6" entrytime="00:05:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kupiszek" birthdate="1984-05-06" gender="M" nation="POL" athleteid="8668">
              <RESULTS>
                <RESULT eventid="6077" points="433" reactiontime="+74" swimtime="00:00:29.10" resultid="8669" heatid="11411" lane="0" entrytime="00:00:30.03" entrycourse="SCM" />
                <RESULT eventid="6238" points="345" reactiontime="+75" swimtime="00:00:34.89" resultid="8670" heatid="11448" lane="9" entrytime="00:00:34.30" entrycourse="SCM" />
                <RESULT eventid="6306" points="428" reactiontime="+74" swimtime="00:01:05.47" resultid="8671" heatid="11473" lane="3" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="351" reactiontime="+78" swimtime="00:01:20.47" resultid="8672" heatid="11492" lane="2" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="8673" heatid="11551" lane="6" entrytime="00:01:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Kapałczyński" birthdate="1964-11-03" gender="M" nation="POL" athleteid="8674">
              <RESULTS>
                <RESULT eventid="6111" points="537" reactiontime="+81" swimtime="00:02:54.57" resultid="8675" heatid="11429" lane="5" entrytime="00:02:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:21.44" />
                    <SPLIT distance="150" swimtime="00:02:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="632" swimtime="00:03:08.71" resultid="8676" heatid="11458" lane="1" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:27.30" />
                    <SPLIT distance="150" swimtime="00:02:17.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="398" reactiontime="+84" swimtime="00:03:08.92" resultid="8677" heatid="11502" lane="5" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                    <SPLIT distance="150" swimtime="00:02:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="452" reactiontime="+94" swimtime="00:06:35.98" resultid="8678" heatid="11578" lane="9" entrytime="00:06:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:27.46" />
                    <SPLIT distance="150" swimtime="00:02:17.05" />
                    <SPLIT distance="200" swimtime="00:03:10.92" />
                    <SPLIT distance="250" swimtime="00:04:06.11" />
                    <SPLIT distance="300" swimtime="00:05:02.32" />
                    <SPLIT distance="350" swimtime="00:05:50.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="487" reactiontime="+88" swimtime="00:01:20.14" resultid="8679" heatid="11592" lane="7" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKKON" nation="POL" clubid="9731" name="IKS Konstancin">
          <ATHLETES>
            <ATHLETE firstname="Rafal" lastname="Juchno" birthdate="1976-10-30" gender="M" nation="POL" license="103714700079" swrid="4992759" athleteid="9732">
              <RESULTS>
                <RESULT eventid="6077" points="534" reactiontime="+85" swimtime="00:00:29.42" resultid="9733" heatid="11411" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="6169" points="375" reactiontime="+99" swimtime="00:12:00.43" resultid="9734" heatid="11647" lane="4" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:22.23" />
                    <SPLIT distance="150" swimtime="00:02:07.59" />
                    <SPLIT distance="200" swimtime="00:02:53.66" />
                    <SPLIT distance="250" swimtime="00:03:39.65" />
                    <SPLIT distance="300" swimtime="00:04:25.77" />
                    <SPLIT distance="350" swimtime="00:05:11.80" />
                    <SPLIT distance="400" swimtime="00:05:57.82" />
                    <SPLIT distance="450" swimtime="00:06:43.89" />
                    <SPLIT distance="500" swimtime="00:07:30.27" />
                    <SPLIT distance="550" swimtime="00:08:17.42" />
                    <SPLIT distance="600" swimtime="00:09:04.31" />
                    <SPLIT distance="650" swimtime="00:09:50.20" />
                    <SPLIT distance="700" swimtime="00:10:35.93" />
                    <SPLIT distance="750" swimtime="00:11:22.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02211" nation="POL" clubid="6800" name="Muks Gilus Gilowice">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" swrid="4292540" athleteid="6900">
              <RESULTS>
                <RESULT eventid="6111" points="757" reactiontime="+75" swimtime="00:02:24.74" resultid="6901" heatid="11432" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6272" points="1091" reactiontime="+74" swimtime="00:02:30.31" resultid="6902" heatid="11460" lane="7" entrytime="00:02:35.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6433" points="981" reactiontime="+71" swimtime="00:01:07.58" resultid="6903" heatid="11520" lane="5" entrytime="00:01:10.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6704" points="1010" reactiontime="+69" swimtime="00:00:30.65" resultid="6904" heatid="11622" lane="3" entrytime="00:00:31.90" />
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="9839" heatid="11579" lane="7" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" clubid="7879" name="Mks Swim Academy Termy Jakuba Oława">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Chorąży" birthdate="1978-09-27" gender="F" nation="POL" license="104501600044" swrid="5506627" athleteid="7880">
              <RESULTS>
                <RESULT eventid="6255" points="677" reactiontime="+93" swimtime="00:03:09.16" resultid="7881" heatid="11454" lane="8" entrytime="00:03:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                    <SPLIT distance="150" swimtime="00:02:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="706" reactiontime="+86" swimtime="00:01:16.49" resultid="7882" heatid="11485" lane="8" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="726" reactiontime="+75" swimtime="00:01:24.21" resultid="7883" heatid="11512" lane="9" entrytime="00:01:25.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="681" reactiontime="+87" swimtime="00:00:33.29" resultid="7884" heatid="11527" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="6687" points="758" reactiontime="+84" swimtime="00:00:37.66" resultid="7885" heatid="11612" lane="0" entrytime="00:00:38.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6844" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-01-01" gender="M" nation="POL" swrid="5416779" athleteid="6843">
              <RESULTS>
                <RESULT eventid="6111" points="236" reactiontime="+97" swimtime="00:03:49.31" resultid="6845" heatid="11427" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.57" />
                    <SPLIT distance="100" swimtime="00:01:57.70" />
                    <SPLIT distance="150" swimtime="00:02:58.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" reactiontime="+109" status="OTL" swimtime="00:00:00.00" resultid="6846" heatid="11647" lane="0" entrytime="00:14:29.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:38.68" />
                    <SPLIT distance="250" swimtime="00:04:32.45" />
                    <SPLIT distance="300" swimtime="00:05:29.95" />
                    <SPLIT distance="400" swimtime="00:07:23.62" />
                    <SPLIT distance="550" swimtime="00:10:14.66" />
                    <SPLIT distance="600" swimtime="00:11:11.45" />
                    <SPLIT distance="650" swimtime="00:12:08.86" />
                    <SPLIT distance="750" swimtime="00:14:01.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="286" reactiontime="+93" swimtime="00:01:28.01" resultid="6847" heatid="11469" lane="0" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" status="DNS" swimtime="00:00:00.00" resultid="6848" heatid="11501" lane="1" entrytime="00:04:20.00" />
                <RESULT eventid="6535" points="250" reactiontime="+93" swimtime="00:03:21.11" resultid="6849" heatid="11563" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                    <SPLIT distance="100" swimtime="00:01:37.22" />
                    <SPLIT distance="150" swimtime="00:02:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="6850" heatid="11576" lane="5" entrytime="00:08:15.00" />
                <RESULT eventid="6636" points="154" reactiontime="+96" swimtime="00:01:57.50" resultid="6851" heatid="11590" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="245" reactiontime="+102" swimtime="00:07:10.84" resultid="6852" heatid="11631" lane="1" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7181" name="Uśks Ostroleka">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Ambroziak" birthdate="1964-05-21" gender="M" nation="POL" athleteid="7182">
              <RESULTS>
                <RESULT eventid="6169" points="333" reactiontime="+88" swimtime="00:13:25.04" resultid="7184" heatid="11648" lane="3" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                    <SPLIT distance="150" swimtime="00:02:22.93" />
                    <SPLIT distance="200" swimtime="00:03:13.54" />
                    <SPLIT distance="250" swimtime="00:04:05.06" />
                    <SPLIT distance="300" swimtime="00:04:55.79" />
                    <SPLIT distance="350" swimtime="00:05:46.57" />
                    <SPLIT distance="400" swimtime="00:06:37.12" />
                    <SPLIT distance="450" swimtime="00:07:28.28" />
                    <SPLIT distance="500" swimtime="00:08:19.62" />
                    <SPLIT distance="550" swimtime="00:09:11.65" />
                    <SPLIT distance="600" swimtime="00:10:03.30" />
                    <SPLIT distance="650" swimtime="00:10:55.95" />
                    <SPLIT distance="700" swimtime="00:11:47.21" />
                    <SPLIT distance="750" swimtime="00:12:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7185" heatid="11563" lane="3" entrytime="00:03:16.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="7186" heatid="11631" lane="2" entrytime="00:07:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Janczewski" birthdate="1990-12-06" gender="M" nation="POL" swrid="5552298" athleteid="7290">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7291" heatid="11417" lane="2" entrytime="00:00:25.00" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7292" heatid="11433" lane="3" entrytime="00:02:18.00" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7293" heatid="11478" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7294" heatid="11541" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7295" heatid="11570" lane="4" entrytime="00:02:04.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8440" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Ptak" birthdate="1983-01-01" gender="M" nation="POL" swrid="4060463" athleteid="8439">
              <RESULTS>
                <RESULT eventid="6272" points="793" reactiontime="+77" swimtime="00:02:31.87" resultid="8441" heatid="11460" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="805" reactiontime="+72" swimtime="00:01:08.25" resultid="8442" heatid="11520" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="794" reactiontime="+77" swimtime="00:00:31.16" resultid="8443" heatid="11622" lane="2" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="8984" name="KS Neptun Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Żukowski" birthdate="1993-04-26" gender="M" nation="POL" license="104901700097" swrid="4087259" athleteid="8985">
              <RESULTS>
                <RESULT eventid="6077" points="884" reactiontime="+75" swimtime="00:00:23.79" resultid="8986" heatid="11419" lane="8" entrytime="00:00:23.50" />
                <RESULT eventid="6340" points="822" reactiontime="+76" swimtime="00:00:58.92" resultid="8987" heatid="11497" lane="6" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="931" reactiontime="+76" swimtime="00:01:03.52" resultid="8988" heatid="11521" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="935" reactiontime="+75" swimtime="00:00:28.90" resultid="8989" heatid="11623" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02902" nation="POL" region="02" clubid="9520" name="Uks Czwórka Nakło">
          <ATHLETES>
            <ATHLETE firstname="Radosław" lastname="Staszkiewicz" birthdate="1968-04-21" gender="M" nation="POL" license="102902700326" swrid="5337392" athleteid="9521">
              <RESULTS>
                <RESULT eventid="6111" points="477" reactiontime="+142" swimtime="00:02:48.86" resultid="9522" heatid="11430" lane="7" entrytime="00:02:47.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="503" swimtime="00:21:19.28" resultid="9523" heatid="11652" lane="9" entrytime="00:21:33.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:53.91" />
                    <SPLIT distance="200" swimtime="00:02:35.84" />
                    <SPLIT distance="250" swimtime="00:03:17.93" />
                    <SPLIT distance="300" swimtime="00:04:00.44" />
                    <SPLIT distance="350" swimtime="00:04:43.06" />
                    <SPLIT distance="400" swimtime="00:05:25.99" />
                    <SPLIT distance="450" swimtime="00:06:09.10" />
                    <SPLIT distance="500" swimtime="00:06:52.34" />
                    <SPLIT distance="550" swimtime="00:07:35.92" />
                    <SPLIT distance="600" swimtime="00:08:18.99" />
                    <SPLIT distance="650" swimtime="00:09:02.12" />
                    <SPLIT distance="700" swimtime="00:09:45.45" />
                    <SPLIT distance="750" swimtime="00:10:28.98" />
                    <SPLIT distance="800" swimtime="00:11:12.61" />
                    <SPLIT distance="850" swimtime="00:11:56.39" />
                    <SPLIT distance="900" swimtime="00:12:39.80" />
                    <SPLIT distance="950" swimtime="00:13:22.99" />
                    <SPLIT distance="1000" swimtime="00:14:06.28" />
                    <SPLIT distance="1050" swimtime="00:14:49.86" />
                    <SPLIT distance="1100" swimtime="00:15:33.72" />
                    <SPLIT distance="1150" swimtime="00:16:17.15" />
                    <SPLIT distance="1200" swimtime="00:17:00.86" />
                    <SPLIT distance="1250" swimtime="00:17:44.33" />
                    <SPLIT distance="1300" swimtime="00:18:28.33" />
                    <SPLIT distance="1350" swimtime="00:19:11.63" />
                    <SPLIT distance="1400" swimtime="00:19:55.02" />
                    <SPLIT distance="1450" swimtime="00:20:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="461" reactiontime="+116" swimtime="00:01:16.75" resultid="9524" heatid="11492" lane="1" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="500" reactiontime="+129" swimtime="00:02:55.03" resultid="9525" heatid="11503" lane="3" entrytime="00:02:51.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:18.44" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="552" reactiontime="+143" swimtime="00:00:32.67" resultid="9526" heatid="11535" lane="7" entrytime="00:00:33.72" />
                <RESULT eventid="6569" points="556" reactiontime="+137" swimtime="00:06:04.02" resultid="9527" heatid="11578" lane="7" entrytime="00:05:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:02:07.05" />
                    <SPLIT distance="200" swimtime="00:02:54.27" />
                    <SPLIT distance="250" swimtime="00:03:48.04" />
                    <SPLIT distance="300" swimtime="00:04:42.16" />
                    <SPLIT distance="350" swimtime="00:05:23.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="544" reactiontime="+103" swimtime="00:01:13.09" resultid="9528" heatid="11593" lane="1" entrytime="00:01:12.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="523" reactiontime="+135" swimtime="00:05:23.22" resultid="9529" heatid="11634" lane="5" entrytime="00:05:23.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                    <SPLIT distance="200" swimtime="00:02:34.88" />
                    <SPLIT distance="250" swimtime="00:03:17.09" />
                    <SPLIT distance="300" swimtime="00:03:59.34" />
                    <SPLIT distance="350" swimtime="00:04:42.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Spychalski" birthdate="1980-09-05" gender="M" nation="POL" license="102902700357" swrid="5337379" athleteid="9530">
              <RESULTS>
                <RESULT eventid="6203" points="522" reactiontime="+85" swimtime="00:20:37.75" resultid="9531" heatid="11652" lane="8" entrytime="00:21:01.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:53.09" />
                    <SPLIT distance="200" swimtime="00:02:34.00" />
                    <SPLIT distance="250" swimtime="00:03:15.59" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                    <SPLIT distance="350" swimtime="00:04:37.97" />
                    <SPLIT distance="400" swimtime="00:05:19.55" />
                    <SPLIT distance="450" swimtime="00:06:01.41" />
                    <SPLIT distance="500" swimtime="00:06:43.15" />
                    <SPLIT distance="550" swimtime="00:07:24.63" />
                    <SPLIT distance="600" swimtime="00:08:06.51" />
                    <SPLIT distance="650" swimtime="00:08:47.91" />
                    <SPLIT distance="700" swimtime="00:09:29.83" />
                    <SPLIT distance="750" swimtime="00:10:11.17" />
                    <SPLIT distance="800" swimtime="00:10:52.66" />
                    <SPLIT distance="850" swimtime="00:11:34.06" />
                    <SPLIT distance="900" swimtime="00:12:15.42" />
                    <SPLIT distance="950" swimtime="00:12:56.87" />
                    <SPLIT distance="1000" swimtime="00:13:38.29" />
                    <SPLIT distance="1050" swimtime="00:14:20.55" />
                    <SPLIT distance="1100" swimtime="00:15:02.60" />
                    <SPLIT distance="1150" swimtime="00:15:44.80" />
                    <SPLIT distance="1200" swimtime="00:16:27.07" />
                    <SPLIT distance="1250" swimtime="00:17:09.66" />
                    <SPLIT distance="1300" swimtime="00:17:52.84" />
                    <SPLIT distance="1350" swimtime="00:18:35.43" />
                    <SPLIT distance="1400" swimtime="00:19:18.33" />
                    <SPLIT distance="1450" swimtime="00:19:59.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8453" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Polowski" birthdate="2000-01-01" gender="M" nation="POL" swrid="4613096" athleteid="8452">
              <RESULTS>
                <RESULT eventid="6272" points="680" reactiontime="+72" swimtime="00:02:35.81" resultid="8454" heatid="11460" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="648" reactiontime="+66" swimtime="00:01:04.96" resultid="8455" heatid="11496" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="760" reactiontime="+72" swimtime="00:01:07.64" resultid="8456" heatid="11521" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="655" reactiontime="+67" swimtime="00:00:28.30" resultid="8457" heatid="11541" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="6704" points="817" reactiontime="+67" swimtime="00:00:30.22" resultid="8458" heatid="11623" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8459" heatid="11638" lane="8" entrytime="00:04:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8546" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-01-01" gender="F" nation="POL" athleteid="8545">
              <RESULTS>
                <RESULT eventid="6059" points="477" reactiontime="+79" swimtime="00:00:36.19" resultid="8547" heatid="11397" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="6145" points="374" reactiontime="+72" swimtime="00:13:31.64" resultid="8548" heatid="11644" lane="7" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:01:33.56" />
                    <SPLIT distance="150" swimtime="00:02:23.91" />
                    <SPLIT distance="200" swimtime="00:03:14.37" />
                    <SPLIT distance="250" swimtime="00:04:05.49" />
                    <SPLIT distance="300" swimtime="00:04:57.61" />
                    <SPLIT distance="350" swimtime="00:05:48.94" />
                    <SPLIT distance="400" swimtime="00:06:40.89" />
                    <SPLIT distance="450" swimtime="00:07:32.25" />
                    <SPLIT distance="500" swimtime="00:08:24.02" />
                    <SPLIT distance="550" swimtime="00:09:15.15" />
                    <SPLIT distance="600" swimtime="00:10:06.84" />
                    <SPLIT distance="650" swimtime="00:10:57.43" />
                    <SPLIT distance="700" swimtime="00:11:49.11" />
                    <SPLIT distance="750" swimtime="00:12:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="415" reactiontime="+74" swimtime="00:01:21.70" resultid="8549" heatid="11463" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="408" reactiontime="+77" swimtime="00:01:33.05" resultid="8550" heatid="11484" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="465" swimtime="00:00:40.20" resultid="8551" heatid="11525" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="6518" points="364" reactiontime="+73" swimtime="00:03:07.44" resultid="8552" heatid="11558" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="150" swimtime="00:02:19.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="505815" nation="POL" clubid="8589" name="Tm Barracuda Kalisz">
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Radomska" birthdate="1982-04-12" gender="F" nation="POL" athleteid="8590">
              <RESULTS>
                <RESULT eventid="6059" points="433" reactiontime="+84" swimtime="00:00:34.72" resultid="8591" heatid="11397" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="6145" reactiontime="+66" status="OTL" swimtime="00:00:00.00" resultid="8592" heatid="11643" lane="9" entrytime="00:12:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:27.11" />
                    <SPLIT distance="150" swimtime="00:02:15.22" />
                    <SPLIT distance="200" swimtime="00:03:04.72" />
                    <SPLIT distance="250" swimtime="00:03:53.70" />
                    <SPLIT distance="300" swimtime="00:04:43.26" />
                    <SPLIT distance="350" swimtime="00:05:33.37" />
                    <SPLIT distance="400" swimtime="00:06:23.64" />
                    <SPLIT distance="450" swimtime="00:07:14.86" />
                    <SPLIT distance="500" swimtime="00:08:05.38" />
                    <SPLIT distance="550" swimtime="00:08:54.93" />
                    <SPLIT distance="600" swimtime="00:09:44.74" />
                    <SPLIT distance="650" swimtime="00:10:34.40" />
                    <SPLIT distance="700" swimtime="00:11:23.79" />
                    <SPLIT distance="750" swimtime="00:12:15.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="410" reactiontime="+92" swimtime="00:01:18.67" resultid="8593" heatid="11463" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="357" reactiontime="+83" swimtime="00:01:36.00" resultid="8594" heatid="11483" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="409" swimtime="00:02:54.21" resultid="8595" heatid="11556" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:22.12" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="413" reactiontime="+104" swimtime="00:06:11.84" resultid="8596" heatid="11626" lane="9" entrytime="00:06:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:11.15" />
                    <SPLIT distance="200" swimtime="00:02:59.76" />
                    <SPLIT distance="250" swimtime="00:03:48.92" />
                    <SPLIT distance="300" swimtime="00:04:37.34" />
                    <SPLIT distance="350" swimtime="00:05:26.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="7859" name="Swim Masters Zlin">
          <ATHLETES>
            <ATHLETE firstname="Karel" lastname="Steker" birthdate="1981-08-12" gender="M" nation="CZE" swrid="5029799" athleteid="7860">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7861" heatid="11412" lane="3" entrytime="00:00:28.52" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7862" heatid="11430" lane="5" entrytime="00:02:43.94" />
                <RESULT eventid="6238" points="521" reactiontime="+70" swimtime="00:00:33.74" resultid="7863" heatid="11447" lane="6" entrytime="00:00:34.77" />
                <RESULT eventid="6374" points="465" reactiontime="+83" swimtime="00:02:42.63" resultid="7864" heatid="11504" lane="9" entrytime="00:02:45.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="536" reactiontime="+81" swimtime="00:00:30.92" resultid="7865" heatid="11537" lane="1" entrytime="00:00:30.79" />
                <RESULT eventid="6535" points="542" reactiontime="+79" swimtime="00:02:18.59" resultid="7866" heatid="11568" lane="1" entrytime="00:02:19.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="543" reactiontime="+71" swimtime="00:01:09.39" resultid="7867" heatid="11593" lane="4" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="512" reactiontime="+81" swimtime="00:05:00.75" resultid="7868" heatid="11635" lane="5" entrytime="00:05:05.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:49.32" />
                    <SPLIT distance="200" swimtime="00:02:29.08" />
                    <SPLIT distance="250" swimtime="00:03:08.54" />
                    <SPLIT distance="300" swimtime="00:03:47.82" />
                    <SPLIT distance="350" swimtime="00:04:26.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Prilucik" birthdate="1966-09-28" gender="M" nation="CZE" swrid="4934037" athleteid="7869">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7870" heatid="11409" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="6306" points="392" reactiontime="+86" swimtime="00:01:19.27" resultid="7871" heatid="11471" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="6704" status="DSQ" swimtime="00:00:00.00" resultid="7872" heatid="11617" lane="2" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8687" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Kuśmider" birthdate="1989-01-01" gender="M" nation="POL" athleteid="8686">
              <RESULTS>
                <RESULT eventid="6203" points="560" reactiontime="+90" swimtime="00:19:50.39" resultid="8688" heatid="11652" lane="7" entrytime="00:20:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                    <SPLIT distance="200" swimtime="00:02:32.14" />
                    <SPLIT distance="250" swimtime="00:03:11.97" />
                    <SPLIT distance="300" swimtime="00:03:52.05" />
                    <SPLIT distance="350" swimtime="00:04:31.60" />
                    <SPLIT distance="400" swimtime="00:05:11.38" />
                    <SPLIT distance="450" swimtime="00:05:51.27" />
                    <SPLIT distance="500" swimtime="00:06:31.54" />
                    <SPLIT distance="550" swimtime="00:07:10.71" />
                    <SPLIT distance="600" swimtime="00:07:50.29" />
                    <SPLIT distance="650" swimtime="00:08:30.16" />
                    <SPLIT distance="700" swimtime="00:09:10.40" />
                    <SPLIT distance="750" swimtime="00:09:50.58" />
                    <SPLIT distance="800" swimtime="00:10:30.65" />
                    <SPLIT distance="850" swimtime="00:11:10.69" />
                    <SPLIT distance="900" swimtime="00:11:50.68" />
                    <SPLIT distance="950" swimtime="00:12:30.82" />
                    <SPLIT distance="1000" swimtime="00:13:11.15" />
                    <SPLIT distance="1050" swimtime="00:13:51.13" />
                    <SPLIT distance="1100" swimtime="00:14:31.28" />
                    <SPLIT distance="1150" swimtime="00:15:11.10" />
                    <SPLIT distance="1200" swimtime="00:15:51.40" />
                    <SPLIT distance="1250" swimtime="00:16:31.30" />
                    <SPLIT distance="1300" swimtime="00:17:11.54" />
                    <SPLIT distance="1350" swimtime="00:17:52.02" />
                    <SPLIT distance="1400" swimtime="00:18:32.56" />
                    <SPLIT distance="1450" swimtime="00:19:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="434" reactiontime="+85" swimtime="00:01:04.74" resultid="8689" heatid="11474" lane="5" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="442" swimtime="00:02:19.82" resultid="8690" heatid="11567" lane="4" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8691" heatid="11635" lane="6" entrytime="00:05:08.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="11" clubid="8792" name="AZS AWF Katowice">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Sordyl" birthdate="1999-07-05" gender="M" nation="POL" license="100611700329" swrid="4292584" athleteid="8793">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="8794" heatid="11417" lane="3" entrytime="00:00:24.96" entrycourse="SCM" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="8795" heatid="11450" lane="3" entrytime="00:00:25.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8383" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Cygankiewicz" birthdate="1986-01-01" gender="M" nation="POL" athleteid="8382">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="8384" heatid="11408" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="8385" heatid="11472" lane="1" entrytime="00:01:12.00" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="8386" heatid="11535" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="8387" heatid="11565" lane="5" entrytime="00:02:45.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8388" heatid="11634" lane="0" entrytime="00:05:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6892" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Marciniszko" birthdate="1944-01-01" gender="M" nation="POL" swrid="4992778" athleteid="6891">
              <RESULTS>
                <RESULT eventid="6077" points="75" reactiontime="+123" swimtime="00:01:14.11" resultid="6893" heatid="11404" lane="7" entrytime="00:01:04.12" />
                <RESULT eventid="6238" points="110" reactiontime="+113" swimtime="00:01:15.99" resultid="6894" heatid="11444" lane="8" entrytime="00:01:17.91" />
                <RESULT eventid="6501" points="89" reactiontime="+117" swimtime="00:03:02.49" resultid="6895" heatid="11548" lane="5" entrytime="00:03:08.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="88" reactiontime="+117" swimtime="00:06:44.31" resultid="6896" heatid="11602" lane="1" entrytime="00:05:36.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.61" />
                    <SPLIT distance="100" swimtime="00:03:23.22" />
                    <SPLIT distance="150" swimtime="00:05:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="188" reactiontime="+87" swimtime="00:01:08.40" resultid="6897" heatid="11615" lane="6" entrytime="00:01:04.80" />
                <RESULT eventid="6433" points="128" reactiontime="+105" swimtime="00:02:51.86" resultid="6898" heatid="11515" lane="9" entrytime="00:02:48.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="112" reactiontime="+98" swimtime="00:06:45.46" resultid="6899" heatid="11456" lane="0" entrytime="00:05:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.12" />
                    <SPLIT distance="100" swimtime="00:03:09.32" />
                    <SPLIT distance="150" swimtime="00:04:57.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14814" nation="POL" region="14" clubid="9419" name="Stowarzyszenie Pływackie Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" license="514814700003" swrid="4992696" athleteid="9420">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="9421" heatid="11406" lane="7" entrytime="00:00:36.23" entrycourse="SCM" />
                <RESULT eventid="6203" points="384" reactiontime="+95" swimtime="00:27:37.42" resultid="9422" heatid="11654" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:02:31.23" />
                    <SPLIT distance="150" swimtime="00:03:26.41" />
                    <SPLIT distance="200" swimtime="00:04:21.55" />
                    <SPLIT distance="250" swimtime="00:05:18.70" />
                    <SPLIT distance="300" swimtime="00:06:14.65" />
                    <SPLIT distance="350" swimtime="00:07:10.01" />
                    <SPLIT distance="400" swimtime="00:08:05.71" />
                    <SPLIT distance="450" swimtime="00:09:01.87" />
                    <SPLIT distance="500" swimtime="00:09:57.51" />
                    <SPLIT distance="550" swimtime="00:10:54.38" />
                    <SPLIT distance="600" swimtime="00:11:50.06" />
                    <SPLIT distance="650" swimtime="00:12:46.15" />
                    <SPLIT distance="700" swimtime="00:13:41.90" />
                    <SPLIT distance="750" swimtime="00:14:37.34" />
                    <SPLIT distance="800" swimtime="00:15:34.32" />
                    <SPLIT distance="850" swimtime="00:16:30.79" />
                    <SPLIT distance="900" swimtime="00:17:28.44" />
                    <SPLIT distance="950" swimtime="00:18:23.85" />
                    <SPLIT distance="1000" swimtime="00:19:19.43" />
                    <SPLIT distance="1050" swimtime="00:20:15.91" />
                    <SPLIT distance="1100" swimtime="00:21:12.08" />
                    <SPLIT distance="1150" swimtime="00:22:07.07" />
                    <SPLIT distance="1200" swimtime="00:23:02.61" />
                    <SPLIT distance="1250" swimtime="00:23:58.46" />
                    <SPLIT distance="1300" swimtime="00:24:54.09" />
                    <SPLIT distance="1350" swimtime="00:25:52.34" />
                    <SPLIT distance="1400" swimtime="00:26:47.23" />
                    <SPLIT distance="1450" swimtime="00:27:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="471" reactiontime="+81" swimtime="00:00:42.82" resultid="9423" heatid="11446" lane="9" entrytime="00:00:42.92" entrycourse="SCM" />
                <RESULT eventid="6306" points="437" swimtime="00:01:20.49" resultid="9424" heatid="11470" lane="9" entrytime="00:01:24.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="388" reactiontime="+81" swimtime="00:01:39.16" resultid="9425" heatid="11547" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="415" reactiontime="+102" swimtime="00:03:06.80" resultid="9426" heatid="11562" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:18.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="382" reactiontime="+94" swimtime="00:03:37.16" resultid="9427" heatid="11601" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                    <SPLIT distance="100" swimtime="00:01:45.38" />
                    <SPLIT distance="150" swimtime="00:02:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="424" reactiontime="+82" swimtime="00:06:45.91" resultid="9428" heatid="11630" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:01:32.23" />
                    <SPLIT distance="150" swimtime="00:02:24.38" />
                    <SPLIT distance="200" swimtime="00:03:17.20" />
                    <SPLIT distance="250" swimtime="00:04:09.95" />
                    <SPLIT distance="300" swimtime="00:05:02.91" />
                    <SPLIT distance="350" swimtime="00:05:56.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Wilczęga" birthdate="1981-10-24" gender="M" nation="POL" license="514814700009" swrid="4992879" athleteid="9429">
              <RESULTS>
                <RESULT eventid="6077" points="651" swimtime="00:00:26.77" resultid="9430" heatid="11415" lane="4" entrytime="00:00:26.39" />
                <RESULT eventid="6306" points="655" reactiontime="+68" swimtime="00:00:59.03" resultid="9431" heatid="11477" lane="1" entrytime="00:00:59.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8533" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kowalski" birthdate="1996-01-01" gender="M" nation="POL" swrid="4282377" athleteid="8532">
              <RESULTS>
                <RESULT eventid="6077" points="692" reactiontime="+65" swimtime="00:00:25.82" resultid="8534" heatid="11416" lane="5" entrytime="00:00:25.80" />
                <RESULT eventid="6340" points="557" reactiontime="+63" swimtime="00:01:07.08" resultid="8535" heatid="11495" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="561" reactiontime="+56" swimtime="00:00:28.72" resultid="8536" heatid="11540" lane="1" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7102" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Rusłana" lastname="Dembecka" birthdate="1957-01-01" gender="F" nation="POL" athleteid="7101">
              <RESULTS>
                <RESULT eventid="6059" points="255" reactiontime="+112" swimtime="00:00:50.81" resultid="7103" heatid="11395" lane="7" />
                <RESULT eventid="6255" points="368" reactiontime="+116" swimtime="00:04:40.11" resultid="7104" heatid="11451" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.58" />
                    <SPLIT distance="100" swimtime="00:02:16.07" />
                    <SPLIT distance="150" swimtime="00:03:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="294" reactiontime="+106" swimtime="00:02:12.98" resultid="7105" heatid="11508" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="275" reactiontime="+103" swimtime="00:00:59.79" resultid="7106" heatid="11608" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9736" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Wypych" birthdate="1991-01-01" gender="M" nation="POL" swrid="4072458" athleteid="9735">
              <RESULTS>
                <RESULT eventid="6077" points="912" swimtime="00:00:22.82" resultid="9737" heatid="11419" lane="4" entrytime="00:00:21.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" clubid="7355" name="KS Masters Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Zygmunt" lastname="Pawlaczek" birthdate="1949-05-26" gender="M" nation="POL" athleteid="7409">
              <RESULTS>
                <RESULT eventid="6077" points="393" reactiontime="+105" swimtime="00:00:38.76" resultid="7410" heatid="11405" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="6169" points="345" reactiontime="+112" swimtime="00:16:20.87" resultid="7411" heatid="11648" lane="7" entrytime="00:16:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:44.84" />
                    <SPLIT distance="150" swimtime="00:02:44.01" />
                    <SPLIT distance="200" swimtime="00:03:43.99" />
                    <SPLIT distance="250" swimtime="00:04:46.57" />
                    <SPLIT distance="300" swimtime="00:05:50.25" />
                    <SPLIT distance="350" swimtime="00:06:54.09" />
                    <SPLIT distance="400" swimtime="00:07:56.93" />
                    <SPLIT distance="450" swimtime="00:08:59.88" />
                    <SPLIT distance="500" swimtime="00:10:03.48" />
                    <SPLIT distance="550" swimtime="00:11:07.51" />
                    <SPLIT distance="600" swimtime="00:12:10.66" />
                    <SPLIT distance="650" swimtime="00:13:15.90" />
                    <SPLIT distance="700" swimtime="00:14:19.86" />
                    <SPLIT distance="750" swimtime="00:15:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="380" reactiontime="+100" swimtime="00:04:15.71" resultid="7412" heatid="11456" lane="8" entrytime="00:04:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.75" />
                    <SPLIT distance="100" swimtime="00:02:00.74" />
                    <SPLIT distance="150" swimtime="00:03:07.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="395" reactiontime="+98" swimtime="00:01:28.06" resultid="7413" heatid="11469" lane="1" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="399" reactiontime="+116" swimtime="00:01:51.92" resultid="7414" heatid="11516" lane="0" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7415" heatid="11563" lane="8" entrytime="00:03:50.00" entrycourse="SCM" />
                <RESULT eventid="6704" points="390" reactiontime="+104" swimtime="00:00:48.60" resultid="7416" heatid="11616" lane="7" entrytime="00:00:48.00" entrycourse="SCM" />
                <RESULT eventid="6738" points="329" reactiontime="+116" swimtime="00:07:54.62" resultid="7417" heatid="11630" lane="4" entrytime="00:08:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                    <SPLIT distance="100" swimtime="00:01:46.11" />
                    <SPLIT distance="150" swimtime="00:02:45.23" />
                    <SPLIT distance="200" swimtime="00:03:47.14" />
                    <SPLIT distance="250" swimtime="00:04:49.95" />
                    <SPLIT distance="300" swimtime="00:05:53.56" />
                    <SPLIT distance="350" swimtime="00:06:55.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Kawula" birthdate="1941-10-02" gender="F" nation="POL" athleteid="7362">
              <RESULTS>
                <RESULT eventid="6059" points="94" swimtime="00:01:32.59" resultid="7363" heatid="11395" lane="9" />
                <RESULT eventid="6289" points="85" swimtime="00:03:21.85" resultid="7364" heatid="11461" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="51" swimtime="00:04:44.54" resultid="7365" heatid="11509" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:19.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="46" swimtime="00:02:17.11" resultid="7366" heatid="11608" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Jawor" birthdate="1947-04-23" gender="M" nation="POL" swrid="4754745" athleteid="7402">
              <RESULTS>
                <RESULT eventid="6238" points="215" reactiontime="+125" swimtime="00:01:00.73" resultid="7403" heatid="11443" lane="4" />
                <RESULT eventid="6340" points="226" reactiontime="+90" swimtime="00:02:16.99" resultid="7404" heatid="11488" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="278" reactiontime="+88" swimtime="00:02:12.79" resultid="7405" heatid="11514" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="202" reactiontime="+101" swimtime="00:02:19.05" resultid="7406" heatid="11548" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="282" reactiontime="+123" swimtime="00:04:34.47" resultid="7407" heatid="11601" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.26" />
                    <SPLIT distance="100" swimtime="00:02:14.32" />
                    <SPLIT distance="150" swimtime="00:03:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="274" reactiontime="+88" swimtime="00:01:00.31" resultid="7408" heatid="11614" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Regina" lastname="Mładszew" birthdate="1952-07-15" gender="F" nation="POL" athleteid="7367">
              <RESULTS>
                <RESULT eventid="6059" points="97" reactiontime="+126" swimtime="00:01:12.36" resultid="7368" heatid="11394" lane="5" />
                <RESULT eventid="6220" points="100" reactiontime="+149" swimtime="00:01:29.99" resultid="7369" heatid="11438" lane="4" />
                <RESULT eventid="6323" points="91" swimtime="00:03:05.35" resultid="7370" heatid="11480" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="64" swimtime="00:01:31.66" resultid="7371" heatid="11523" lane="2" />
                <RESULT eventid="6484" points="134" reactiontime="+134" swimtime="00:02:54.06" resultid="7372" heatid="11544" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="175" reactiontime="+70" swimtime="00:05:53.09" resultid="7373" heatid="11598" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.57" />
                    <SPLIT distance="100" swimtime="00:02:55.85" />
                    <SPLIT distance="150" swimtime="00:04:26.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="114" swimtime="00:01:28.92" resultid="7374" heatid="11607" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gizela" lastname="Wójcik" birthdate="1949-11-16" gender="F" nation="POL" athleteid="7380">
              <RESULTS>
                <RESULT eventid="6059" points="111" swimtime="00:01:09.31" resultid="7381" heatid="11393" lane="4" />
                <RESULT eventid="6220" points="211" reactiontime="+147" swimtime="00:01:10.17" resultid="7382" heatid="11438" lane="8" />
                <RESULT eventid="6255" points="252" swimtime="00:05:37.21" resultid="7383" heatid="11451" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.73" />
                    <SPLIT distance="100" swimtime="00:02:42.73" />
                    <SPLIT distance="150" swimtime="00:04:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="226" swimtime="00:02:39.34" resultid="7384" heatid="11509" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach." eventid="6484" reactiontime="+120" status="DSQ" swimtime="00:00:00.00" resultid="7385" heatid="11544" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="182" swimtime="00:01:16.06" resultid="7386" heatid="11607" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Ołpiński" birthdate="1991-04-26" gender="M" nation="POL" swrid="4217107" athleteid="7356">
              <RESULTS>
                <RESULT eventid="6077" points="535" reactiontime="+75" swimtime="00:00:27.25" resultid="7357" heatid="11416" lane="8" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="6111" points="398" reactiontime="+82" swimtime="00:02:40.52" resultid="7358" heatid="11428" lane="5" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:02:01.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="484" reactiontime="+82" swimtime="00:01:02.44" resultid="7359" heatid="11471" lane="5" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="490" swimtime="00:00:28.99" resultid="7360" heatid="11538" lane="8" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="6535" points="381" reactiontime="+78" swimtime="00:02:26.83" resultid="7361" heatid="11565" lane="0" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:48.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Zając" birthdate="1946-01-02" gender="M" nation="POL" athleteid="7394">
              <RESULTS>
                <RESULT eventid="6077" points="160" swimtime="00:00:57.59" resultid="7395" heatid="11403" lane="7" />
                <RESULT eventid="6238" points="116" reactiontime="+96" swimtime="00:01:14.61" resultid="7396" heatid="11443" lane="1" />
                <RESULT eventid="6306" points="145" swimtime="00:02:15.22" resultid="7397" heatid="11467" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="174" swimtime="00:02:35.39" resultid="7398" heatid="11514" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="96" reactiontime="+116" swimtime="00:02:58.11" resultid="7399" heatid="11548" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="7400" heatid="11601" lane="6" />
                <RESULT eventid="6704" points="153" swimtime="00:01:13.21" resultid="7401" heatid="11614" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janina" lastname="Zając" birthdate="1946-08-16" gender="F" nation="POL" athleteid="7387">
              <RESULTS>
                <RESULT eventid="6059" points="114" swimtime="00:01:11.15" resultid="7388" heatid="11395" lane="0" />
                <RESULT eventid="6220" points="140" reactiontime="+130" swimtime="00:01:23.99" resultid="7389" heatid="11438" lane="6" />
                <RESULT eventid="6289" points="96" swimtime="00:02:52.20" resultid="7390" heatid="11461" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="150" reactiontime="+95" swimtime="00:02:55.97" resultid="7391" heatid="11543" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="161" reactiontime="+95" swimtime="00:06:11.81" resultid="7392" heatid="11598" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.61" />
                    <SPLIT distance="100" swimtime="00:02:59.21" />
                    <SPLIT distance="150" swimtime="00:04:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="71" swimtime="00:01:53.80" resultid="7393" heatid="11608" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pavlo" lastname="Vechirko" birthdate="1968-01-02" gender="M" nation="POL" athleteid="7418">
              <RESULTS>
                <RESULT eventid="6433" points="493" reactiontime="+90" swimtime="00:01:24.96" resultid="7419" heatid="11518" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="435" reactiontime="+94" swimtime="00:01:19.79" resultid="7420" heatid="11551" lane="9" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="534" swimtime="00:00:37.90" resultid="7421" heatid="11619" lane="4" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Józefa" lastname="Wołoszczuk" birthdate="1953-01-23" gender="F" nation="POL" athleteid="7375">
              <RESULTS>
                <RESULT eventid="6220" points="179" reactiontime="+86" swimtime="00:01:10.93" resultid="7376" heatid="11438" lane="1" />
                <RESULT eventid="6289" points="135" swimtime="00:02:18.22" resultid="7377" heatid="11461" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="182" reactiontime="+94" swimtime="00:02:34.37" resultid="7378" heatid="11544" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="191" reactiontime="+92" swimtime="00:05:26.93" resultid="7379" heatid="11598" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.30" />
                    <SPLIT distance="100" swimtime="00:02:43.59" />
                    <SPLIT distance="150" swimtime="00:04:07.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6820" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Łopuszyński" birthdate="1969-01-01" gender="M" nation="POL" athleteid="6819">
              <RESULTS>
                <RESULT eventid="6111" points="184" reactiontime="+89" swimtime="00:03:51.92" resultid="6821" heatid="11427" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:53.24" />
                    <SPLIT distance="150" swimtime="00:02:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="209" reactiontime="+110" swimtime="00:03:53.97" resultid="6822" heatid="11501" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.12" />
                    <SPLIT distance="100" swimtime="00:01:50.17" />
                    <SPLIT distance="150" swimtime="00:02:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="159" reactiontime="+115" swimtime="00:00:49.39" resultid="6823" heatid="11532" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="6569" points="219" reactiontime="+104" swimtime="00:08:16.61" resultid="6824" heatid="11576" lane="6" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                    <SPLIT distance="100" swimtime="00:01:51.76" />
                    <SPLIT distance="150" swimtime="00:02:57.70" />
                    <SPLIT distance="200" swimtime="00:04:01.99" />
                    <SPLIT distance="250" swimtime="00:05:11.75" />
                    <SPLIT distance="300" swimtime="00:06:23.16" />
                    <SPLIT distance="350" swimtime="00:07:19.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="172" swimtime="00:01:47.14" resultid="6825" heatid="11590" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" clubid="7030" name="Motyl Masters">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Lorkowski" birthdate="1960-02-27" gender="M" nation="POL" swrid="4992838" athleteid="7031">
              <RESULTS>
                <RESULT eventid="6077" points="636" swimtime="00:00:31.20" resultid="7032" heatid="11410" lane="9" entrytime="00:00:31.99" />
                <RESULT eventid="6111" points="624" reactiontime="+83" swimtime="00:02:58.93" resultid="7033" heatid="11429" lane="3" entrytime="00:02:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:24.85" />
                    <SPLIT distance="150" swimtime="00:02:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="629" reactiontime="+87" swimtime="00:01:09.84" resultid="7034" heatid="11472" lane="3" entrytime="00:01:10.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="508" reactiontime="+92" swimtime="00:03:20.13" resultid="7035" heatid="11502" lane="1" entrytime="00:03:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="150" swimtime="00:02:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="645" reactiontime="+90" swimtime="00:02:37.91" resultid="7036" heatid="11566" lane="6" entrytime="00:02:39.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="594" reactiontime="+95" swimtime="00:06:25.28" resultid="7037" heatid="11577" lane="6" entrytime="00:06:29.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:02:21.92" />
                    <SPLIT distance="200" swimtime="00:03:08.75" />
                    <SPLIT distance="250" swimtime="00:04:04.63" />
                    <SPLIT distance="300" swimtime="00:05:00.24" />
                    <SPLIT distance="350" swimtime="00:05:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="680" reactiontime="+94" swimtime="00:02:58.49" resultid="7038" heatid="11604" lane="9" entrytime="00:03:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:27.11" />
                    <SPLIT distance="150" swimtime="00:02:13.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="621" reactiontime="+92" swimtime="00:05:41.33" resultid="7039" heatid="11633" lane="3" entrytime="00:05:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:03.52" />
                    <SPLIT distance="200" swimtime="00:02:48.06" />
                    <SPLIT distance="250" swimtime="00:03:32.41" />
                    <SPLIT distance="300" swimtime="00:04:16.66" />
                    <SPLIT distance="350" swimtime="00:04:59.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Pawłowski" birthdate="1977-06-26" gender="M" nation="POL" swrid="4992839" athleteid="7055">
              <RESULTS>
                <RESULT eventid="6169" points="494" reactiontime="+87" swimtime="00:10:57.20" resultid="7056" heatid="11646" lane="7" entrytime="00:11:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                    <SPLIT distance="150" swimtime="00:01:55.27" />
                    <SPLIT distance="200" swimtime="00:02:36.76" />
                    <SPLIT distance="250" swimtime="00:03:18.00" />
                    <SPLIT distance="300" swimtime="00:03:59.50" />
                    <SPLIT distance="350" swimtime="00:04:40.90" />
                    <SPLIT distance="400" swimtime="00:05:22.56" />
                    <SPLIT distance="450" swimtime="00:06:04.27" />
                    <SPLIT distance="500" swimtime="00:06:45.82" />
                    <SPLIT distance="550" swimtime="00:07:28.14" />
                    <SPLIT distance="600" swimtime="00:08:10.73" />
                    <SPLIT distance="650" swimtime="00:08:52.82" />
                    <SPLIT distance="700" swimtime="00:09:34.80" />
                    <SPLIT distance="750" swimtime="00:10:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="606" reactiontime="+80" swimtime="00:00:32.92" resultid="7057" heatid="11447" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="6272" points="545" reactiontime="+80" swimtime="00:03:00.72" resultid="7058" heatid="11458" lane="8" entrytime="00:03:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                    <SPLIT distance="150" swimtime="00:02:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="569" reactiontime="+85" swimtime="00:01:11.66" resultid="7059" heatid="11551" lane="2" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="530" reactiontime="+84" swimtime="00:05:57.11" resultid="7060" heatid="11578" lane="0" entrytime="00:06:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:02:12.27" />
                    <SPLIT distance="200" swimtime="00:02:57.47" />
                    <SPLIT distance="250" swimtime="00:03:47.20" />
                    <SPLIT distance="300" swimtime="00:04:36.67" />
                    <SPLIT distance="350" swimtime="00:05:16.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="539" reactiontime="+78" swimtime="00:02:41.60" resultid="7061" heatid="11605" lane="0" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:02:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7062" heatid="11620" lane="8" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Przybylski" birthdate="1967-03-12" gender="M" nation="POL" athleteid="7047">
              <RESULTS>
                <RESULT eventid="6077" points="723" reactiontime="+83" swimtime="00:00:28.99" resultid="7048" heatid="11412" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7049" heatid="11474" lane="4" entrytime="00:01:04.01" />
                <RESULT eventid="6374" points="366" swimtime="00:03:14.22" resultid="7050" heatid="11503" lane="9" entrytime="00:03:05.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:20.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="630" reactiontime="+89" swimtime="00:00:32.71" resultid="7051" heatid="11536" lane="0" entrytime="00:00:32.51" />
                <RESULT eventid="6501" points="510" reactiontime="+76" swimtime="00:01:21.02" resultid="7052" heatid="11550" lane="4" entrytime="00:01:18.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="7053" heatid="11592" lane="1" entrytime="00:01:20.07" />
                <RESULT eventid="6670" points="530" reactiontime="+82" swimtime="00:02:56.94" resultid="7054" heatid="11604" lane="7" entrytime="00:02:55.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:11.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" swrid="4791744" athleteid="7040">
              <RESULTS>
                <RESULT eventid="6111" points="767" reactiontime="+79" swimtime="00:02:24.61" resultid="7041" heatid="11433" lane="2" entrytime="00:02:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="762" reactiontime="+79" swimtime="00:01:05.64" resultid="7042" heatid="11496" lane="3" entrytime="00:01:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="713" reactiontime="+74" swimtime="00:00:28.74" resultid="7043" heatid="11540" lane="5" entrytime="00:00:27.69" />
                <RESULT eventid="6535" points="731" reactiontime="+83" swimtime="00:02:07.31" resultid="7044" heatid="11570" lane="1" entrytime="00:02:05.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="796" reactiontime="+66" swimtime="00:01:03.16" resultid="7045" heatid="11596" lane="6" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="702" swimtime="00:04:36.60" resultid="7046" heatid="11638" lane="0" entrytime="00:04:31.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:42.00" />
                    <SPLIT distance="200" swimtime="00:02:17.46" />
                    <SPLIT distance="250" swimtime="00:02:52.68" />
                    <SPLIT distance="300" swimtime="00:03:27.79" />
                    <SPLIT distance="350" swimtime="00:04:02.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+83" swimtime="00:01:57.27" resultid="9837" heatid="11583" lane="5" entrytime="00:01:58.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="150" swimtime="00:01:30.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7047" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="7055" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="7031" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="7040" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+79" swimtime="00:02:13.41" resultid="9838" heatid="12331" lane="6" entrytime="00:02:07.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:41.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7047" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="7055" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="7040" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="7031" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7911" name="Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" swrid="4302086" athleteid="7912">
              <RESULTS>
                <RESULT eventid="6077" points="194" reactiontime="+115" swimtime="00:00:55.34" resultid="7913" heatid="11404" lane="3" entrytime="00:00:52.50" />
                <RESULT eventid="6111" points="212" swimtime="00:05:46.18" resultid="7914" heatid="11427" lane="1" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.07" />
                    <SPLIT distance="100" swimtime="00:03:06.00" />
                    <SPLIT distance="150" swimtime="00:04:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="203" reactiontime="+110" swimtime="00:01:05.71" resultid="7915" heatid="11444" lane="7" entrytime="00:01:01.50" />
                <RESULT eventid="6340" points="235" reactiontime="+119" swimtime="00:02:23.35" resultid="7916" heatid="11488" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="310" swimtime="00:02:23.11" resultid="7917" heatid="11515" lane="8" entrytime="00:02:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="214" reactiontime="+107" swimtime="00:02:33.69" resultid="7918" heatid="11548" lane="4" entrytime="00:02:15.00" />
                <RESULT eventid="6704" points="403" swimtime="00:00:58.16" resultid="7919" heatid="11615" lane="4" entrytime="00:00:57.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Heisler" birthdate="1951-01-01" gender="F" nation="POL" swrid="4191114" athleteid="7930">
              <RESULTS>
                <RESULT eventid="6059" points="376" reactiontime="+90" swimtime="00:00:46.19" resultid="7931" heatid="11396" lane="6" entrytime="00:00:44.50" />
                <RESULT eventid="6220" status="DNS" swimtime="00:00:00.00" resultid="7932" heatid="11439" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="6323" points="279" reactiontime="+84" swimtime="00:02:07.61" resultid="7933" heatid="11482" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="325" swimtime="00:02:21.18" resultid="7934" heatid="11510" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="169" swimtime="00:01:06.25" resultid="7935" heatid="11524" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="6687" points="329" reactiontime="+94" swimtime="00:01:02.50" resultid="7936" heatid="11609" lane="6" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gorbaczow" birthdate="1958-01-01" gender="M" nation="POL" swrid="4191113" athleteid="7920">
              <RESULTS>
                <RESULT eventid="6077" points="694" reactiontime="+85" swimtime="00:00:30.31" resultid="7921" heatid="11409" lane="2" entrytime="00:00:32.20" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="7922" heatid="11447" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="6306" points="650" reactiontime="+89" swimtime="00:01:09.08" resultid="7923" heatid="11473" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="727" reactiontime="+99" swimtime="00:00:32.41" resultid="7924" heatid="11536" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7925" heatid="11566" lane="7" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Gorbaczow" birthdate="1987-01-01" gender="M" nation="POL" athleteid="7926">
              <RESULTS>
                <RESULT eventid="6077" points="306" swimtime="00:00:32.66" resultid="7927" heatid="11407" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="6306" points="275" reactiontime="+94" swimtime="00:01:15.88" resultid="7928" heatid="11471" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="220" reactiontime="+101" swimtime="00:00:39.09" resultid="7929" heatid="11534" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7013" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Wilmowicz" birthdate="1979-01-01" gender="M" nation="POL" athleteid="7012">
              <RESULTS>
                <RESULT eventid="6077" points="522" swimtime="00:00:28.81" resultid="7014" heatid="11411" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="6203" points="583" reactiontime="+76" swimtime="00:19:53.11" resultid="7015" heatid="11652" lane="1" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                    <SPLIT distance="200" swimtime="00:02:25.52" />
                    <SPLIT distance="250" swimtime="00:03:04.47" />
                    <SPLIT distance="300" swimtime="00:03:43.62" />
                    <SPLIT distance="350" swimtime="00:04:22.94" />
                    <SPLIT distance="400" swimtime="00:05:02.60" />
                    <SPLIT distance="450" swimtime="00:05:42.22" />
                    <SPLIT distance="500" swimtime="00:06:21.97" />
                    <SPLIT distance="550" swimtime="00:07:01.49" />
                    <SPLIT distance="600" swimtime="00:07:41.05" />
                    <SPLIT distance="650" swimtime="00:08:20.67" />
                    <SPLIT distance="700" swimtime="00:09:00.50" />
                    <SPLIT distance="750" swimtime="00:09:40.46" />
                    <SPLIT distance="800" swimtime="00:10:20.74" />
                    <SPLIT distance="850" swimtime="00:11:00.85" />
                    <SPLIT distance="900" swimtime="00:11:40.92" />
                    <SPLIT distance="950" swimtime="00:12:22.34" />
                    <SPLIT distance="1000" swimtime="00:13:02.47" />
                    <SPLIT distance="1050" swimtime="00:13:42.99" />
                    <SPLIT distance="1100" swimtime="00:14:23.59" />
                    <SPLIT distance="1150" swimtime="00:15:05.00" />
                    <SPLIT distance="1200" swimtime="00:15:45.20" />
                    <SPLIT distance="1250" swimtime="00:16:26.31" />
                    <SPLIT distance="1300" swimtime="00:17:08.23" />
                    <SPLIT distance="1350" swimtime="00:17:49.10" />
                    <SPLIT distance="1400" swimtime="00:18:30.27" />
                    <SPLIT distance="1450" swimtime="00:19:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="547" reactiontime="+78" swimtime="00:01:02.69" resultid="7016" heatid="11474" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z2 - Pływak pokonał jednym stylem więcej niż 1 dystansu." eventid="6340" reactiontime="+75" status="DSQ" swimtime="00:00:00.00" resultid="7017" heatid="11494" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="550" reactiontime="+83" swimtime="00:02:17.93" resultid="7018" heatid="11568" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="529" reactiontime="+85" swimtime="00:04:57.42" resultid="7019" heatid="11636" lane="8" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:09.92" />
                    <SPLIT distance="150" swimtime="00:01:47.65" />
                    <SPLIT distance="200" swimtime="00:02:26.05" />
                    <SPLIT distance="250" swimtime="00:03:04.94" />
                    <SPLIT distance="300" swimtime="00:03:43.88" />
                    <SPLIT distance="350" swimtime="00:04:21.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6914" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Pietruszewski-Gil" birthdate="1986-01-01" gender="M" nation="POL" athleteid="6913">
              <RESULTS>
                <RESULT eventid="6077" points="366" reactiontime="+90" swimtime="00:00:30.79" resultid="6915" heatid="11411" lane="6" entrytime="00:00:29.99" />
                <RESULT eventid="6306" points="374" swimtime="00:01:08.47" resultid="6916" heatid="11473" lane="4" entrytime="00:01:06.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9738" name="5 Styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-01-01" gender="M" nation="POL" swrid="4273597" athleteid="9759">
              <RESULTS>
                <RESULT eventid="6111" points="668" swimtime="00:02:15.10" resultid="9760" heatid="11433" lane="1" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                    <SPLIT distance="150" swimtime="00:01:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="857" swimtime="00:02:27.93" resultid="9761" heatid="11460" lane="1" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="705" reactiontime="+67" swimtime="00:01:01.77" resultid="9762" heatid="11496" lane="8" entrytime="00:01:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="780" reactiontime="+68" swimtime="00:01:06.63" resultid="9763" heatid="11520" lane="3" entrytime="00:01:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="749" reactiontime="+70" swimtime="00:04:53.90" resultid="9764" heatid="11579" lane="2" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                    <SPLIT distance="200" swimtime="00:02:23.99" />
                    <SPLIT distance="250" swimtime="00:03:03.57" />
                    <SPLIT distance="300" swimtime="00:03:44.75" />
                    <SPLIT distance="350" swimtime="00:04:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="615" reactiontime="+75" swimtime="00:01:01.88" resultid="9765" heatid="11595" lane="7" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="722" swimtime="00:00:30.99" resultid="9766" heatid="11622" lane="8" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Kozyra" birthdate="1959-12-25" gender="M" nation="POL" athleteid="9803">
              <RESULTS>
                <RESULT eventid="6077" points="378" reactiontime="+92" swimtime="00:00:37.10" resultid="9804" heatid="11407" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="6111" points="320" reactiontime="+98" swimtime="00:03:43.45" resultid="9805" heatid="11427" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:44.00" />
                    <SPLIT distance="150" swimtime="00:02:53.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="333" reactiontime="+93" swimtime="00:01:38.50" resultid="9806" heatid="11489" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="318" reactiontime="+88" swimtime="00:00:42.70" resultid="9807" heatid="11533" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="6535" points="368" reactiontime="+101" swimtime="00:03:10.40" resultid="9808" heatid="11563" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:30.47" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wziątek" birthdate="1988-01-01" gender="M" nation="POL" athleteid="9739">
              <RESULTS>
                <RESULT eventid="6169" reactiontime="+81" status="OTL" swimtime="00:00:00.00" resultid="9740" heatid="11647" lane="6" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:19.25" />
                    <SPLIT distance="150" swimtime="00:02:04.80" />
                    <SPLIT distance="200" swimtime="00:02:51.11" />
                    <SPLIT distance="250" swimtime="00:03:37.83" />
                    <SPLIT distance="300" swimtime="00:04:25.25" />
                    <SPLIT distance="350" swimtime="00:05:13.29" />
                    <SPLIT distance="400" swimtime="00:06:02.11" />
                    <SPLIT distance="450" swimtime="00:06:51.82" />
                    <SPLIT distance="500" swimtime="00:07:41.63" />
                    <SPLIT distance="550" swimtime="00:08:30.86" />
                    <SPLIT distance="600" swimtime="00:09:20.79" />
                    <SPLIT distance="650" swimtime="00:10:11.01" />
                    <SPLIT distance="700" swimtime="00:11:00.19" />
                    <SPLIT distance="750" swimtime="00:11:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="349" reactiontime="+84" swimtime="00:01:09.60" resultid="9741" heatid="11471" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="323" reactiontime="+86" swimtime="00:02:35.20" resultid="9742" heatid="11566" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:53.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="296" reactiontime="+86" swimtime="00:01:18.92" resultid="9743" heatid="11592" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="371" reactiontime="+78" swimtime="00:05:34.12" resultid="9744" heatid="11632" lane="5" entrytime="00:06:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:56.87" />
                    <SPLIT distance="200" swimtime="00:02:39.59" />
                    <SPLIT distance="250" swimtime="00:03:23.53" />
                    <SPLIT distance="300" swimtime="00:04:07.91" />
                    <SPLIT distance="350" swimtime="00:04:52.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Cieślak" birthdate="1992-01-01" gender="M" nation="POL" swrid="4071989" athleteid="9780">
              <RESULTS>
                <RESULT eventid="6077" points="937" reactiontime="+66" swimtime="00:00:22.61" resultid="9781" heatid="11419" lane="3" entrytime="00:00:22.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6238" points="1167" reactiontime="+66" swimtime="00:00:25.17" resultid="9782" heatid="11450" lane="5" entrytime="00:00:25.50" />
                <RESULT eventid="6467" points="904" reactiontime="+64" swimtime="00:00:23.65" resultid="9783" heatid="11542" lane="4" entrytime="00:00:23.12" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9784" heatid="11597" lane="5" entrytime="00:00:52.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-01-10" gender="M" nation="POL" athleteid="9752">
              <RESULTS>
                <RESULT eventid="6077" points="363" reactiontime="+82" swimtime="00:00:32.51" resultid="9753" heatid="11408" lane="5" entrytime="00:00:33.10" />
                <RESULT eventid="6306" points="342" reactiontime="+79" swimtime="00:01:13.28" resultid="9754" heatid="11471" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="333" swimtime="00:01:26.30" resultid="9755" heatid="11490" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="369" reactiontime="+85" swimtime="00:01:28.61" resultid="9756" heatid="11518" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="343" reactiontime="+83" swimtime="00:02:41.46" resultid="9757" heatid="11565" lane="7" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:01:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="371" reactiontime="+78" swimtime="00:00:40.47" resultid="9758" heatid="11618" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Wąsiakowska" birthdate="1990-01-01" gender="F" nation="POL" swrid="4112407" athleteid="9812">
              <RESULTS>
                <RESULT eventid="6059" status="DNS" swimtime="00:00:00.00" resultid="9813" heatid="11400" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Dzikiewicz" birthdate="1990-11-11" gender="M" nation="POL" athleteid="9794">
              <RESULTS>
                <RESULT eventid="6077" points="321" reactiontime="+90" swimtime="00:00:32.30" resultid="9795" heatid="11406" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="6306" points="245" reactiontime="+93" swimtime="00:01:18.28" resultid="9796" heatid="11469" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łatkowska" birthdate="1965-01-01" gender="F" nation="POL" athleteid="9785">
              <RESULTS>
                <RESULT eventid="6059" points="345" swimtime="00:00:40.96" resultid="9786" heatid="11396" lane="4" entrytime="00:00:41.99" />
                <RESULT eventid="6186" points="358" reactiontime="+91" swimtime="00:27:49.28" resultid="9787" heatid="11651" lane="5" entrytime="00:28:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:39.38" />
                    <SPLIT distance="150" swimtime="00:02:33.77" />
                    <SPLIT distance="200" swimtime="00:03:29.47" />
                    <SPLIT distance="250" swimtime="00:04:25.83" />
                    <SPLIT distance="300" swimtime="00:05:21.67" />
                    <SPLIT distance="350" swimtime="00:06:18.43" />
                    <SPLIT distance="400" swimtime="00:07:15.11" />
                    <SPLIT distance="450" swimtime="00:08:11.48" />
                    <SPLIT distance="500" swimtime="00:09:08.11" />
                    <SPLIT distance="550" swimtime="00:10:05.01" />
                    <SPLIT distance="600" swimtime="00:11:02.14" />
                    <SPLIT distance="650" swimtime="00:11:58.49" />
                    <SPLIT distance="700" swimtime="00:12:54.05" />
                    <SPLIT distance="750" swimtime="00:13:51.41" />
                    <SPLIT distance="800" swimtime="00:14:47.71" />
                    <SPLIT distance="850" swimtime="00:15:44.59" />
                    <SPLIT distance="900" swimtime="00:16:41.48" />
                    <SPLIT distance="950" swimtime="00:17:38.39" />
                    <SPLIT distance="1000" swimtime="00:18:35.18" />
                    <SPLIT distance="1050" swimtime="00:19:32.29" />
                    <SPLIT distance="1100" swimtime="00:20:28.66" />
                    <SPLIT distance="1150" swimtime="00:21:24.77" />
                    <SPLIT distance="1200" swimtime="00:22:20.40" />
                    <SPLIT distance="1250" swimtime="00:23:16.25" />
                    <SPLIT distance="1300" swimtime="00:24:12.55" />
                    <SPLIT distance="1350" swimtime="00:25:09.06" />
                    <SPLIT distance="1400" swimtime="00:26:05.16" />
                    <SPLIT distance="1450" swimtime="00:26:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="281" reactiontime="+84" swimtime="00:00:51.65" resultid="9788" heatid="11439" lane="6" entrytime="00:00:52.06" />
                <RESULT eventid="6323" points="317" reactiontime="+86" swimtime="00:01:46.88" resultid="9789" heatid="11482" lane="3" entrytime="00:01:47.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="232" reactiontime="+84" swimtime="00:00:51.98" resultid="9790" heatid="11524" lane="2" entrytime="00:00:51.13" />
                <RESULT eventid="6518" points="303" reactiontime="+104" swimtime="00:03:25.12" resultid="9791" heatid="11556" lane="7" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:38.73" />
                    <SPLIT distance="150" swimtime="00:02:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="9792" heatid="11610" lane="9" entrytime="00:00:55.60" />
                <RESULT eventid="6721" points="284" reactiontime="+89" swimtime="00:07:23.25" resultid="9793" heatid="11625" lane="7" entrytime="00:07:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:42.68" />
                    <SPLIT distance="150" swimtime="00:02:38.60" />
                    <SPLIT distance="200" swimtime="00:03:35.75" />
                    <SPLIT distance="250" swimtime="00:04:33.66" />
                    <SPLIT distance="300" swimtime="00:05:30.93" />
                    <SPLIT distance="350" swimtime="00:06:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Dubiel" birthdate="1987-01-01" gender="M" nation="POL" swrid="4060947" athleteid="9770">
              <RESULTS>
                <RESULT eventid="6238" points="755" reactiontime="+64" swimtime="00:00:26.88" resultid="9771" heatid="11450" lane="8" entrytime="00:00:26.99" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6306" points="829" reactiontime="+75" swimtime="00:00:52.54" resultid="9772" heatid="11479" lane="8" entrytime="00:00:53.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="861" reactiontime="+72" swimtime="00:00:58.78" resultid="9773" heatid="11553" lane="5" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6077" points="761" swimtime="00:00:24.13" resultid="11364" heatid="11418" lane="4" entrytime="00:00:23.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Szydło" birthdate="1992-01-01" gender="F" nation="POL" swrid="4072250" athleteid="9811" />
            <ATHLETE firstname="Paweł" lastname="Korzeniowski" birthdate="1985-10-10" gender="M" nation="POL" swrid="4042751" athleteid="9797">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6077" points="918" reactiontime="+71" swimtime="00:00:22.66" resultid="9798" heatid="11419" lane="5" entrytime="00:00:22.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6238" points="850" reactiontime="+69" swimtime="00:00:25.84" resultid="9799" heatid="11450" lane="6" entrytime="00:00:26.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek., Czas lepszy od Rekordu Świata danej kat. wiek." eventid="6340" points="1109" swimtime="00:00:54.86" resultid="9800" heatid="11497" lane="4" entrytime="00:00:54.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6467" points="932" reactiontime="+70" swimtime="00:00:24.19" resultid="9801" heatid="11542" lane="5" entrytime="00:00:23.12" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9802" heatid="11597" lane="4" entrytime="00:00:52.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Budzis" birthdate="1990-01-01" gender="F" nation="POL" swrid="4060627" athleteid="9809">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6220" points="843" reactiontime="+70" swimtime="00:00:31.57" resultid="9810" heatid="11441" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-01-01" gender="M" nation="POL" athleteid="9745">
              <RESULTS>
                <RESULT eventid="6077" points="531" reactiontime="+73" swimtime="00:00:28.20" resultid="9746" heatid="11412" lane="6" entrytime="00:00:28.70" />
                <RESULT eventid="6306" points="466" reactiontime="+76" swimtime="00:01:02.63" resultid="9748" heatid="11475" lane="1" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="578" reactiontime="+74" swimtime="00:02:13.42" resultid="9749" heatid="11569" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:04.02" />
                    <SPLIT distance="150" swimtime="00:01:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9750" heatid="11592" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="6738" points="669" reactiontime="+73" swimtime="00:04:36.90" resultid="9751" heatid="11636" lane="4" entrytime="00:04:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:40.81" />
                    <SPLIT distance="200" swimtime="00:02:15.85" />
                    <SPLIT distance="250" swimtime="00:02:51.12" />
                    <SPLIT distance="300" swimtime="00:03:26.57" />
                    <SPLIT distance="350" swimtime="00:04:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" points="691" reactiontime="+79" swimtime="00:09:38.07" resultid="9823" heatid="11645" lane="7" entrytime="00:09:59.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:41.98" />
                    <SPLIT distance="200" swimtime="00:02:18.13" />
                    <SPLIT distance="250" swimtime="00:02:54.52" />
                    <SPLIT distance="300" swimtime="00:03:31.16" />
                    <SPLIT distance="350" swimtime="00:04:07.60" />
                    <SPLIT distance="400" swimtime="00:04:44.25" />
                    <SPLIT distance="450" swimtime="00:05:20.83" />
                    <SPLIT distance="500" swimtime="00:05:57.69" />
                    <SPLIT distance="550" swimtime="00:06:34.08" />
                    <SPLIT distance="600" swimtime="00:07:10.93" />
                    <SPLIT distance="650" swimtime="00:07:47.79" />
                    <SPLIT distance="700" swimtime="00:08:24.67" />
                    <SPLIT distance="750" swimtime="00:09:01.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Pilarska" birthdate="1997-01-01" gender="F" nation="POL" swrid="4282150" athleteid="9767">
              <RESULTS>
                <RESULT eventid="6059" points="783" reactiontime="+72" swimtime="00:00:27.43" resultid="9768" heatid="11401" lane="0" entrytime="00:00:28.30" />
                <RESULT eventid="6450" points="831" reactiontime="+73" swimtime="00:00:29.34" resultid="9769" heatid="11528" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Rybinski" birthdate="1993-10-11" gender="M" nation="POL" swrid="4087262" athleteid="9774">
              <RESULTS>
                <RESULT eventid="6077" points="814" swimtime="00:00:24.46" resultid="9775" heatid="11419" lane="1" entrytime="00:00:23.50" />
                <RESULT eventid="6306" points="715" reactiontime="+61" swimtime="00:00:54.31" resultid="9776" heatid="11479" lane="6" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="9777" heatid="11542" lane="2" entrytime="00:00:24.50" />
                <RESULT eventid="6535" points="793" reactiontime="+65" swimtime="00:02:00.08" resultid="9778" heatid="11571" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="100" swimtime="00:00:58.18" />
                    <SPLIT distance="150" swimtime="00:01:29.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="785" reactiontime="+63" swimtime="00:00:58.44" resultid="9779" heatid="11597" lane="8" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6610" reactiontime="+67" swimtime="00:01:32.20" resultid="11371" heatid="11582" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.64" />
                    <SPLIT distance="100" swimtime="00:00:44.89" />
                    <SPLIT distance="150" swimtime="00:01:08.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9780" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="9797" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="9770" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9774" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6779" reactiontime="+77" swimtime="00:01:43.30" resultid="11375" heatid="12332" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                    <SPLIT distance="100" swimtime="00:00:54.73" />
                    <SPLIT distance="150" swimtime="00:01:20.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9797" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="9780" number="2" reactiontime="+194" />
                    <RELAYPOSITION athleteid="9774" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="9770" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+90" swimtime="00:01:59.59" resultid="11372" heatid="11582" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="150" swimtime="00:01:31.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9794" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="9752" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="9759" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="9745" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G3" eventid="6779" reactiontime="+81" status="DSQ" swimtime="00:00:00.00" resultid="11376" heatid="12332" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:44.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9759" number="1" reactiontime="+81" status="DSQ" />
                    <RELAYPOSITION athleteid="9752" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="9739" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="9745" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+79" swimtime="00:01:55.38" resultid="11370" heatid="11580" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="100" swimtime="00:00:56.86" />
                    <SPLIT distance="150" swimtime="00:01:28.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9809" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="9812" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="9811" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="9767" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" reactiontime="+76" swimtime="00:02:09.13" resultid="11374" heatid="11639" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:40.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9809" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="9811" number="2" />
                    <RELAYPOSITION athleteid="9767" number="3" />
                    <RELAYPOSITION athleteid="9812" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+74" swimtime="00:01:53.42" resultid="9816" heatid="11435" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.49" />
                    <SPLIT distance="100" swimtime="00:00:44.95" />
                    <SPLIT distance="150" swimtime="00:01:25.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9797" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="9780" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="9785" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="9767" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6391" reactiontime="+75" swimtime="00:01:53.31" resultid="9818" heatid="11506" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="100" swimtime="00:00:55.07" />
                    <SPLIT distance="150" swimtime="00:01:24.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9797" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9780" number="2" />
                    <RELAYPOSITION athleteid="9767" number="3" />
                    <RELAYPOSITION athleteid="9812" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+75" swimtime="00:02:10.42" resultid="11366" heatid="11505" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="150" swimtime="00:01:29.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9809" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9774" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="9770" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="9785" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8492" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Zuzanna" lastname="Janecka" birthdate="1999-01-01" gender="F" nation="POL" swrid="4853973" athleteid="8491">
              <RESULTS>
                <RESULT eventid="6220" points="527" reactiontime="+88" swimtime="00:00:35.90" resultid="8493" heatid="11440" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="6289" points="678" swimtime="00:01:05.80" resultid="8494" heatid="11465" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="611" reactiontime="+77" swimtime="00:02:25.12" resultid="8495" heatid="11559" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="477" reactiontime="+100" swimtime="00:02:48.60" resultid="8496" heatid="11600" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="576" reactiontime="+74" swimtime="00:05:08.52" resultid="8497" heatid="11628" lane="6" entrytime="00:05:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:50.64" />
                    <SPLIT distance="200" swimtime="00:02:29.47" />
                    <SPLIT distance="250" swimtime="00:03:09.18" />
                    <SPLIT distance="300" swimtime="00:03:49.13" />
                    <SPLIT distance="350" swimtime="00:04:29.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11390" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="1978-01-01" gender="M" nation="POL" athleteid="11389">
              <RESULTS>
                <RESULT eventid="6077" points="500" swimtime="00:00:29.23" resultid="11391" heatid="11410" lane="4" entrytime="00:00:30.68" />
                <RESULT eventid="6306" points="460" reactiontime="+83" swimtime="00:01:06.40" resultid="11392" heatid="11473" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7142" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Wiatrowski" birthdate="1996-01-01" gender="M" nation="POL" swrid="4290292" athleteid="7141">
              <RESULTS>
                <RESULT eventid="6077" points="599" reactiontime="+83" swimtime="00:00:27.09" resultid="7143" heatid="11413" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="6111" points="514" swimtime="00:02:30.43" resultid="7144" heatid="11427" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:08.66" />
                    <SPLIT distance="150" swimtime="00:01:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="430" reactiontime="+80" swimtime="00:00:33.18" resultid="7145" heatid="11448" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="6340" points="545" reactiontime="+74" swimtime="00:01:07.56" resultid="7146" heatid="11494" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="538" reactiontime="+71" swimtime="00:00:29.13" resultid="7147" heatid="11537" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="6704" points="569" reactiontime="+68" swimtime="00:00:34.09" resultid="7148" heatid="11619" lane="0" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8681" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Juruć" birthdate="1996-01-01" gender="M" nation="POL" swrid="4195546" athleteid="8680">
              <RESULTS>
                <RESULT eventid="6203" points="630" reactiontime="+70" swimtime="00:18:49.41" resultid="8682" heatid="11652" lane="3" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:04.29" />
                    <SPLIT distance="150" swimtime="00:01:40.12" />
                    <SPLIT distance="200" swimtime="00:02:16.45" />
                    <SPLIT distance="250" swimtime="00:02:53.74" />
                    <SPLIT distance="300" swimtime="00:03:30.78" />
                    <SPLIT distance="350" swimtime="00:04:08.25" />
                    <SPLIT distance="400" swimtime="00:04:45.79" />
                    <SPLIT distance="450" swimtime="00:05:23.39" />
                    <SPLIT distance="500" swimtime="00:06:01.03" />
                    <SPLIT distance="550" swimtime="00:06:38.48" />
                    <SPLIT distance="600" swimtime="00:07:16.04" />
                    <SPLIT distance="650" swimtime="00:07:53.47" />
                    <SPLIT distance="700" swimtime="00:08:30.81" />
                    <SPLIT distance="750" swimtime="00:09:08.81" />
                    <SPLIT distance="800" swimtime="00:09:46.79" />
                    <SPLIT distance="850" swimtime="00:10:25.84" />
                    <SPLIT distance="900" swimtime="00:11:05.01" />
                    <SPLIT distance="950" swimtime="00:11:44.24" />
                    <SPLIT distance="1000" swimtime="00:12:22.60" />
                    <SPLIT distance="1050" swimtime="00:13:01.49" />
                    <SPLIT distance="1100" swimtime="00:13:40.78" />
                    <SPLIT distance="1150" swimtime="00:14:20.06" />
                    <SPLIT distance="1200" swimtime="00:14:59.03" />
                    <SPLIT distance="1250" swimtime="00:15:37.70" />
                    <SPLIT distance="1300" swimtime="00:16:16.85" />
                    <SPLIT distance="1350" swimtime="00:16:56.05" />
                    <SPLIT distance="1400" swimtime="00:17:34.35" />
                    <SPLIT distance="1450" swimtime="00:18:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="8683" heatid="11477" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8684" heatid="11606" lane="0" entrytime="00:02:30.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8685" heatid="11637" lane="3" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" clubid="8692" name="UKS Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Tadeusz" lastname="Gołembiewski" birthdate="1985-03-14" gender="M" nation="POL" license="503415700164" swrid="4061025" athleteid="9513">
              <RESULTS>
                <RESULT eventid="6467" points="497" reactiontime="+82" swimtime="00:00:29.82" resultid="9514" heatid="11539" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="6535" points="576" reactiontime="+90" swimtime="00:02:13.95" resultid="9515" heatid="11570" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9516" heatid="11595" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9517" heatid="11637" lane="6" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Rybak-Starczak" birthdate="1975-01-16" gender="F" nation="POL" license="503415600144" swrid="5439532" athleteid="9495">
              <RESULTS>
                <RESULT eventid="6094" points="516" reactiontime="+100" swimtime="00:03:07.02" resultid="9496" heatid="11422" lane="5" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:31.56" />
                    <SPLIT distance="150" swimtime="00:02:23.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="605" reactiontime="+99" swimtime="00:03:20.03" resultid="9497" heatid="11454" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:36.36" />
                    <SPLIT distance="150" swimtime="00:02:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="526" reactiontime="+121" swimtime="00:01:25.63" resultid="9498" heatid="11484" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="578" swimtime="00:01:33.05" resultid="9499" heatid="11511" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Jaruga" birthdate="1974-08-05" gender="F" nation="POL" athleteid="8693">
              <RESULTS>
                <RESULT eventid="6186" points="537" swimtime="00:23:52.67" resultid="8694" heatid="11650" lane="0" entrytime="00:26:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:27.77" />
                    <SPLIT distance="150" swimtime="00:02:14.86" />
                    <SPLIT distance="200" swimtime="00:03:02.30" />
                    <SPLIT distance="250" swimtime="00:03:50.04" />
                    <SPLIT distance="300" swimtime="00:04:38.50" />
                    <SPLIT distance="350" swimtime="00:05:26.80" />
                    <SPLIT distance="400" swimtime="00:06:15.28" />
                    <SPLIT distance="450" swimtime="00:07:03.57" />
                    <SPLIT distance="500" swimtime="00:07:52.07" />
                    <SPLIT distance="550" swimtime="00:08:40.55" />
                    <SPLIT distance="600" swimtime="00:09:29.09" />
                    <SPLIT distance="650" swimtime="00:10:17.74" />
                    <SPLIT distance="700" swimtime="00:11:06.15" />
                    <SPLIT distance="750" swimtime="00:11:54.60" />
                    <SPLIT distance="800" swimtime="00:12:42.92" />
                    <SPLIT distance="850" swimtime="00:13:31.44" />
                    <SPLIT distance="900" swimtime="00:14:19.55" />
                    <SPLIT distance="950" swimtime="00:15:07.57" />
                    <SPLIT distance="1000" swimtime="00:15:55.73" />
                    <SPLIT distance="1050" swimtime="00:16:43.91" />
                    <SPLIT distance="1100" swimtime="00:17:32.41" />
                    <SPLIT distance="1150" swimtime="00:18:20.62" />
                    <SPLIT distance="1200" swimtime="00:19:08.64" />
                    <SPLIT distance="1250" swimtime="00:19:56.41" />
                    <SPLIT distance="1300" swimtime="00:20:43.89" />
                    <SPLIT distance="1350" swimtime="00:21:31.80" />
                    <SPLIT distance="1400" swimtime="00:22:19.45" />
                    <SPLIT distance="1450" swimtime="00:23:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="418" reactiontime="+85" swimtime="00:02:54.45" resultid="8695" heatid="11556" lane="5" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:08.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="407" reactiontime="+97" swimtime="00:07:16.26" resultid="8696" heatid="11573" lane="2" entrytime="00:08:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:51.91" />
                    <SPLIT distance="150" swimtime="00:02:50.25" />
                    <SPLIT distance="200" swimtime="00:03:46.55" />
                    <SPLIT distance="250" swimtime="00:04:44.66" />
                    <SPLIT distance="300" swimtime="00:05:44.19" />
                    <SPLIT distance="350" swimtime="00:06:32.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" license="503415700180" swrid="4754708" athleteid="9500">
              <RESULTS>
                <RESULT eventid="6203" points="560" reactiontime="+69" swimtime="00:28:00.25" resultid="9501" heatid="11653" lane="9" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.65" />
                    <SPLIT distance="100" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:45.15" />
                    <SPLIT distance="200" swimtime="00:03:40.81" />
                    <SPLIT distance="250" swimtime="00:04:36.48" />
                    <SPLIT distance="300" swimtime="00:05:31.99" />
                    <SPLIT distance="350" swimtime="00:06:28.52" />
                    <SPLIT distance="400" swimtime="00:07:23.74" />
                    <SPLIT distance="450" swimtime="00:08:20.11" />
                    <SPLIT distance="500" swimtime="00:09:16.09" />
                    <SPLIT distance="550" swimtime="00:10:12.16" />
                    <SPLIT distance="600" swimtime="00:11:08.81" />
                    <SPLIT distance="650" swimtime="00:12:04.94" />
                    <SPLIT distance="700" swimtime="00:13:00.76" />
                    <SPLIT distance="750" swimtime="00:13:56.92" />
                    <SPLIT distance="800" swimtime="00:14:53.16" />
                    <SPLIT distance="850" swimtime="00:15:49.25" />
                    <SPLIT distance="900" swimtime="00:16:45.96" />
                    <SPLIT distance="950" swimtime="00:17:42.36" />
                    <SPLIT distance="1000" swimtime="00:18:38.54" />
                    <SPLIT distance="1050" swimtime="00:19:35.64" />
                    <SPLIT distance="1100" swimtime="00:20:31.73" />
                    <SPLIT distance="1150" swimtime="00:21:28.34" />
                    <SPLIT distance="1200" swimtime="00:22:25.47" />
                    <SPLIT distance="1250" swimtime="00:23:21.86" />
                    <SPLIT distance="1300" swimtime="00:24:18.76" />
                    <SPLIT distance="1350" swimtime="00:25:14.72" />
                    <SPLIT distance="1400" swimtime="00:26:10.47" />
                    <SPLIT distance="1450" swimtime="00:27:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="376" reactiontime="+90" swimtime="00:00:48.04" resultid="9502" heatid="11445" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="6501" points="331" reactiontime="+91" swimtime="00:01:48.49" resultid="9503" heatid="11549" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="489" reactiontime="+105" swimtime="00:03:50.88" resultid="9504" heatid="11602" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                    <SPLIT distance="100" swimtime="00:01:55.69" />
                    <SPLIT distance="150" swimtime="00:02:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="9505" heatid="11631" lane="8" entrytime="00:07:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska-Błachowicz" birthdate="1954-07-13" gender="F" nation="POL" license="503415600184" swrid="5471727" athleteid="9506">
              <RESULTS>
                <RESULT eventid="6220" points="314" reactiontime="+96" swimtime="00:00:58.85" resultid="9507" heatid="11439" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="6323" points="253" reactiontime="+100" swimtime="00:02:09.37" resultid="9508" heatid="11482" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="188" swimtime="00:01:01.75" resultid="9509" heatid="11524" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="6484" points="271" reactiontime="+99" swimtime="00:02:15.23" resultid="9510" heatid="11544" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M3 - Pływak obrócił się na plecy w czasie wyścigu (z wyjątkiem wykonywania nawrotu, po dotknięciu dłońmi, a przed opuszczeniem ściany)." eventid="6618" reactiontime="+107" status="DSQ" swimtime="00:00:00.00" resultid="9511" heatid="11586" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="303" reactiontime="+105" swimtime="00:00:57.89" resultid="9512" heatid="11609" lane="2" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Miśkiewicz" birthdate="1959-03-24" gender="M" nation="POL" license="503415700185" swrid="4920302" athleteid="9489">
              <RESULTS>
                <RESULT eventid="6077" points="267" reactiontime="+115" swimtime="00:00:41.64" resultid="9490" heatid="11405" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="6238" points="292" reactiontime="+97" swimtime="00:00:47.34" resultid="9491" heatid="11445" lane="0" entrytime="00:00:47.00" />
                <RESULT eventid="6340" points="243" swimtime="00:01:49.39" resultid="9492" heatid="11489" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="274" reactiontime="+91" swimtime="00:01:43.98" resultid="9493" heatid="11550" lane="0" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="322" reactiontime="+103" swimtime="00:03:49.06" resultid="9494" heatid="11603" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                    <SPLIT distance="100" swimtime="00:01:54.15" />
                    <SPLIT distance="150" swimtime="00:02:53.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" swimtime="00:02:52.58" resultid="9518" heatid="11435" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                    <SPLIT distance="100" swimtime="00:01:34.72" />
                    <SPLIT distance="150" swimtime="00:02:11.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9489" number="1" />
                    <RELAYPOSITION athleteid="9506" number="2" />
                    <RELAYPOSITION athleteid="9495" number="3" />
                    <RELAYPOSITION athleteid="9500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+99" swimtime="00:03:04.85" resultid="9519" heatid="11505" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:44.54" />
                    <SPLIT distance="150" swimtime="00:02:39.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9489" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="9506" number="2" />
                    <RELAYPOSITION athleteid="9495" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="9500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8121" name="Delfin Masters Łódź" />
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="9548" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Monika" lastname="Dargas-Miszczak" birthdate="1981-09-06" gender="F" nation="POL" license="504214600090" swrid="5486407" athleteid="9555">
              <RESULTS>
                <RESULT eventid="6059" points="492" reactiontime="+84" swimtime="00:00:33.28" resultid="9556" heatid="11394" lane="3" />
                <RESULT eventid="6289" points="499" reactiontime="+80" swimtime="00:01:13.72" resultid="9557" heatid="11461" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="536" reactiontime="+67" swimtime="00:00:36.07" resultid="9558" heatid="11523" lane="6" />
                <RESULT eventid="6518" points="516" swimtime="00:02:41.20" resultid="9559" heatid="11554" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:16.49" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="389" swimtime="00:01:28.45" resultid="9560" heatid="11585" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="504" swimtime="00:05:47.97" resultid="9561" heatid="11624" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:02:04.36" />
                    <SPLIT distance="200" swimtime="00:02:49.84" />
                    <SPLIT distance="250" swimtime="00:03:35.15" />
                    <SPLIT distance="300" swimtime="00:04:20.93" />
                    <SPLIT distance="350" swimtime="00:05:05.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Sutowski" birthdate="1959-12-03" gender="M" nation="POL" license="104214700079" swrid="4992657" athleteid="9610">
              <RESULTS>
                <RESULT eventid="6077" points="253" reactiontime="+100" swimtime="00:00:42.39" resultid="9611" heatid="11405" lane="0" entrytime="00:00:43.15" entrycourse="SCM" />
                <RESULT eventid="6169" points="428" reactiontime="+105" swimtime="00:13:41.98" resultid="9612" heatid="11649" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:37.01" />
                    <SPLIT distance="150" swimtime="00:02:29.55" />
                    <SPLIT distance="200" swimtime="00:03:21.75" />
                    <SPLIT distance="250" swimtime="00:04:14.69" />
                    <SPLIT distance="300" swimtime="00:05:08.13" />
                    <SPLIT distance="350" swimtime="00:06:00.31" />
                    <SPLIT distance="400" swimtime="00:06:51.82" />
                    <SPLIT distance="450" swimtime="00:07:44.14" />
                    <SPLIT distance="500" swimtime="00:08:35.55" />
                    <SPLIT distance="550" swimtime="00:09:26.81" />
                    <SPLIT distance="600" swimtime="00:10:18.01" />
                    <SPLIT distance="650" swimtime="00:11:10.76" />
                    <SPLIT distance="700" swimtime="00:12:02.93" />
                    <SPLIT distance="750" swimtime="00:12:54.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="350" reactiontime="+104" swimtime="00:01:24.89" resultid="9613" heatid="11469" lane="8" entrytime="00:01:28.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="181" reactiontime="+100" swimtime="00:00:51.52" resultid="9614" heatid="11530" lane="0" />
                <RESULT eventid="6535" points="390" reactiontime="+106" swimtime="00:03:06.75" resultid="9615" heatid="11562" lane="3" entrytime="00:06:49.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                    <SPLIT distance="150" swimtime="00:02:21.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" license="104214700039" swrid="5552366" athleteid="9597">
              <RESULTS>
                <RESULT eventid="6077" points="465" reactiontime="+89" swimtime="00:00:30.80" resultid="9598" heatid="11403" lane="2" />
                <RESULT eventid="6169" points="449" reactiontime="+92" swimtime="00:11:18.72" resultid="9599" heatid="11649" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:56.86" />
                    <SPLIT distance="200" swimtime="00:02:38.21" />
                    <SPLIT distance="250" swimtime="00:03:20.46" />
                    <SPLIT distance="300" swimtime="00:04:03.56" />
                    <SPLIT distance="350" swimtime="00:04:47.08" />
                    <SPLIT distance="400" swimtime="00:05:31.27" />
                    <SPLIT distance="450" swimtime="00:06:15.03" />
                    <SPLIT distance="500" swimtime="00:06:58.80" />
                    <SPLIT distance="550" swimtime="00:07:42.65" />
                    <SPLIT distance="600" swimtime="00:08:26.20" />
                    <SPLIT distance="650" swimtime="00:09:09.37" />
                    <SPLIT distance="700" swimtime="00:09:52.75" />
                    <SPLIT distance="750" swimtime="00:10:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="460" reactiontime="+87" swimtime="00:01:17.69" resultid="9600" heatid="11492" lane="8" entrytime="00:01:18.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="623" reactiontime="+88" swimtime="00:01:17.33" resultid="9601" heatid="11514" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="479" reactiontime="+92" swimtime="00:02:26.59" resultid="9602" heatid="11562" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="462" reactiontime="+91" swimtime="00:05:17.99" resultid="9603" heatid="11635" lane="8" entrytime="00:05:19.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:13.41" />
                    <SPLIT distance="150" swimtime="00:01:53.27" />
                    <SPLIT distance="200" swimtime="00:02:34.34" />
                    <SPLIT distance="250" swimtime="00:03:16.16" />
                    <SPLIT distance="300" swimtime="00:03:57.05" />
                    <SPLIT distance="350" swimtime="00:04:38.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Nowak" birthdate="1952-12-17" gender="M" nation="POL" license="504214700029" swrid="4302652" athleteid="9660">
              <RESULTS>
                <RESULT eventid="6111" points="655" reactiontime="+90" swimtime="00:03:24.61" resultid="9661" heatid="11427" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:43.88" />
                    <SPLIT distance="150" swimtime="00:02:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="763" reactiontime="+86" swimtime="00:03:22.72" resultid="9662" heatid="11455" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:35.29" />
                    <SPLIT distance="150" swimtime="00:02:28.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="783" reactiontime="+89" swimtime="00:01:24.16" resultid="9663" heatid="11487" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="804" reactiontime="+89" swimtime="00:01:28.65" resultid="9664" heatid="11514" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="674" reactiontime="+93" swimtime="00:07:31.85" resultid="9665" heatid="11576" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                    <SPLIT distance="100" swimtime="00:01:50.40" />
                    <SPLIT distance="150" swimtime="00:03:51.64" />
                    <SPLIT distance="200" swimtime="00:04:49.97" />
                    <SPLIT distance="250" swimtime="00:05:48.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="811" reactiontime="+83" swimtime="00:00:38.10" resultid="9666" heatid="11614" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" license="504214700003" swrid="4270348" athleteid="9654">
              <RESULTS>
                <RESULT eventid="6111" points="624" reactiontime="+87" swimtime="00:02:34.90" resultid="9655" heatid="11426" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:01:59.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="501" reactiontime="+103" swimtime="00:20:44.61" resultid="9656" heatid="11654" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                    <SPLIT distance="200" swimtime="00:02:41.19" />
                    <SPLIT distance="250" swimtime="00:03:22.92" />
                    <SPLIT distance="300" swimtime="00:04:04.49" />
                    <SPLIT distance="350" swimtime="00:04:46.16" />
                    <SPLIT distance="400" swimtime="00:05:27.91" />
                    <SPLIT distance="450" swimtime="00:06:09.37" />
                    <SPLIT distance="500" swimtime="00:06:50.85" />
                    <SPLIT distance="550" swimtime="00:07:32.31" />
                    <SPLIT distance="600" swimtime="00:08:14.29" />
                    <SPLIT distance="650" swimtime="00:08:56.51" />
                    <SPLIT distance="700" swimtime="00:09:38.75" />
                    <SPLIT distance="750" swimtime="00:10:20.79" />
                    <SPLIT distance="800" swimtime="00:11:02.91" />
                    <SPLIT distance="850" swimtime="00:11:45.30" />
                    <SPLIT distance="900" swimtime="00:12:27.56" />
                    <SPLIT distance="950" swimtime="00:13:09.71" />
                    <SPLIT distance="1000" swimtime="00:13:52.01" />
                    <SPLIT distance="1050" swimtime="00:14:34.51" />
                    <SPLIT distance="1100" swimtime="00:15:16.85" />
                    <SPLIT distance="1150" swimtime="00:15:58.99" />
                    <SPLIT distance="1200" swimtime="00:16:41.40" />
                    <SPLIT distance="1250" swimtime="00:17:23.70" />
                    <SPLIT distance="1300" swimtime="00:18:05.53" />
                    <SPLIT distance="1350" swimtime="00:18:46.98" />
                    <SPLIT distance="1400" swimtime="00:19:27.94" />
                    <SPLIT distance="1450" swimtime="00:20:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="670" reactiontime="+88" swimtime="00:02:48.72" resultid="9657" heatid="11459" lane="6" entrytime="00:02:50.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:05.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="9658" heatid="11519" lane="2" entrytime="00:01:18.83" entrycourse="SCM" />
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="9659" heatid="11575" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kozak" birthdate="1986-02-13" gender="M" nation="POL" license="504214700012" swrid="4992669" athleteid="9592">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="9593" heatid="11402" lane="1" />
                <RESULT eventid="6272" points="630" reactiontime="+91" swimtime="00:02:43.98" resultid="9594" heatid="11455" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:02:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="697" reactiontime="+81" swimtime="00:01:11.60" resultid="9595" heatid="11514" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="727" reactiontime="+81" swimtime="00:00:32.09" resultid="9596" heatid="11615" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" license="504214600017" swrid="4302692" athleteid="9562">
              <RESULTS>
                <RESULT eventid="6059" points="192" swimtime="00:00:57.71" resultid="9563" heatid="11394" lane="8" />
                <RESULT eventid="6145" points="373" swimtime="00:18:08.02" resultid="9564" heatid="11644" lane="8" entrytime="00:18:26.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.30" />
                    <SPLIT distance="150" swimtime="00:03:25.17" />
                    <SPLIT distance="200" swimtime="00:04:34.62" />
                    <SPLIT distance="250" swimtime="00:05:43.73" />
                    <SPLIT distance="300" swimtime="00:06:53.05" />
                    <SPLIT distance="350" swimtime="00:08:00.95" />
                    <SPLIT distance="400" swimtime="00:10:15.47" />
                    <SPLIT distance="450" swimtime="00:11:23.49" />
                    <SPLIT distance="500" swimtime="00:12:31.93" />
                    <SPLIT distance="550" swimtime="00:13:39.86" />
                    <SPLIT distance="600" swimtime="00:14:47.31" />
                    <SPLIT distance="650" swimtime="00:15:56.04" />
                    <SPLIT distance="700" swimtime="00:17:04.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="223" swimtime="00:02:03.02" resultid="9565" heatid="11462" lane="7" entrytime="00:03:40.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="356" swimtime="00:08:55.58" resultid="9566" heatid="11625" lane="1" entrytime="00:08:42.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.22" />
                    <SPLIT distance="100" swimtime="00:02:12.62" />
                    <SPLIT distance="150" swimtime="00:03:21.62" />
                    <SPLIT distance="200" swimtime="00:04:30.06" />
                    <SPLIT distance="250" swimtime="00:05:37.75" />
                    <SPLIT distance="300" swimtime="00:06:44.41" />
                    <SPLIT distance="350" swimtime="00:07:51.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Bielecka" birthdate="1988-04-07" gender="F" nation="POL" license="504214600154" athleteid="9647">
              <RESULTS>
                <RESULT eventid="6094" points="641" reactiontime="+62" swimtime="00:02:45.74" resultid="9648" heatid="11420" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="543" reactiontime="+80" swimtime="00:22:30.77" resultid="9649" heatid="11651" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:23.69" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                    <SPLIT distance="200" swimtime="00:02:54.10" />
                    <SPLIT distance="250" swimtime="00:03:39.08" />
                    <SPLIT distance="300" swimtime="00:04:24.70" />
                    <SPLIT distance="350" swimtime="00:05:09.54" />
                    <SPLIT distance="400" swimtime="00:05:54.84" />
                    <SPLIT distance="450" swimtime="00:06:40.28" />
                    <SPLIT distance="500" swimtime="00:07:26.26" />
                    <SPLIT distance="550" swimtime="00:08:11.53" />
                    <SPLIT distance="600" swimtime="00:08:57.20" />
                    <SPLIT distance="650" swimtime="00:09:42.61" />
                    <SPLIT distance="700" swimtime="00:10:28.37" />
                    <SPLIT distance="750" swimtime="00:11:14.07" />
                    <SPLIT distance="800" swimtime="00:11:59.33" />
                    <SPLIT distance="850" swimtime="00:12:44.81" />
                    <SPLIT distance="900" swimtime="00:13:29.74" />
                    <SPLIT distance="950" swimtime="00:14:14.89" />
                    <SPLIT distance="1000" swimtime="00:15:00.05" />
                    <SPLIT distance="1050" swimtime="00:15:45.35" />
                    <SPLIT distance="1100" swimtime="00:16:30.37" />
                    <SPLIT distance="1150" swimtime="00:17:15.21" />
                    <SPLIT distance="1200" swimtime="00:18:01.59" />
                    <SPLIT distance="1250" swimtime="00:18:46.96" />
                    <SPLIT distance="1300" swimtime="00:19:32.24" />
                    <SPLIT distance="1350" swimtime="00:20:17.54" />
                    <SPLIT distance="1400" swimtime="00:21:03.02" />
                    <SPLIT distance="1450" swimtime="00:21:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="489" swimtime="00:03:01.17" resultid="9650" heatid="11498" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="600" reactiontime="+72" swimtime="00:00:33.41" resultid="9651" heatid="11523" lane="5" />
                <RESULT eventid="6552" status="DNS" swimtime="00:00:00.00" resultid="9652" heatid="11572" lane="3" />
                <RESULT eventid="6618" points="514" reactiontime="+69" swimtime="00:01:18.13" resultid="9653" heatid="11585" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kośla" birthdate="1993-01-05" gender="F" nation="POL" license="104214600085" swrid="4086961" athleteid="9579">
              <RESULTS>
                <RESULT eventid="6059" points="644" reactiontime="+79" swimtime="00:00:29.28" resultid="9580" heatid="11393" lane="5" />
                <RESULT eventid="6220" points="750" reactiontime="+72" swimtime="00:00:32.50" resultid="9581" heatid="11438" lane="3" />
                <RESULT eventid="6289" status="DNS" swimtime="00:00:00.00" resultid="9582" heatid="11462" lane="0" />
                <RESULT eventid="6484" points="756" reactiontime="+72" swimtime="00:01:09.99" resultid="9583" heatid="11544" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Sobczak-Porada" birthdate="1987-07-20" gender="F" nation="POL" license="504214600056" athleteid="9567">
              <RESULTS>
                <RESULT eventid="6059" points="206" reactiontime="+96" swimtime="00:00:44.30" resultid="9568" heatid="11394" lane="2" />
                <RESULT eventid="6289" points="179" reactiontime="+99" swimtime="00:01:42.53" resultid="9569" heatid="11461" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" status="DNS" swimtime="00:00:00.00" resultid="9570" heatid="11555" lane="3" />
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="9571" heatid="11608" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szymański" birthdate="1980-10-04" gender="M" nation="POL" license="504214700028" swrid="4542528" athleteid="9584">
              <RESULTS>
                <RESULT eventid="6077" points="891" swimtime="00:00:24.12" resultid="9585" heatid="11417" lane="4" entrytime="00:00:24.88" entrycourse="SCM" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="9586" heatid="11426" lane="9" />
                <RESULT eventid="6238" points="944" reactiontime="+75" swimtime="00:00:27.67" resultid="9587" heatid="11450" lane="9" entrytime="00:00:27.92" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6340" points="944" reactiontime="+68" swimtime="00:01:00.98" resultid="9588" heatid="11497" lane="0" entrytime="00:01:01.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="848" swimtime="00:00:26.54" resultid="9589" heatid="11529" lane="4" />
                <RESULT eventid="6501" points="949" reactiontime="+71" swimtime="00:01:00.08" resultid="9590" heatid="11553" lane="1" entrytime="00:01:04.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="801" reactiontime="+76" swimtime="00:00:31.31" resultid="9591" heatid="11614" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" license="104214700058" swrid="5506638" athleteid="9616">
              <RESULTS>
                <RESULT eventid="6077" points="531" reactiontime="+70" swimtime="00:00:27.19" resultid="9617" heatid="11404" lane="0" />
                <RESULT eventid="6111" points="610" reactiontime="+84" swimtime="00:02:30.11" resultid="9618" heatid="11426" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="673" reactiontime="+75" swimtime="00:02:40.40" resultid="9619" heatid="11460" lane="8" entrytime="00:02:38.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="9620" heatid="11487" lane="5" />
                <RESULT eventid="6433" points="621" reactiontime="+76" swimtime="00:01:14.42" resultid="9621" heatid="11513" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="535" reactiontime="+77" swimtime="00:02:17.25" resultid="9622" heatid="11561" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9623" heatid="11589" lane="7" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="9624" heatid="11615" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymański" birthdate="1981-11-04" gender="M" nation="POL" license="504214700060" swrid="4542568" athleteid="9625">
              <RESULTS>
                <RESULT eventid="6077" points="600" reactiontime="+82" swimtime="00:00:27.51" resultid="9626" heatid="11403" lane="3" />
                <RESULT eventid="6238" points="573" reactiontime="+93" swimtime="00:00:32.68" resultid="9627" heatid="11443" lane="7" />
                <RESULT eventid="6340" points="543" reactiontime="+91" swimtime="00:01:13.30" resultid="9628" heatid="11488" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="607" swimtime="00:00:29.67" resultid="9629" heatid="11530" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Petryszyn" birthdate="1994-07-31" gender="F" nation="POL" license="104214600156" swrid="4369524" athleteid="9572">
              <RESULTS>
                <RESULT eventid="6059" points="719" reactiontime="+73" swimtime="00:00:28.22" resultid="9573" heatid="11394" lane="7" />
                <RESULT eventid="6220" points="758" reactiontime="+84" swimtime="00:00:32.39" resultid="9574" heatid="11438" lane="2" />
                <RESULT eventid="6289" points="713" reactiontime="+74" swimtime="00:01:02.81" resultid="9575" heatid="11461" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="750" reactiontime="+76" swimtime="00:00:30.36" resultid="9576" heatid="11524" lane="9" />
                <RESULT eventid="6484" points="724" reactiontime="+80" swimtime="00:01:10.99" resultid="9577" heatid="11543" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="616" reactiontime="+95" swimtime="00:02:40.34" resultid="9578" heatid="11598" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:17.15" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" license="504214700005" swrid="4183799" athleteid="9630">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="9631" heatid="11414" lane="9" entrytime="00:00:27.89" entrycourse="SCM" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="9632" heatid="11426" lane="2" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="9633" heatid="11475" lane="6" entrytime="00:01:02.66" entrycourse="SCM" />
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="9634" heatid="11493" lane="4" entrytime="00:01:11.11" entrycourse="SCM" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="9635" heatid="11536" lane="1" entrytime="00:00:32.17" entrycourse="SCM" />
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="9636" heatid="11575" lane="5" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="9637" heatid="11589" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Sutowski" birthdate="1993-02-18" gender="M" nation="POL" license="504214700099" swrid="4073514" athleteid="9604">
              <RESULTS>
                <RESULT eventid="6077" points="512" swimtime="00:00:28.54" resultid="9605" heatid="11412" lane="9" entrytime="00:00:29.42" entrycourse="SCM" />
                <RESULT eventid="6306" points="447" reactiontime="+79" swimtime="00:01:03.49" resultid="9606" heatid="11473" lane="8" entrytime="00:01:08.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="346" reactiontime="+84" swimtime="00:01:18.58" resultid="9607" heatid="11487" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="380" swimtime="00:00:32.72" resultid="9608" heatid="11534" lane="4" entrytime="00:00:34.49" entrycourse="SCM" />
                <RESULT eventid="6535" points="402" reactiontime="+79" swimtime="00:02:30.63" resultid="9609" heatid="11561" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:51.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" license="504214700091" swrid="5506635" athleteid="9638">
              <RESULTS>
                <RESULT eventid="6077" points="766" reactiontime="+69" swimtime="00:00:26.08" resultid="9639" heatid="11416" lane="0" entrytime="00:00:26.01" entrycourse="SCM" />
                <RESULT eventid="6169" points="522" reactiontime="+78" swimtime="00:10:45.25" resultid="9640" heatid="11649" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:02:34.25" />
                    <SPLIT distance="250" swimtime="00:03:15.02" />
                    <SPLIT distance="300" swimtime="00:03:55.59" />
                    <SPLIT distance="350" swimtime="00:04:36.19" />
                    <SPLIT distance="400" swimtime="00:05:16.98" />
                    <SPLIT distance="450" swimtime="00:05:57.86" />
                    <SPLIT distance="500" swimtime="00:06:38.72" />
                    <SPLIT distance="550" swimtime="00:07:20.00" />
                    <SPLIT distance="600" swimtime="00:08:01.74" />
                    <SPLIT distance="650" swimtime="00:08:43.81" />
                    <SPLIT distance="700" swimtime="00:09:26.32" />
                    <SPLIT distance="750" swimtime="00:10:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="588" reactiontime="+77" swimtime="00:00:33.25" resultid="9641" heatid="11443" lane="6" />
                <RESULT eventid="6306" points="716" swimtime="00:00:59.13" resultid="9642" heatid="11467" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="813" reactiontime="+77" swimtime="00:01:10.78" resultid="9643" heatid="11520" lane="7" entrytime="00:01:12.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="674" reactiontime="+71" swimtime="00:00:29.28" resultid="9644" heatid="11538" lane="6" entrytime="00:00:29.31" entrycourse="SCM" />
                <RESULT eventid="6704" points="817" reactiontime="+69" swimtime="00:00:32.39" resultid="9645" heatid="11622" lane="5" entrytime="00:00:31.89" entrycourse="SCM" />
                <RESULT eventid="6738" points="470" reactiontime="+74" swimtime="00:05:16.11" resultid="9646" heatid="11629" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="150" swimtime="00:01:50.54" />
                    <SPLIT distance="200" swimtime="00:02:31.45" />
                    <SPLIT distance="250" swimtime="00:03:13.37" />
                    <SPLIT distance="300" swimtime="00:03:55.93" />
                    <SPLIT distance="350" swimtime="00:04:35.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olga" lastname="Krysiak" birthdate="1991-06-07" gender="F" nation="POL" license="104214600021" athleteid="9549">
              <RESULTS>
                <RESULT eventid="6059" points="690" swimtime="00:00:29.30" resultid="9550" heatid="11394" lane="1" />
                <RESULT eventid="6289" points="657" reactiontime="+67" swimtime="00:01:06.08" resultid="9552" heatid="11462" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="666" reactiontime="+70" swimtime="00:02:23.88" resultid="9553" heatid="11555" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="647" reactiontime="+73" swimtime="00:05:11.48" resultid="9554" heatid="11624" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:51.16" />
                    <SPLIT distance="200" swimtime="00:02:31.90" />
                    <SPLIT distance="250" swimtime="00:03:12.77" />
                    <SPLIT distance="300" swimtime="00:03:53.44" />
                    <SPLIT distance="350" swimtime="00:04:33.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+71" swimtime="00:01:44.61" resultid="9672" heatid="11582" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.18" />
                    <SPLIT distance="100" swimtime="00:00:52.05" />
                    <SPLIT distance="150" swimtime="00:01:19.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9584" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="9592" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9625" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="9638" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+69" swimtime="00:02:05.49" resultid="9674" heatid="12331" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:39.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9584" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="9660" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="9597" number="3" reactiontime="+90" />
                    <RELAYPOSITION athleteid="9638" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6586" reactiontime="+194" swimtime="00:01:55.47" resultid="9671" heatid="11580" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:00:59.09" />
                    <SPLIT distance="150" swimtime="00:01:27.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9647" number="1" reactiontime="+194" />
                    <RELAYPOSITION athleteid="9549" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="9579" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9572" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" reactiontime="+80" swimtime="00:02:13.37" resultid="9673" heatid="11639" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:44.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9572" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="9647" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="9555" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="9549" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+70" swimtime="00:01:46.67" resultid="9667" heatid="11434" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.16" />
                    <SPLIT distance="100" swimtime="00:00:50.17" />
                    <SPLIT distance="150" swimtime="00:01:18.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9584" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="9638" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="9549" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9572" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+70" swimtime="00:01:58.42" resultid="9669" heatid="11505" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="150" swimtime="00:01:34.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9579" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="9638" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="9572" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9584" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+72" swimtime="00:01:54.81" resultid="9668" heatid="11434" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.62" />
                    <SPLIT distance="100" swimtime="00:00:56.33" />
                    <SPLIT distance="150" swimtime="00:01:26.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9616" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9579" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="9647" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="9604" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+92" swimtime="00:02:07.60" resultid="9670" heatid="11506" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:38.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9625" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="9592" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="9647" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="9549" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="7271" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrii" lastname="Lobanov" birthdate="1962-01-01" gender="M" nation="UKR" athleteid="7270">
              <RESULTS>
                <RESULT eventid="6272" points="551" swimtime="00:03:22.30" resultid="7272" heatid="11456" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="100" swimtime="00:01:37.44" />
                    <SPLIT distance="150" swimtime="00:02:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="7273" heatid="11490" lane="9" entrytime="00:01:35.00" />
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="7274" heatid="11517" lane="0" entrytime="00:01:40.00" />
                <RESULT eventid="6704" points="485" swimtime="00:00:41.65" resultid="7275" heatid="11616" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6808" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Aleksy" lastname="Wierzchoń" birthdate="1962-01-01" gender="M" nation="POL" athleteid="6807">
              <RESULTS>
                <RESULT eventid="6077" points="475" swimtime="00:00:34.38" resultid="6809" heatid="11411" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="6203" points="484" reactiontime="+103" swimtime="00:24:56.35" resultid="6810" heatid="11654" lane="4" entrytime="00:29:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                    <SPLIT distance="100" swimtime="00:01:28.18" />
                    <SPLIT distance="150" swimtime="00:02:17.49" />
                    <SPLIT distance="200" swimtime="00:03:08.18" />
                    <SPLIT distance="250" swimtime="00:03:58.57" />
                    <SPLIT distance="300" swimtime="00:04:49.07" />
                    <SPLIT distance="350" swimtime="00:05:39.40" />
                    <SPLIT distance="400" swimtime="00:06:29.59" />
                    <SPLIT distance="450" swimtime="00:07:20.53" />
                    <SPLIT distance="500" swimtime="00:08:10.78" />
                    <SPLIT distance="550" swimtime="00:09:01.12" />
                    <SPLIT distance="600" swimtime="00:09:51.66" />
                    <SPLIT distance="650" swimtime="00:10:41.58" />
                    <SPLIT distance="700" swimtime="00:11:31.79" />
                    <SPLIT distance="750" swimtime="00:12:21.84" />
                    <SPLIT distance="800" swimtime="00:13:12.76" />
                    <SPLIT distance="850" swimtime="00:14:03.49" />
                    <SPLIT distance="900" swimtime="00:14:53.11" />
                    <SPLIT distance="950" swimtime="00:15:44.29" />
                    <SPLIT distance="1000" swimtime="00:16:34.19" />
                    <SPLIT distance="1050" swimtime="00:17:24.37" />
                    <SPLIT distance="1100" swimtime="00:18:14.71" />
                    <SPLIT distance="1150" swimtime="00:19:05.20" />
                    <SPLIT distance="1200" swimtime="00:19:55.56" />
                    <SPLIT distance="1250" swimtime="00:20:46.66" />
                    <SPLIT distance="1300" swimtime="00:21:36.48" />
                    <SPLIT distance="1350" swimtime="00:22:26.76" />
                    <SPLIT distance="1400" swimtime="00:23:17.56" />
                    <SPLIT distance="1450" swimtime="00:24:08.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="101806" nation="POL" clubid="6811" name="Towarzystwo Sportowe Wisła Kraków">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Krokoszyński" birthdate="1930-05-04" gender="M" nation="POL" license="501806700062" swrid="4302634" athleteid="6812">
              <RESULTS>
                <RESULT eventid="6077" points="427" reactiontime="+121" swimtime="00:00:57.30" resultid="6813" heatid="11404" lane="2" entrytime="00:00:58.07" />
                <RESULT eventid="6238" points="396" reactiontime="+87" swimtime="00:01:12.50" resultid="6814" heatid="11444" lane="1" entrytime="00:01:05.70" />
                <RESULT eventid="6306" points="400" reactiontime="+125" swimtime="00:02:09.12" resultid="6815" heatid="11468" lane="9" entrytime="00:01:58.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="286" reactiontime="+113" swimtime="00:02:56.96" resultid="6816" heatid="11515" lane="0" entrytime="00:02:40.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="6817" heatid="11548" lane="6" entrytime="00:04:10.78" />
                <RESULT eventid="6535" points="315" swimtime="00:05:04.15" resultid="6818" heatid="11562" lane="4" entrytime="00:04:12.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.09" />
                    <SPLIT distance="100" swimtime="00:02:20.14" />
                    <SPLIT distance="150" swimtime="00:03:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7471" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dawid" lastname="Teodorczyk" birthdate="1985-01-01" gender="M" nation="POL" athleteid="7470">
              <RESULTS>
                <RESULT eventid="6077" points="520" swimtime="00:00:27.39" resultid="7472" heatid="11403" lane="1" />
                <RESULT eventid="6340" points="541" reactiontime="+79" swimtime="00:01:09.70" resultid="7473" heatid="11488" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7474" heatid="11530" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8411" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Koba-Gołaszewska" birthdate="1986-01-01" gender="F" nation="POL" athleteid="8410">
              <RESULTS>
                <RESULT eventid="6059" points="584" reactiontime="+77" swimtime="00:00:31.31" resultid="8412" heatid="11399" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="6289" points="528" reactiontime="+81" swimtime="00:01:11.46" resultid="8413" heatid="11465" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="447" reactiontime="+86" swimtime="00:00:37.18" resultid="8414" heatid="11526" lane="7" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8423" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Musiałowski" birthdate="1995-01-01" gender="M" nation="POL" swrid="4258691" athleteid="8422">
              <RESULTS>
                <RESULT eventid="6077" points="719" reactiontime="+71" swimtime="00:00:25.49" resultid="8424" heatid="11416" lane="3" entrytime="00:00:25.86" />
                <RESULT eventid="6111" points="617" reactiontime="+74" swimtime="00:02:21.57" resultid="8425" heatid="11433" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="649" reactiontime="+74" swimtime="00:00:56.09" resultid="8426" heatid="11477" lane="5" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="683" reactiontime="+75" swimtime="00:01:02.66" resultid="8427" heatid="11497" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="635" reactiontime="+79" swimtime="00:01:12.16" resultid="8428" heatid="11520" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="695" reactiontime="+70" swimtime="00:00:26.75" resultid="8429" heatid="11541" lane="4" entrytime="00:00:26.40" />
                <RESULT eventid="6636" points="728" reactiontime="+74" swimtime="00:00:59.93" resultid="8430" heatid="11596" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="618" reactiontime="+75" swimtime="00:00:33.17" resultid="8431" heatid="11621" lane="3" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8538" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jędrzej" lastname="Karpisz" birthdate="1999-01-01" gender="M" nation="POL" swrid="4641502" athleteid="8537">
              <RESULTS>
                <RESULT eventid="6238" points="433" reactiontime="+70" swimtime="00:00:33.61" resultid="8539" heatid="11446" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="6272" points="446" swimtime="00:02:59.34" resultid="8540" heatid="11460" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:21.48" />
                    <SPLIT distance="150" swimtime="00:02:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="529" reactiontime="+68" swimtime="00:01:16.31" resultid="8541" heatid="11519" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="383" reactiontime="+74" swimtime="00:01:15.44" resultid="8542" heatid="11552" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="594" reactiontime="+68" swimtime="00:00:33.61" resultid="8543" heatid="11621" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8544" heatid="11636" lane="6" entrytime="00:04:57.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UKGRO" nation="POL" clubid="7065" name="UKS Sparta Grodzisk Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Jarosław" lastname="Plich" birthdate="1978-06-21" gender="M" nation="POL" athleteid="7077">
              <RESULTS>
                <RESULT eventid="6238" points="472" reactiontime="+89" swimtime="00:00:34.85" resultid="7078" heatid="11448" lane="0" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="6340" points="474" reactiontime="+82" swimtime="00:01:16.67" resultid="7079" heatid="11492" lane="6" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="444" reactiontime="+107" swimtime="00:01:17.40" resultid="7080" heatid="11551" lane="3" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="428" reactiontime="+110" swimtime="00:02:53.11" resultid="7081" heatid="11604" lane="8" entrytime="00:02:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:26.84" />
                    <SPLIT distance="150" swimtime="00:02:12.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Głowa" birthdate="1979-10-08" gender="M" nation="POL" athleteid="7082">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="6306" reactiontime="+65" status="DSQ" swimtime="00:00:00.00" resultid="7083" heatid="11474" lane="2" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="576" swimtime="00:02:15.84" resultid="7084" heatid="11568" lane="4" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="477" reactiontime="+97" swimtime="00:01:12.42" resultid="7085" heatid="11594" lane="8" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Zieliński" birthdate="1980-05-18" gender="M" nation="POL" athleteid="7066">
              <RESULTS>
                <RESULT eventid="6340" points="534" reactiontime="+96" swimtime="00:01:13.71" resultid="7067" heatid="11493" lane="2" entrytime="00:01:12.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="539" reactiontime="+88" swimtime="00:01:18.10" resultid="7068" heatid="11519" lane="4" entrytime="00:01:17.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="578" reactiontime="+74" swimtime="00:00:34.91" resultid="7069" heatid="11620" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="6272" points="550" reactiontime="+87" swimtime="00:02:54.39" resultid="11377" heatid="11455" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:22.59" />
                    <SPLIT distance="150" swimtime="00:02:07.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Milewski" birthdate="1992-03-04" gender="M" nation="POL" swrid="4124793" athleteid="7070">
              <RESULTS>
                <RESULT eventid="6077" points="620" reactiontime="+79" swimtime="00:00:25.95" resultid="7071" heatid="11417" lane="6" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="6111" points="446" reactiontime="+84" swimtime="00:02:34.56" resultid="7072" heatid="11432" lane="0" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:59.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="631" swimtime="00:00:57.16" resultid="7073" heatid="11477" lane="4" entrytime="00:00:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="527" reactiontime="+87" swimtime="00:00:28.31" resultid="7074" heatid="11541" lane="7" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="6535" points="505" reactiontime="+91" swimtime="00:02:13.75" resultid="7075" heatid="11570" lane="7" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:01:00.88" />
                    <SPLIT distance="150" swimtime="00:01:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="471" reactiontime="+84" swimtime="00:01:07.63" resultid="7076" heatid="11595" lane="8" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+87" swimtime="00:01:50.11" resultid="9863" heatid="11584" lane="1" entrytime="00:01:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="100" swimtime="00:00:55.02" />
                    <SPLIT distance="150" swimtime="00:01:23.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7070" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="7066" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="7077" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="7082" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8568" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-01-01" gender="M" nation="POL" swrid="5435204" athleteid="8567">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G7" eventid="6111" reactiontime="+86" status="DSQ" swimtime="00:00:00.00" resultid="8569" heatid="11427" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                    <SPLIT distance="100" swimtime="00:01:50.01" />
                    <SPLIT distance="150" swimtime="00:02:58.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="349" reactiontime="+94" swimtime="00:27:48.31" resultid="8570" heatid="11653" lane="8" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="100" swimtime="00:01:38.23" />
                    <SPLIT distance="150" swimtime="00:02:31.96" />
                    <SPLIT distance="200" swimtime="00:03:26.07" />
                    <SPLIT distance="250" swimtime="00:04:20.91" />
                    <SPLIT distance="300" swimtime="00:05:16.14" />
                    <SPLIT distance="350" swimtime="00:06:10.36" />
                    <SPLIT distance="400" swimtime="00:07:04.59" />
                    <SPLIT distance="450" swimtime="00:07:58.94" />
                    <SPLIT distance="500" swimtime="00:08:52.78" />
                    <SPLIT distance="550" swimtime="00:09:46.65" />
                    <SPLIT distance="600" swimtime="00:10:41.00" />
                    <SPLIT distance="650" swimtime="00:11:35.18" />
                    <SPLIT distance="700" swimtime="00:12:29.57" />
                    <SPLIT distance="750" swimtime="00:13:23.76" />
                    <SPLIT distance="800" swimtime="00:14:19.34" />
                    <SPLIT distance="850" swimtime="00:16:12.28" />
                    <SPLIT distance="900" swimtime="00:17:09.02" />
                    <SPLIT distance="950" swimtime="00:18:05.69" />
                    <SPLIT distance="1000" swimtime="00:19:01.63" />
                    <SPLIT distance="1050" swimtime="00:20:55.88" />
                    <SPLIT distance="1100" swimtime="00:21:53.72" />
                    <SPLIT distance="1150" swimtime="00:22:51.04" />
                    <SPLIT distance="1200" swimtime="00:23:49.67" />
                    <SPLIT distance="1250" swimtime="00:24:48.77" />
                    <SPLIT distance="1300" swimtime="00:25:47.78" />
                    <SPLIT distance="1350" swimtime="00:26:49.37" />
                    <SPLIT distance="1400" swimtime="00:27:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="205" swimtime="00:01:55.62" resultid="8571" heatid="11489" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="315" reactiontime="+130" swimtime="00:03:54.56" resultid="8572" heatid="11502" lane="9" entrytime="00:03:50.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:49.94" />
                    <SPLIT distance="150" swimtime="00:02:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="6467" reactiontime="+92" status="DSQ" swimtime="00:00:41.28" resultid="8573" heatid="11532" lane="5" entrytime="00:00:41.75" entrycourse="SCM" />
                <RESULT eventid="6569" points="228" reactiontime="+91" swimtime="00:08:50.23" resultid="8574" heatid="11576" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                    <SPLIT distance="100" swimtime="00:01:54.99" />
                    <SPLIT distance="150" swimtime="00:03:11.44" />
                    <SPLIT distance="200" swimtime="00:04:28.92" />
                    <SPLIT distance="250" swimtime="00:05:44.90" />
                    <SPLIT distance="300" swimtime="00:07:01.63" />
                    <SPLIT distance="350" swimtime="00:07:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="248" reactiontime="+108" swimtime="00:01:47.16" resultid="8575" heatid="11591" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8576" heatid="11631" lane="3" entrytime="00:06:54.51" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="9454" name="Towarzystwo Pływackie ,,Masters&apos;&apos; Opole">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" license="100607700003" swrid="4843497" athleteid="9455">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6077" points="975" reactiontime="+76" swimtime="00:00:27.06" resultid="9456" heatid="11402" lane="3" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6238" points="1063" reactiontime="+65" swimtime="00:00:30.77" resultid="9457" heatid="11449" lane="9" entrytime="00:00:31.17" entrycourse="SCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6501" points="1101" reactiontime="+62" swimtime="00:01:05.46" resultid="9458" heatid="11552" lane="6" entrytime="00:01:07.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6670" points="1320" reactiontime="+64" swimtime="00:02:23.12" resultid="9459" heatid="11606" lane="6" entrytime="00:02:24.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:46.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Vogel" birthdate="1981-09-20" gender="M" nation="POL" license="100607700016" swrid="5506641" athleteid="9460">
              <RESULTS>
                <RESULT eventid="6340" points="617" reactiontime="+73" swimtime="00:01:10.23" resultid="9461" heatid="11488" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="659" reactiontime="+75" swimtime="00:00:28.87" resultid="9462" heatid="11538" lane="3" entrytime="00:00:29.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7092" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Babica" birthdate="1979-01-01" gender="F" nation="POL" athleteid="7091">
              <RESULTS>
                <RESULT eventid="6094" points="557" reactiontime="+99" swimtime="00:02:58.41" resultid="7093" heatid="11422" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:19.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="601" reactiontime="+96" swimtime="00:22:07.56" resultid="7094" heatid="11650" lane="8" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:16.88" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                    <SPLIT distance="200" swimtime="00:02:42.67" />
                    <SPLIT distance="250" swimtime="00:03:26.43" />
                    <SPLIT distance="300" swimtime="00:04:10.28" />
                    <SPLIT distance="350" swimtime="00:04:54.17" />
                    <SPLIT distance="400" swimtime="00:05:38.72" />
                    <SPLIT distance="450" swimtime="00:06:23.39" />
                    <SPLIT distance="500" swimtime="00:07:07.80" />
                    <SPLIT distance="550" swimtime="00:07:52.37" />
                    <SPLIT distance="600" swimtime="00:08:36.88" />
                    <SPLIT distance="650" swimtime="00:09:21.59" />
                    <SPLIT distance="700" swimtime="00:10:06.79" />
                    <SPLIT distance="750" swimtime="00:10:51.55" />
                    <SPLIT distance="800" swimtime="00:11:36.72" />
                    <SPLIT distance="850" swimtime="00:12:21.98" />
                    <SPLIT distance="900" swimtime="00:13:07.02" />
                    <SPLIT distance="950" swimtime="00:13:52.70" />
                    <SPLIT distance="1000" swimtime="00:14:37.70" />
                    <SPLIT distance="1050" swimtime="00:15:23.41" />
                    <SPLIT distance="1100" swimtime="00:16:09.19" />
                    <SPLIT distance="1150" swimtime="00:16:55.00" />
                    <SPLIT distance="1200" swimtime="00:17:40.91" />
                    <SPLIT distance="1250" swimtime="00:18:25.83" />
                    <SPLIT distance="1300" swimtime="00:19:11.47" />
                    <SPLIT distance="1350" swimtime="00:19:56.32" />
                    <SPLIT distance="1400" swimtime="00:20:41.99" />
                    <SPLIT distance="1450" swimtime="00:21:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="402" reactiontime="+106" swimtime="00:01:27.51" resultid="7095" heatid="11586" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="564" reactiontime="+95" swimtime="00:05:35.14" resultid="7096" heatid="11626" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                    <SPLIT distance="200" swimtime="00:02:42.55" />
                    <SPLIT distance="250" swimtime="00:03:26.42" />
                    <SPLIT distance="300" swimtime="00:04:09.94" />
                    <SPLIT distance="350" swimtime="00:04:53.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8505" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Kotulski" birthdate="1981-01-01" gender="M" nation="POL" athleteid="8504">
              <RESULTS>
                <RESULT eventid="6077" points="433" swimtime="00:00:30.67" resultid="8506" heatid="11408" lane="4" entrytime="00:00:33.10" />
                <RESULT eventid="6306" points="322" swimtime="00:01:14.80" resultid="8507" heatid="11471" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="261" reactiontime="+77" swimtime="00:02:56.70" resultid="8508" heatid="11564" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:02:09.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8482" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Opałko" birthdate="1999-01-01" gender="F" nation="POL" swrid="4493246" athleteid="8481">
              <RESULTS>
                <RESULT eventid="6059" points="570" reactiontime="+77" swimtime="00:00:31.37" resultid="8483" heatid="11399" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="6094" points="470" reactiontime="+79" swimtime="00:02:57.54" resultid="8484" heatid="11423" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:13.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="486" reactiontime="+73" swimtime="00:00:36.87" resultid="8485" heatid="11440" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="6323" points="544" reactiontime="+76" swimtime="00:01:17.38" resultid="8486" heatid="11485" lane="1" entrytime="00:01:18.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="500" swimtime="00:00:35.10" resultid="8487" heatid="11527" lane="8" entrytime="00:00:33.72" entrycourse="SCM" />
                <RESULT eventid="6552" points="428" reactiontime="+82" swimtime="00:06:40.24" resultid="8488" heatid="11574" lane="3" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:30.05" />
                    <SPLIT distance="150" swimtime="00:02:21.72" />
                    <SPLIT distance="200" swimtime="00:03:13.45" />
                    <SPLIT distance="250" swimtime="00:04:07.32" />
                    <SPLIT distance="300" swimtime="00:05:03.89" />
                    <SPLIT distance="350" swimtime="00:05:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="361" swimtime="00:01:27.21" resultid="8489" heatid="11588" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="545" reactiontime="+80" swimtime="00:00:39.79" resultid="8490" heatid="11611" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8376" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Mela" birthdate="1984-01-01" gender="M" nation="POL" athleteid="8375">
              <RESULTS>
                <RESULT eventid="6077" points="346" reactiontime="+86" swimtime="00:00:31.38" resultid="8377" heatid="11407" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="6169" reactiontime="+114" status="OTL" swimtime="00:00:00.00" resultid="8378" heatid="11646" lane="2" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:08.09" />
                    <SPLIT distance="550" swimtime="00:09:19.23" />
                    <SPLIT distance="700" swimtime="00:10:54.84" />
                    <SPLIT distance="750" swimtime="00:11:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="321" reactiontime="+97" swimtime="00:01:12.09" resultid="8379" heatid="11473" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="330" reactiontime="+88" swimtime="00:02:41.15" resultid="8380" heatid="11566" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="327" reactiontime="+90" swimtime="00:05:51.76" resultid="8381" heatid="11634" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:03.45" />
                    <SPLIT distance="200" swimtime="00:02:48.58" />
                    <SPLIT distance="250" swimtime="00:03:34.14" />
                    <SPLIT distance="300" swimtime="00:04:20.75" />
                    <SPLIT distance="350" swimtime="00:05:07.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7509" name="Weteran Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" license="102611600016" swrid="4792005" athleteid="7549">
              <RESULTS>
                <RESULT eventid="6145" points="772" reactiontime="+84" swimtime="00:10:37.70" resultid="7550" heatid="11643" lane="5" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:02:35.84" />
                    <SPLIT distance="250" swimtime="00:03:15.55" />
                    <SPLIT distance="300" swimtime="00:03:55.91" />
                    <SPLIT distance="350" swimtime="00:04:36.12" />
                    <SPLIT distance="400" swimtime="00:05:16.46" />
                    <SPLIT distance="450" swimtime="00:05:56.89" />
                    <SPLIT distance="500" swimtime="00:06:37.24" />
                    <SPLIT distance="550" swimtime="00:07:17.49" />
                    <SPLIT distance="600" swimtime="00:07:57.86" />
                    <SPLIT distance="650" swimtime="00:08:38.05" />
                    <SPLIT distance="700" swimtime="00:09:18.58" />
                    <SPLIT distance="750" swimtime="00:09:58.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" status="DNS" swimtime="00:00:00.00" resultid="7551" heatid="11454" lane="7" entrytime="00:03:06.00" />
                <RESULT eventid="6289" points="662" swimtime="00:01:09.91" resultid="7552" heatid="11465" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="758" reactiontime="+72" swimtime="00:02:26.86" resultid="7553" heatid="11559" lane="8" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:50.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6721" points="805" swimtime="00:05:07.78" resultid="7554" heatid="11628" lane="8" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                    <SPLIT distance="200" swimtime="00:02:31.83" />
                    <SPLIT distance="250" swimtime="00:03:11.30" />
                    <SPLIT distance="300" swimtime="00:03:50.97" />
                    <SPLIT distance="350" swimtime="00:04:30.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" license="102611700035" swrid="5464152" athleteid="7521">
              <RESULTS>
                <RESULT eventid="6077" points="485" reactiontime="+94" swimtime="00:00:35.10" resultid="7522" heatid="11406" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="6169" points="463" swimtime="00:13:35.75" resultid="7523" heatid="11647" lane="1" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:14.15" />
                    <SPLIT distance="200" swimtime="00:03:03.72" />
                    <SPLIT distance="250" swimtime="00:03:53.48" />
                    <SPLIT distance="300" swimtime="00:04:44.35" />
                    <SPLIT distance="400" swimtime="00:06:27.82" />
                    <SPLIT distance="450" swimtime="00:07:19.88" />
                    <SPLIT distance="500" swimtime="00:08:13.28" />
                    <SPLIT distance="550" swimtime="00:09:07.17" />
                    <SPLIT distance="600" swimtime="00:10:01.81" />
                    <SPLIT distance="650" swimtime="00:10:57.20" />
                    <SPLIT distance="700" swimtime="00:11:50.54" />
                    <SPLIT distance="750" swimtime="00:12:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="447" reactiontime="+74" swimtime="00:00:43.57" resultid="7524" heatid="11445" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="6306" points="486" swimtime="00:01:17.68" resultid="7525" heatid="11470" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="430" reactiontime="+78" swimtime="00:01:35.86" resultid="7526" heatid="11549" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="497" reactiontime="+90" swimtime="00:02:55.96" resultid="7527" heatid="11564" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:02:09.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="400" reactiontime="+79" swimtime="00:03:33.91" resultid="7528" heatid="11603" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                    <SPLIT distance="100" swimtime="00:01:42.93" />
                    <SPLIT distance="150" swimtime="00:02:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="512" reactiontime="+106" swimtime="00:06:21.14" resultid="7529" heatid="11632" lane="7" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:02:12.48" />
                    <SPLIT distance="200" swimtime="00:03:01.82" />
                    <SPLIT distance="250" swimtime="00:03:51.62" />
                    <SPLIT distance="300" swimtime="00:04:41.57" />
                    <SPLIT distance="350" swimtime="00:05:32.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" license="102611600029" swrid="5464154" athleteid="7535">
              <RESULTS>
                <RESULT eventid="6059" points="218" swimtime="00:00:55.32" resultid="7536" heatid="11395" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="6220" points="285" reactiontime="+77" swimtime="00:01:03.48" resultid="7537" heatid="11439" lane="0" entrytime="00:01:12.00" />
                <RESULT eventid="6289" points="208" swimtime="00:02:05.95" resultid="7538" heatid="11463" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="236" reactiontime="+77" swimtime="00:02:24.01" resultid="7539" heatid="11544" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="239" swimtime="00:04:30.15" resultid="7540" heatid="11555" lane="4" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:02:09.83" />
                    <SPLIT distance="150" swimtime="00:03:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="267" reactiontime="+83" swimtime="00:05:07.14" resultid="7541" heatid="11599" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.47" />
                    <SPLIT distance="100" swimtime="00:02:33.56" />
                    <SPLIT distance="150" swimtime="00:03:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="306" swimtime="00:09:23.33" resultid="7542" heatid="11625" lane="9" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.82" />
                    <SPLIT distance="100" swimtime="00:02:11.34" />
                    <SPLIT distance="150" swimtime="00:03:24.87" />
                    <SPLIT distance="200" swimtime="00:04:37.15" />
                    <SPLIT distance="250" swimtime="00:05:49.46" />
                    <SPLIT distance="300" swimtime="00:07:00.95" />
                    <SPLIT distance="350" swimtime="00:08:12.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" license="102611700032" swrid="4792004" athleteid="7530">
              <RESULTS>
                <RESULT eventid="6238" points="477" reactiontime="+88" swimtime="00:00:46.57" resultid="7531" heatid="11445" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="6467" points="424" reactiontime="+87" swimtime="00:00:45.23" resultid="7532" heatid="11532" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="6501" points="462" reactiontime="+83" swimtime="00:01:45.57" resultid="7533" heatid="11549" lane="2" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="474" reactiontime="+84" swimtime="00:03:51.01" resultid="7534" heatid="11602" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                    <SPLIT distance="100" swimtime="00:01:50.29" />
                    <SPLIT distance="150" swimtime="00:02:51.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-18" gender="F" nation="POL" license="102611600033" swrid="4655173" athleteid="7543">
              <RESULTS>
                <RESULT eventid="6059" points="239" swimtime="00:00:53.67" resultid="7544" heatid="11396" lane="9" entrytime="00:00:56.00" />
                <RESULT eventid="6255" points="266" swimtime="00:05:31.40" resultid="7545" heatid="11452" lane="0" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.54" />
                    <SPLIT distance="100" swimtime="00:02:39.98" />
                    <SPLIT distance="150" swimtime="00:04:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="216" swimtime="00:02:18.89" resultid="7546" heatid="11482" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="243" reactiontime="+91" swimtime="00:02:35.47" resultid="7547" heatid="11509" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="297" swimtime="00:01:04.67" resultid="7548" heatid="11609" lane="1" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wjciech" lastname="Kosiak" birthdate="1940-04-20" gender="M" nation="POL" license="102611700027" athleteid="7515">
              <RESULTS>
                <RESULT eventid="6077" points="332" reactiontime="+94" swimtime="00:00:46.27" resultid="7516" heatid="11405" lane="9" entrytime="00:00:44.47" />
                <RESULT eventid="6306" points="321" reactiontime="+96" swimtime="00:01:47.62" resultid="7517" heatid="11468" lane="2" entrytime="00:01:44.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7518" heatid="11531" lane="5" entrytime="00:01:07.00" />
                <RESULT eventid="6535" points="302" reactiontime="+111" swimtime="00:04:08.11" resultid="7519" heatid="11563" lane="9" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.31" />
                    <SPLIT distance="100" swimtime="00:02:04.29" />
                    <SPLIT distance="150" swimtime="00:03:10.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="355" reactiontime="+100" swimtime="00:08:28.53" resultid="7520" heatid="11630" lane="3" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.68" />
                    <SPLIT distance="100" swimtime="00:02:03.27" />
                    <SPLIT distance="150" swimtime="00:03:09.68" />
                    <SPLIT distance="200" swimtime="00:04:15.01" />
                    <SPLIT distance="250" swimtime="00:05:20.27" />
                    <SPLIT distance="300" swimtime="00:06:25.79" />
                    <SPLIT distance="350" swimtime="00:07:30.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" license="102611700015" swrid="4137183" athleteid="7510">
              <RESULTS>
                <RESULT eventid="6077" points="595" reactiontime="+87" swimtime="00:00:33.76" resultid="7511" heatid="11409" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="6306" points="519" reactiontime="+88" swimtime="00:01:20.39" resultid="7512" heatid="11470" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="598" reactiontime="+90" swimtime="00:00:38.00" resultid="7513" heatid="11534" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="6704" points="417" reactiontime="+91" swimtime="00:00:47.54" resultid="7514" heatid="11616" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+101" swimtime="00:02:32.26" resultid="9912" heatid="11583" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7521" number="1" reactiontime="+101" />
                    <RELAYPOSITION athleteid="7530" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="7515" number="3" />
                    <RELAYPOSITION athleteid="7510" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+84" swimtime="00:02:59.83" resultid="9913" heatid="12331" lane="1" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:15.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7521" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="7510" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="7530" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7515" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" clubid="7020" name="UKS ENERGETYK Zgorzelec">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Daszyński" birthdate="1948-11-29" gender="M" nation="POL" swrid="4361205" athleteid="7021">
              <RESULTS>
                <RESULT eventid="6111" points="284" reactiontime="+99" swimtime="00:04:30.34" resultid="7022" heatid="11427" lane="7" entrytime="00:04:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.08" />
                    <SPLIT distance="100" swimtime="00:02:13.61" />
                    <SPLIT distance="150" swimtime="00:03:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" points="306" swimtime="00:17:00.00" resultid="7023" heatid="11648" lane="1" entrytime="00:16:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.40" />
                    <SPLIT distance="100" swimtime="00:02:01.13" />
                    <SPLIT distance="150" swimtime="00:03:04.33" />
                    <SPLIT distance="200" swimtime="00:04:08.69" />
                    <SPLIT distance="250" swimtime="00:05:13.00" />
                    <SPLIT distance="300" swimtime="00:06:17.17" />
                    <SPLIT distance="350" swimtime="00:07:21.64" />
                    <SPLIT distance="400" swimtime="00:08:26.19" />
                    <SPLIT distance="450" swimtime="00:09:30.66" />
                    <SPLIT distance="500" swimtime="00:10:35.52" />
                    <SPLIT distance="550" swimtime="00:11:40.48" />
                    <SPLIT distance="600" swimtime="00:12:45.19" />
                    <SPLIT distance="650" swimtime="00:13:49.02" />
                    <SPLIT distance="700" swimtime="00:14:53.92" />
                    <SPLIT distance="750" swimtime="00:15:59.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="274" reactiontime="+95" swimtime="00:00:53.34" resultid="7024" heatid="11444" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="6374" points="177" reactiontime="+100" swimtime="00:05:16.45" resultid="7025" heatid="11501" lane="8" entrytime="00:05:15.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.93" />
                    <SPLIT distance="100" swimtime="00:02:32.73" />
                    <SPLIT distance="150" swimtime="00:03:57.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="279" reactiontime="+89" swimtime="00:01:54.84" resultid="7026" heatid="11549" lane="0" entrytime="00:01:59.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="329" reactiontime="+97" swimtime="00:09:33.61" resultid="7027" heatid="11576" lane="7" entrytime="00:09:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.58" />
                    <SPLIT distance="100" swimtime="00:02:31.17" />
                    <SPLIT distance="150" swimtime="00:03:42.30" />
                    <SPLIT distance="200" swimtime="00:04:51.12" />
                    <SPLIT distance="250" swimtime="00:06:12.81" />
                    <SPLIT distance="300" swimtime="00:07:33.18" />
                    <SPLIT distance="350" swimtime="00:08:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="378" swimtime="00:04:11.63" resultid="7028" heatid="11602" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:03:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="283" reactiontime="+95" swimtime="00:08:19.12" resultid="7029" heatid="11630" lane="5" entrytime="00:08:22.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.38" />
                    <SPLIT distance="100" swimtime="00:01:58.60" />
                    <SPLIT distance="150" swimtime="00:03:03.61" />
                    <SPLIT distance="200" swimtime="00:04:07.78" />
                    <SPLIT distance="250" swimtime="00:05:11.90" />
                    <SPLIT distance="300" swimtime="00:06:15.64" />
                    <SPLIT distance="350" swimtime="00:07:19.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6973" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Jankowski" birthdate="1995-01-01" gender="M" nation="POL" swrid="4112623" athleteid="6972">
              <RESULTS>
                <RESULT eventid="6077" points="881" reactiontime="+68" swimtime="00:00:23.82" resultid="6974" heatid="11418" lane="5" entrytime="00:00:24.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6238" points="887" reactiontime="+61" swimtime="00:00:26.07" resultid="6975" heatid="11450" lane="7" entrytime="00:00:26.50" />
                <RESULT eventid="6306" points="853" reactiontime="+71" swimtime="00:00:51.21" resultid="6976" heatid="11478" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6501" points="929" reactiontime="+59" swimtime="00:00:56.40" resultid="6977" heatid="11553" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="740" reactiontime="+67" swimtime="00:02:08.47" resultid="6978" heatid="11606" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:01.69" />
                    <SPLIT distance="150" swimtime="00:01:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7130" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Sędrowicz" birthdate="1997-01-01" gender="M" nation="POL" swrid="4878673" athleteid="7122">
              <RESULTS>
                <RESULT eventid="6077" points="472" reactiontime="+75" swimtime="00:00:29.32" resultid="7123" heatid="11412" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="6111" points="315" reactiontime="+74" swimtime="00:02:57.12" resultid="7124" heatid="11430" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:23.51" />
                    <SPLIT distance="150" swimtime="00:02:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="432" swimtime="00:03:02.97" resultid="7125" heatid="11458" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                    <SPLIT distance="150" swimtime="00:02:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="7126" heatid="11492" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="6433" points="467" reactiontime="+74" swimtime="00:01:19.93" resultid="7127" heatid="11518" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="380" swimtime="00:00:32.70" resultid="7128" heatid="11535" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="7129" heatid="11601" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02207" nation="POL" region="07" clubid="8784" name="&quot;Masters Zdzieszowice&quot;">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" license="502207600005" swrid="4992846" athleteid="8785">
              <RESULTS>
                <RESULT eventid="6323" points="520" reactiontime="+89" swimtime="00:01:25.94" resultid="8786" heatid="11481" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="396" reactiontime="+92" swimtime="00:03:19.28" resultid="8787" heatid="11498" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:34.80" />
                    <SPLIT distance="150" swimtime="00:02:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="510" reactiontime="+91" swimtime="00:00:37.56" resultid="8788" heatid="11522" lane="3" />
                <RESULT eventid="6552" points="525" swimtime="00:06:40.87" resultid="8789" heatid="11572" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                    <SPLIT distance="150" swimtime="00:02:24.94" />
                    <SPLIT distance="200" swimtime="00:03:14.29" />
                    <SPLIT distance="250" swimtime="00:04:12.23" />
                    <SPLIT distance="300" swimtime="00:05:10.18" />
                    <SPLIT distance="350" swimtime="00:05:57.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="432" reactiontime="+94" swimtime="00:01:27.33" resultid="8790" heatid="11586" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="591" reactiontime="+85" swimtime="00:03:03.17" resultid="8791" heatid="11598" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:17.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8449" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mareks" lastname="Treščinskis" birthdate="1991-01-01" gender="M" nation="POL" athleteid="8448">
              <RESULTS>
                <RESULT eventid="6306" points="496" reactiontime="+73" swimtime="00:01:01.92" resultid="8450" heatid="11476" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="385" reactiontime="+74" swimtime="00:02:26.32" resultid="8451" heatid="11569" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:46.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8525" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Korniak" birthdate="1990-01-01" gender="F" nation="POL" athleteid="8524">
              <RESULTS>
                <RESULT eventid="6059" points="376" swimtime="00:00:35.87" resultid="8526" heatid="11398" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="6220" points="321" reactiontime="+67" swimtime="00:00:43.55" resultid="8527" heatid="11440" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="6289" points="341" reactiontime="+101" swimtime="00:01:22.26" resultid="8528" heatid="11465" lane="7" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="304" reactiontime="+84" swimtime="00:01:42.93" resultid="8529" heatid="11512" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="319" reactiontime="+74" swimtime="00:01:34.09" resultid="8530" heatid="11546" lane="0" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="298" reactiontime="+88" swimtime="00:00:46.91" resultid="8531" heatid="11611" lane="6" entrytime="00:00:40.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8243" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Dusza" birthdate="1983-10-11" gender="F" nation="POL" athleteid="8283">
              <RESULTS>
                <RESULT eventid="6094" points="363" reactiontime="+91" swimtime="00:03:23.58" resultid="8284" heatid="11422" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:37.77" />
                    <SPLIT distance="150" swimtime="00:02:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="421" reactiontime="+95" swimtime="00:24:29.04" resultid="8285" heatid="11650" lane="1" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="150" swimtime="00:02:15.67" />
                    <SPLIT distance="200" swimtime="00:03:03.72" />
                    <SPLIT distance="250" swimtime="00:03:51.31" />
                    <SPLIT distance="300" swimtime="00:04:40.01" />
                    <SPLIT distance="350" swimtime="00:05:28.51" />
                    <SPLIT distance="400" swimtime="00:06:17.11" />
                    <SPLIT distance="450" swimtime="00:07:05.87" />
                    <SPLIT distance="500" swimtime="00:07:54.76" />
                    <SPLIT distance="550" swimtime="00:08:43.69" />
                    <SPLIT distance="600" swimtime="00:09:33.41" />
                    <SPLIT distance="650" swimtime="00:10:23.39" />
                    <SPLIT distance="700" swimtime="00:11:12.94" />
                    <SPLIT distance="750" swimtime="00:12:03.63" />
                    <SPLIT distance="800" swimtime="00:12:53.69" />
                    <SPLIT distance="850" swimtime="00:13:44.22" />
                    <SPLIT distance="900" swimtime="00:14:34.47" />
                    <SPLIT distance="950" swimtime="00:15:24.49" />
                    <SPLIT distance="1000" swimtime="00:16:14.46" />
                    <SPLIT distance="1050" swimtime="00:17:04.21" />
                    <SPLIT distance="1100" swimtime="00:17:54.32" />
                    <SPLIT distance="1150" swimtime="00:18:44.24" />
                    <SPLIT distance="1200" swimtime="00:19:33.91" />
                    <SPLIT distance="1250" swimtime="00:20:23.20" />
                    <SPLIT distance="1300" swimtime="00:21:12.43" />
                    <SPLIT distance="1350" swimtime="00:22:01.53" />
                    <SPLIT distance="1400" swimtime="00:22:51.14" />
                    <SPLIT distance="1450" swimtime="00:23:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="346" reactiontime="+89" swimtime="00:01:22.24" resultid="8286" heatid="11464" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="361" reactiontime="+89" swimtime="00:01:32.90" resultid="8287" heatid="11483" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="387" reactiontime="+91" swimtime="00:02:55.68" resultid="8288" heatid="11557" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:11.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="399" reactiontime="+89" swimtime="00:07:08.65" resultid="8289" heatid="11574" lane="0" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="100" swimtime="00:01:46.50" />
                    <SPLIT distance="150" swimtime="00:02:41.06" />
                    <SPLIT distance="200" swimtime="00:03:33.82" />
                    <SPLIT distance="250" swimtime="00:04:31.19" />
                    <SPLIT distance="300" swimtime="00:05:30.15" />
                    <SPLIT distance="350" swimtime="00:06:20.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="391" reactiontime="+89" swimtime="00:06:13.36" resultid="8290" heatid="11626" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:26.07" />
                    <SPLIT distance="150" swimtime="00:02:13.64" />
                    <SPLIT distance="200" swimtime="00:03:02.18" />
                    <SPLIT distance="250" swimtime="00:03:50.38" />
                    <SPLIT distance="300" swimtime="00:04:38.56" />
                    <SPLIT distance="350" swimtime="00:05:26.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Burandt" birthdate="1972-12-15" gender="F" nation="POL" swrid="5471721" athleteid="8330">
              <RESULTS>
                <RESULT eventid="6289" points="547" reactiontime="+77" swimtime="00:01:14.51" resultid="8331" heatid="11464" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="539" swimtime="00:01:24.84" resultid="8332" heatid="11484" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="589" reactiontime="+86" swimtime="00:00:37.15" resultid="8333" heatid="11525" lane="4" entrytime="00:00:36.78" />
                <RESULT eventid="6518" points="527" swimtime="00:02:45.74" resultid="8334" heatid="11557" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                    <SPLIT distance="150" swimtime="00:02:01.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="474" swimtime="00:00:45.91" resultid="8335" heatid="11611" lane="7" entrytime="00:00:41.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Zwierzyński" birthdate="1960-05-10" gender="M" nation="POL" athleteid="8254">
              <RESULTS>
                <RESULT eventid="6077" points="192" swimtime="00:00:46.48" resultid="8255" heatid="11404" lane="4" entrytime="00:00:47.04" />
                <RESULT eventid="6203" reactiontime="+96" status="OTL" swimtime="00:00:00.00" resultid="8256" heatid="11654" lane="5" entrytime="00:29:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:51.66" />
                    <SPLIT distance="150" swimtime="00:02:56.40" />
                    <SPLIT distance="200" swimtime="00:04:01.71" />
                    <SPLIT distance="250" swimtime="00:05:07.61" />
                    <SPLIT distance="300" swimtime="00:06:14.25" />
                    <SPLIT distance="350" swimtime="00:07:20.87" />
                    <SPLIT distance="400" swimtime="00:08:27.40" />
                    <SPLIT distance="450" swimtime="00:09:33.84" />
                    <SPLIT distance="500" swimtime="00:10:40.17" />
                    <SPLIT distance="550" swimtime="00:11:48.03" />
                    <SPLIT distance="600" swimtime="00:12:54.61" />
                    <SPLIT distance="650" swimtime="00:14:02.14" />
                    <SPLIT distance="700" swimtime="00:15:07.84" />
                    <SPLIT distance="750" swimtime="00:16:14.19" />
                    <SPLIT distance="800" swimtime="00:17:19.27" />
                    <SPLIT distance="850" swimtime="00:18:26.94" />
                    <SPLIT distance="900" swimtime="00:19:34.20" />
                    <SPLIT distance="950" swimtime="00:20:45.58" />
                    <SPLIT distance="1000" swimtime="00:21:54.07" />
                    <SPLIT distance="1050" swimtime="00:23:01.53" />
                    <SPLIT distance="1100" swimtime="00:24:06.36" />
                    <SPLIT distance="1150" swimtime="00:25:13.39" />
                    <SPLIT distance="1200" swimtime="00:26:22.03" />
                    <SPLIT distance="1250" swimtime="00:27:31.28" />
                    <SPLIT distance="1300" swimtime="00:28:37.39" />
                    <SPLIT distance="1350" swimtime="00:29:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="214" reactiontime="+78" swimtime="00:04:37.00" resultid="8257" heatid="11456" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.05" />
                    <SPLIT distance="100" swimtime="00:02:08.93" />
                    <SPLIT distance="150" swimtime="00:03:24.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="172" reactiontime="+90" swimtime="00:01:47.53" resultid="8258" heatid="11468" lane="8" entrytime="00:01:49.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="204" reactiontime="+110" swimtime="00:02:05.39" resultid="8259" heatid="11515" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="182" reactiontime="+84" swimtime="00:04:00.83" resultid="8260" heatid="11563" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:53.06" />
                    <SPLIT distance="150" swimtime="00:02:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="223" reactiontime="+78" swimtime="00:00:53.95" resultid="8261" heatid="11616" lane="9" entrytime="00:00:56.27" />
                <RESULT eventid="6738" points="186" reactiontime="+83" swimtime="00:08:29.99" resultid="8262" heatid="11631" lane="9" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                    <SPLIT distance="100" swimtime="00:01:56.65" />
                    <SPLIT distance="150" swimtime="00:03:00.70" />
                    <SPLIT distance="200" swimtime="00:04:07.00" />
                    <SPLIT distance="250" swimtime="00:05:14.86" />
                    <SPLIT distance="300" swimtime="00:06:20.92" />
                    <SPLIT distance="350" swimtime="00:07:26.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Chudoba" birthdate="1981-03-04" gender="M" nation="POL" athleteid="8250">
              <RESULTS>
                <RESULT eventid="6374" points="492" reactiontime="+91" swimtime="00:02:39.67" resultid="8251" heatid="11503" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:13.68" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="674" swimtime="00:00:28.65" resultid="8252" heatid="11539" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="6636" points="664" swimtime="00:01:04.87" resultid="8253" heatid="11595" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Bałtóg" birthdate="1972-03-11" gender="F" nation="POL" athleteid="8324">
              <RESULTS>
                <RESULT eventid="6289" points="565" swimtime="00:01:13.71" resultid="8325" heatid="11464" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="532" reactiontime="+84" swimtime="00:01:25.20" resultid="8326" heatid="11483" lane="1" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="556" reactiontime="+80" swimtime="00:00:37.88" resultid="8327" heatid="11525" lane="3" entrytime="00:00:37.53" />
                <RESULT eventid="6518" points="470" swimtime="00:02:52.18" resultid="8328" heatid="11559" lane="9" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="461" reactiontime="+89" swimtime="00:01:27.49" resultid="8329" heatid="11587" lane="8" entrytime="00:01:28.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Chojcan" birthdate="1986-08-04" gender="F" nation="POL" athleteid="8297">
              <RESULTS>
                <RESULT eventid="6094" points="642" reactiontime="+79" swimtime="00:02:48.38" resultid="8298" heatid="11423" lane="7" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:02:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="520" reactiontime="+85" swimtime="00:11:43.80" resultid="8299" heatid="11643" lane="7" entrytime="00:11:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="150" swimtime="00:02:00.69" />
                    <SPLIT distance="200" swimtime="00:02:44.71" />
                    <SPLIT distance="250" swimtime="00:03:29.24" />
                    <SPLIT distance="300" swimtime="00:04:14.30" />
                    <SPLIT distance="350" swimtime="00:04:59.29" />
                    <SPLIT distance="400" swimtime="00:05:44.54" />
                    <SPLIT distance="450" swimtime="00:06:29.76" />
                    <SPLIT distance="500" swimtime="00:07:15.21" />
                    <SPLIT distance="550" swimtime="00:08:00.43" />
                    <SPLIT distance="600" swimtime="00:08:45.50" />
                    <SPLIT distance="650" swimtime="00:09:30.42" />
                    <SPLIT distance="700" swimtime="00:10:15.31" />
                    <SPLIT distance="750" swimtime="00:11:00.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="658" reactiontime="+66" swimtime="00:00:35.51" resultid="8300" heatid="11440" lane="3" entrytime="00:00:35.67" />
                <RESULT eventid="6357" points="457" reactiontime="+87" swimtime="00:03:05.07" resultid="8301" heatid="11499" lane="2" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:23.77" />
                    <SPLIT distance="150" swimtime="00:02:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="562" reactiontime="+75" swimtime="00:00:34.46" resultid="8302" heatid="11526" lane="2" entrytime="00:00:35.27" />
                <RESULT eventid="6484" points="667" reactiontime="+70" swimtime="00:01:15.45" resultid="8303" heatid="11546" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="537" swimtime="00:01:18.43" resultid="8304" heatid="11587" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="608" reactiontime="+72" swimtime="00:02:48.51" resultid="8305" heatid="11600" lane="2" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:02:04.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Podulka" birthdate="1975-09-29" gender="F" nation="POL" athleteid="8312">
              <RESULTS>
                <RESULT eventid="6059" points="585" reactiontime="+87" swimtime="00:00:32.16" resultid="8313" heatid="11399" lane="0" entrytime="00:00:32.32" />
                <RESULT eventid="6289" points="476" reactiontime="+99" swimtime="00:01:16.37" resultid="8314" heatid="11464" lane="6" entrytime="00:01:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="561" reactiontime="+90" swimtime="00:00:36.38" resultid="8315" heatid="11525" lane="6" entrytime="00:00:37.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Kolenkiewicz" birthdate="1977-12-13" gender="M" nation="POL" athleteid="8263">
              <RESULTS>
                <RESULT eventid="6111" points="679" reactiontime="+75" swimtime="00:02:30.59" resultid="8264" heatid="11432" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="688" reactiontime="+88" swimtime="00:02:47.25" resultid="8265" heatid="11459" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:02:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="690" reactiontime="+93" swimtime="00:01:14.74" resultid="8266" heatid="11519" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="673" reactiontime="+81" swimtime="00:00:34.55" resultid="8267" heatid="11620" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radosław" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" swrid="4429483" athleteid="8278">
              <RESULTS>
                <RESULT eventid="6272" points="511" reactiontime="+77" swimtime="00:03:04.61" resultid="8279" heatid="11458" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="489" reactiontime="+99" swimtime="00:01:23.85" resultid="8280" heatid="11519" lane="9" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="358" reactiontime="+97" swimtime="00:02:41.46" resultid="8281" heatid="11567" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:01:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="526" swimtime="00:00:37.51" resultid="8282" heatid="11620" lane="0" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Bąkowski" birthdate="1984-06-20" gender="M" nation="POL" athleteid="8244">
              <RESULTS>
                <RESULT eventid="6077" points="413" reactiontime="+89" swimtime="00:00:29.58" resultid="8245" heatid="11412" lane="0" entrytime="00:00:29.30" />
                <RESULT eventid="6238" points="362" reactiontime="+100" swimtime="00:00:34.32" resultid="8246" heatid="11447" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="6340" points="419" reactiontime="+96" swimtime="00:01:15.89" resultid="8247" heatid="11492" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="429" reactiontime="+94" swimtime="00:01:14.13" resultid="8248" heatid="11551" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="415" reactiontime="+88" swimtime="00:02:42.93" resultid="8249" heatid="11604" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Krowicka" birthdate="1960-05-11" gender="F" nation="POL" athleteid="8316">
              <RESULTS>
                <RESULT eventid="6059" points="480" reactiontime="+71" swimtime="00:00:39.59" resultid="8317" heatid="11397" lane="2" entrytime="00:00:38.90" />
                <RESULT eventid="6094" points="429" reactiontime="+79" swimtime="00:03:50.96" resultid="8318" heatid="11421" lane="7" entrytime="00:03:48.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                    <SPLIT distance="100" swimtime="00:01:55.64" />
                    <SPLIT distance="150" swimtime="00:02:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="519" swimtime="00:03:53.17" resultid="8319" heatid="11453" lane="9" entrytime="00:03:54.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                    <SPLIT distance="100" swimtime="00:01:51.33" />
                    <SPLIT distance="150" swimtime="00:02:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="468" reactiontime="+79" swimtime="00:01:41.84" resultid="8320" heatid="11483" lane="9" entrytime="00:01:40.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="514" swimtime="00:01:46.29" resultid="8321" heatid="11511" lane="9" entrytime="00:01:45.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="328" swimtime="00:00:48.44" resultid="8322" heatid="11524" lane="6" entrytime="00:00:49.19" />
                <RESULT eventid="6687" points="537" swimtime="00:00:46.88" resultid="8323" heatid="11610" lane="6" entrytime="00:00:47.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Michalczuk" birthdate="1970-03-05" gender="M" nation="POL" athleteid="8272">
              <RESULTS>
                <RESULT eventid="6077" points="417" reactiontime="+70" swimtime="00:00:32.77" resultid="8273" heatid="11409" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="6238" points="229" reactiontime="+84" swimtime="00:00:46.34" resultid="8274" heatid="11446" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="6306" points="368" reactiontime="+74" swimtime="00:01:14.07" resultid="8275" heatid="11472" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="269" reactiontime="+87" swimtime="00:01:31.82" resultid="8276" heatid="11490" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="321" reactiontime="+82" swimtime="00:02:52.40" resultid="8277" heatid="11565" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:10.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Wawrzyńczak" birthdate="1990-09-11" gender="F" nation="POL" swrid="4071814" athleteid="8291">
              <RESULTS>
                <RESULT eventid="6059" points="476" swimtime="00:00:33.17" resultid="8292" heatid="11399" lane="1" entrytime="00:00:31.90" />
                <RESULT eventid="6220" points="587" reactiontime="+77" swimtime="00:00:35.61" resultid="8293" heatid="11441" lane="9" entrytime="00:00:35.50" />
                <RESULT eventid="6450" points="565" reactiontime="+70" swimtime="00:00:34.08" resultid="8294" heatid="11527" lane="1" entrytime="00:00:33.60" />
                <RESULT eventid="6484" points="541" reactiontime="+81" swimtime="00:01:18.89" resultid="8295" heatid="11546" lane="1" entrytime="00:01:17.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="498" reactiontime="+79" swimtime="00:01:18.94" resultid="8296" heatid="11588" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Cwojdzińska" birthdate="1992-12-21" gender="F" nation="POL" swrid="4104697" athleteid="8306">
              <RESULTS>
                <RESULT eventid="6094" points="508" reactiontime="+78" swimtime="00:02:59.07" resultid="8307" heatid="11422" lane="4" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="597" reactiontime="+66" swimtime="00:00:35.41" resultid="8308" heatid="11440" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="6323" points="516" swimtime="00:01:20.78" resultid="8309" heatid="11484" lane="4" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="593" reactiontime="+63" swimtime="00:01:16.54" resultid="8310" heatid="11546" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="574" reactiontime="+67" swimtime="00:02:50.38" resultid="8311" heatid="11600" lane="8" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:05.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Maciaszek" birthdate="1991-05-16" gender="M" nation="POL" athleteid="8268">
              <RESULTS>
                <RESULT eventid="6077" points="631" swimtime="00:00:25.79" resultid="8269" heatid="11416" lane="9" entrytime="00:00:26.07" />
                <RESULT eventid="6340" points="510" reactiontime="+81" swimtime="00:01:08.82" resultid="8270" heatid="11493" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="551" reactiontime="+66" swimtime="00:00:27.89" resultid="8271" heatid="11540" lane="0" entrytime="00:00:28.01" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+91" swimtime="00:01:50.21" resultid="9857" heatid="11584" lane="8" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:00:57.22" />
                    <SPLIT distance="150" swimtime="00:01:25.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8244" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="8250" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="8263" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="8268" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" status="DNS" swimtime="00:00:00.00" resultid="9858" heatid="12332" lane="2" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8244" number="1" />
                    <RELAYPOSITION athleteid="8263" number="2" />
                    <RELAYPOSITION athleteid="8250" number="3" />
                    <RELAYPOSITION athleteid="8268" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+83" swimtime="00:02:12.53" resultid="9859" heatid="11581" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:04.92" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8291" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="8297" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="8306" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="8283" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" status="DNS" swimtime="00:00:00.00" resultid="9860" heatid="11639" lane="6" entrytime="00:02:33.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8297" number="1" />
                    <RELAYPOSITION athleteid="8306" number="2" />
                    <RELAYPOSITION athleteid="8291" number="3" />
                    <RELAYPOSITION athleteid="8283" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="6586" reactiontime="+93" swimtime="00:02:18.32" resultid="9861" heatid="11581" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:44.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8324" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="8312" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="8316" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="8330" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6755" status="DNS" swimtime="00:00:00.00" resultid="9862" heatid="11639" lane="2" entrytime="00:02:42.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8324" number="1" />
                    <RELAYPOSITION athleteid="8316" number="2" />
                    <RELAYPOSITION athleteid="8330" number="3" />
                    <RELAYPOSITION athleteid="8312" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+81" swimtime="00:01:56.36" resultid="9852" heatid="11436" lane="7" entrytime="00:01:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="100" swimtime="00:00:52.54" />
                    <SPLIT distance="150" swimtime="00:01:24.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8250" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="8268" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="8297" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="8306" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+64" swimtime="00:02:09.88" resultid="9853" heatid="11507" lane="2" entrytime="00:02:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:38.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8297" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="8263" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="8250" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="8306" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+79" swimtime="00:02:02.74" resultid="9854" heatid="11436" lane="0" entrytime="00:02:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="100" swimtime="00:01:01.38" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8263" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="8291" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="8312" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="8244" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+88" swimtime="00:02:15.15" resultid="9855" heatid="11505" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                    <SPLIT distance="150" swimtime="00:01:43.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8244" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="8268" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="8291" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="8312" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+80" swimtime="00:02:29.84" resultid="9856" heatid="11506" lane="5" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:01:56.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8324" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="8278" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="8330" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="8272" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="7087" name="The swimming and sport Crazy Fish club">
          <ATHLETES>
            <ATHLETE firstname="Svitlana" lastname="Urbanik" birthdate="1985-07-23" gender="F" nation="UKR" license="Poltava" athleteid="7088">
              <RESULTS>
                <RESULT eventid="6094" status="DNS" swimtime="00:00:00.00" resultid="7089" heatid="11421" lane="0" />
                <RESULT eventid="6255" status="DNS" swimtime="00:00:00.00" resultid="7090" heatid="11451" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="9470" name="UKS ,,Jasień&apos;&apos; Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="9471">
              <RESULTS>
                <RESULT eventid="6059" points="714" reactiontime="+77" swimtime="00:00:29.28" resultid="9472" heatid="11400" lane="3" entrytime="00:00:29.84" entrycourse="SCM" />
                <RESULT eventid="6255" points="581" reactiontime="+80" swimtime="00:03:05.90" resultid="9473" heatid="11454" lane="1" entrytime="00:03:07.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:28.79" />
                    <SPLIT distance="150" swimtime="00:02:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="654" reactiontime="+81" swimtime="00:01:16.23" resultid="9474" heatid="11481" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="594" reactiontime="+82" swimtime="00:01:22.13" resultid="9475" heatid="11512" lane="2" entrytime="00:01:22.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="434" reactiontime="+91" swimtime="00:02:49.21" resultid="9476" heatid="11555" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                    <SPLIT distance="150" swimtime="00:02:05.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="732" reactiontime="+78" swimtime="00:00:35.13" resultid="9477" heatid="11612" lane="6" entrytime="00:00:35.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Pytel" birthdate="1979-02-03" gender="F" nation="POL" license="102706600133" athleteid="9478">
              <RESULTS>
                <RESULT eventid="6059" points="245" swimtime="00:00:41.99" resultid="9479" heatid="11394" lane="4" />
                <RESULT eventid="6220" points="253" reactiontime="+70" swimtime="00:00:48.30" resultid="9480" heatid="11437" lane="5" />
                <RESULT eventid="6415" points="277" reactiontime="+81" swimtime="00:01:56.01" resultid="9481" heatid="11509" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="9482" heatid="11522" lane="5" />
                <RESULT eventid="6687" points="364" reactiontime="+80" swimtime="00:00:48.06" resultid="9483" heatid="11608" lane="1" />
                <RESULT eventid="6255" points="270" swimtime="00:04:16.83" resultid="12233" heatid="11451" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                    <SPLIT distance="100" swimtime="00:02:00.49" />
                    <SPLIT distance="150" swimtime="00:03:07.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8558" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-01-01" gender="F" nation="POL" athleteid="8557">
              <RESULTS>
                <RESULT comment="O2 - Pływak nie miał kontaktu ze ścianą podczas nawrotu." eventid="6094" reactiontime="+98" status="DSQ" swimtime="00:00:00.00" resultid="8559" heatid="11421" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                    <SPLIT distance="100" swimtime="00:01:49.13" />
                    <SPLIT distance="150" swimtime="00:02:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="451" reactiontime="+95" swimtime="00:23:55.94" resultid="8560" heatid="11651" lane="4" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:14.84" />
                    <SPLIT distance="200" swimtime="00:03:02.76" />
                    <SPLIT distance="250" swimtime="00:03:50.29" />
                    <SPLIT distance="300" swimtime="00:04:38.16" />
                    <SPLIT distance="350" swimtime="00:05:26.06" />
                    <SPLIT distance="400" swimtime="00:06:13.80" />
                    <SPLIT distance="450" swimtime="00:07:01.49" />
                    <SPLIT distance="500" swimtime="00:07:49.42" />
                    <SPLIT distance="550" swimtime="00:08:37.31" />
                    <SPLIT distance="600" swimtime="00:09:25.47" />
                    <SPLIT distance="650" swimtime="00:10:13.58" />
                    <SPLIT distance="700" swimtime="00:11:01.70" />
                    <SPLIT distance="750" swimtime="00:11:49.96" />
                    <SPLIT distance="800" swimtime="00:12:38.24" />
                    <SPLIT distance="850" swimtime="00:13:26.20" />
                    <SPLIT distance="900" swimtime="00:14:14.79" />
                    <SPLIT distance="950" swimtime="00:15:03.25" />
                    <SPLIT distance="1000" swimtime="00:15:51.39" />
                    <SPLIT distance="1050" swimtime="00:16:39.39" />
                    <SPLIT distance="1100" swimtime="00:17:27.41" />
                    <SPLIT distance="1150" swimtime="00:18:15.60" />
                    <SPLIT distance="1200" swimtime="00:19:04.36" />
                    <SPLIT distance="1250" swimtime="00:19:53.42" />
                    <SPLIT distance="1300" swimtime="00:20:42.64" />
                    <SPLIT distance="1350" swimtime="00:21:31.39" />
                    <SPLIT distance="1400" swimtime="00:22:20.65" />
                    <SPLIT distance="1450" swimtime="00:23:09.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="311" reactiontime="+95" swimtime="00:01:37.60" resultid="8561" heatid="11482" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="268" reactiontime="+99" swimtime="00:03:41.03" resultid="8562" heatid="11499" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="307" reactiontime="+95" swimtime="00:03:09.73" resultid="8563" heatid="11556" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:20.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="377" reactiontime="+103" swimtime="00:07:16.73" resultid="8564" heatid="11573" lane="3" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                    <SPLIT distance="100" swimtime="00:01:46.89" />
                    <SPLIT distance="150" swimtime="00:02:51.04" />
                    <SPLIT distance="200" swimtime="00:03:54.79" />
                    <SPLIT distance="250" swimtime="00:04:49.24" />
                    <SPLIT distance="300" swimtime="00:05:44.18" />
                    <SPLIT distance="350" swimtime="00:06:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="252" swimtime="00:01:40.83" resultid="8565" heatid="11586" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" status="DNS" swimtime="00:00:00.00" resultid="8566" heatid="11626" lane="1" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9700" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Adrian" lastname="Teodorski" birthdate="1990-01-01" gender="M" nation="POL" swrid="4071733" athleteid="9699">
              <RESULTS>
                <RESULT eventid="6111" points="402" reactiontime="+85" swimtime="00:02:39.98" resultid="9701" heatid="11432" lane="7" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" reactiontime="+84" status="DNF" swimtime="00:00:00.00" resultid="9702" heatid="11652" lane="6" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                    <SPLIT distance="200" swimtime="00:02:32.45" />
                    <SPLIT distance="250" swimtime="00:03:12.55" />
                    <SPLIT distance="300" swimtime="00:03:52.50" />
                    <SPLIT distance="350" swimtime="00:04:32.85" />
                    <SPLIT distance="400" swimtime="00:05:12.86" />
                    <SPLIT distance="450" swimtime="00:05:55.47" />
                    <SPLIT distance="500" swimtime="00:06:17.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" status="DNS" swimtime="00:00:00.00" resultid="9703" heatid="11459" lane="0" entrytime="00:02:55.20" />
                <RESULT eventid="6374" points="337" reactiontime="+92" swimtime="00:02:58.14" resultid="9704" heatid="11504" lane="7" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:24.98" />
                    <SPLIT distance="150" swimtime="00:02:16.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="521" reactiontime="+70" swimtime="00:00:28.41" resultid="9705" heatid="11540" lane="6" entrytime="00:00:27.82" />
                <RESULT eventid="6569" points="461" reactiontime="+97" swimtime="00:05:45.41" resultid="9706" heatid="11579" lane="1" entrytime="00:05:25.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:05.97" />
                    <SPLIT distance="200" swimtime="00:02:48.76" />
                    <SPLIT distance="250" swimtime="00:03:40.04" />
                    <SPLIT distance="300" swimtime="00:04:30.51" />
                    <SPLIT distance="350" swimtime="00:05:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="467" reactiontime="+79" swimtime="00:01:07.79" resultid="9707" heatid="11595" lane="5" entrytime="00:01:03.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="491" reactiontime="+88" swimtime="00:05:04.45" resultid="9708" heatid="11636" lane="2" entrytime="00:04:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                    <SPLIT distance="200" swimtime="00:02:30.24" />
                    <SPLIT distance="250" swimtime="00:03:10.39" />
                    <SPLIT distance="300" swimtime="00:03:50.31" />
                    <SPLIT distance="350" swimtime="00:04:28.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6923" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kubiak" birthdate="1989-01-01" gender="M" nation="POL" athleteid="6922">
              <RESULTS>
                <RESULT eventid="6111" points="203" reactiontime="+111" swimtime="00:03:20.78" resultid="6924" heatid="11429" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="150" swimtime="00:02:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" status="OTL" swimtime="00:00:00.00" resultid="6925" heatid="11645" lane="1" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                    <SPLIT distance="200" swimtime="00:02:42.38" />
                    <SPLIT distance="250" swimtime="00:03:25.44" />
                    <SPLIT distance="300" swimtime="00:04:10.03" />
                    <SPLIT distance="350" swimtime="00:04:52.96" />
                    <SPLIT distance="400" swimtime="00:06:21.14" />
                    <SPLIT distance="450" swimtime="00:07:05.94" />
                    <SPLIT distance="500" swimtime="00:07:49.63" />
                    <SPLIT distance="550" swimtime="00:08:34.05" />
                    <SPLIT distance="600" swimtime="00:09:16.14" />
                    <SPLIT distance="650" swimtime="00:09:58.92" />
                    <SPLIT distance="700" swimtime="00:10:41.95" />
                    <SPLIT distance="750" swimtime="00:11:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="306" reactiontime="+111" swimtime="00:01:12.73" resultid="6926" heatid="11472" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="221" swimtime="00:03:25.07" resultid="6927" heatid="11502" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:37.32" />
                    <SPLIT distance="150" swimtime="00:02:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="219" reactiontime="+108" swimtime="00:00:37.90" resultid="6928" heatid="11534" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="6569" points="250" reactiontime="+107" swimtime="00:07:03.63" resultid="6929" heatid="11577" lane="7" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="150" swimtime="00:02:42.51" />
                    <SPLIT distance="200" swimtime="00:03:37.45" />
                    <SPLIT distance="250" swimtime="00:04:39.29" />
                    <SPLIT distance="300" swimtime="00:05:42.94" />
                    <SPLIT distance="350" swimtime="00:06:22.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="168" swimtime="00:01:35.38" resultid="6930" heatid="11591" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="363" reactiontime="+98" swimtime="00:05:36.76" resultid="6931" heatid="11634" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="150" swimtime="00:02:02.33" />
                    <SPLIT distance="200" swimtime="00:02:45.62" />
                    <SPLIT distance="250" swimtime="00:03:29.46" />
                    <SPLIT distance="300" swimtime="00:04:11.70" />
                    <SPLIT distance="350" swimtime="00:04:54.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6960" name="AQUAPARK WROCŁAW">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Witkowski" birthdate="1984-01-01" gender="M" nation="POL" swrid="4036605" athleteid="6959">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6077" points="778" reactiontime="+76" swimtime="00:00:23.95" resultid="6961" heatid="11403" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00304" nation="POL" clubid="7175" name="Towarzystwo Pływackie Zielona Góra">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Karczewski" birthdate="1974-06-11" gender="M" nation="POL" license="100304700490" swrid="5342868" athleteid="7176">
              <RESULTS>
                <RESULT eventid="6077" points="519" swimtime="00:00:29.70" resultid="7177" heatid="11411" lane="9" entrytime="00:00:30.40" />
                <RESULT eventid="6306" points="521" reactiontime="+78" swimtime="00:01:05.73" resultid="7178" heatid="11473" lane="5" entrytime="00:01:06.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="583" swimtime="00:00:30.74" resultid="7179" heatid="11536" lane="4" entrytime="00:00:31.09" />
                <RESULT eventid="6636" points="540" reactiontime="+80" swimtime="00:01:11.87" resultid="7180" heatid="11592" lane="5" entrytime="00:01:16.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7198" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Mazerant" birthdate="1978-01-10" gender="M" nation="POL" athleteid="7197">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7199" heatid="11408" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7200" heatid="11472" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="7201" heatid="11566" lane="3" entrytime="00:02:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7281" name="MASTERS Zdzieszowice">
          <ATHLETES>
            <ATHLETE firstname="Sasha" lastname="Broshevan" birthdate="1986-08-06" gender="M" nation="POL" athleteid="7282">
              <RESULTS>
                <RESULT eventid="6077" points="524" swimtime="00:00:27.31" resultid="7283" heatid="11415" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="6238" points="455" reactiontime="+75" swimtime="00:00:31.81" resultid="7284" heatid="11448" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="6340" points="452" reactiontime="+82" swimtime="00:01:14.01" resultid="7285" heatid="11493" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="532" reactiontime="+84" swimtime="00:00:29.15" resultid="7286" heatid="11530" lane="3" />
                <RESULT eventid="6501" points="417" reactiontime="+73" swimtime="00:01:14.82" resultid="7287" heatid="11551" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="406" reactiontime="+76" swimtime="00:01:14.50" resultid="7288" heatid="11589" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="495" swimtime="00:00:36.46" resultid="7289" heatid="11620" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6854" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Burzyński" birthdate="1962-01-01" gender="M" nation="POL" athleteid="6853">
              <RESULTS>
                <RESULT eventid="6203" points="359" reactiontime="+140" swimtime="00:27:32.42" resultid="6855" heatid="11653" lane="0" entrytime="00:28:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="350" swimtime="00:07:53.30" />
                    <SPLIT distance="400" swimtime="00:08:47.94" />
                    <SPLIT distance="450" swimtime="00:09:43.05" />
                    <SPLIT distance="600" swimtime="00:10:38.00" />
                    <SPLIT distance="650" swimtime="00:11:33.53" />
                    <SPLIT distance="700" swimtime="00:12:29.82" />
                    <SPLIT distance="750" swimtime="00:13:25.76" />
                    <SPLIT distance="800" swimtime="00:14:22.76" />
                    <SPLIT distance="850" swimtime="00:15:18.11" />
                    <SPLIT distance="900" swimtime="00:16:14.22" />
                    <SPLIT distance="950" swimtime="00:17:11.58" />
                    <SPLIT distance="1000" swimtime="00:18:07.92" />
                    <SPLIT distance="1050" swimtime="00:19:04.34" />
                    <SPLIT distance="1100" swimtime="00:20:01.06" />
                    <SPLIT distance="1150" swimtime="00:20:57.94" />
                    <SPLIT distance="1200" swimtime="00:21:54.44" />
                    <SPLIT distance="1250" swimtime="00:22:51.00" />
                    <SPLIT distance="1300" swimtime="00:23:47.38" />
                    <SPLIT distance="1350" swimtime="00:24:44.08" />
                    <SPLIT distance="1400" swimtime="00:25:40.76" />
                    <SPLIT distance="1450" swimtime="00:26:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="230" reactiontime="+129" swimtime="00:04:20.40" resultid="6856" heatid="11501" lane="7" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                    <SPLIT distance="100" swimtime="00:02:02.26" />
                    <SPLIT distance="150" swimtime="00:03:11.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="226" reactiontime="+122" swimtime="00:01:51.98" resultid="6857" heatid="11490" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="290" reactiontime="+134" swimtime="00:08:08.90" resultid="6858" heatid="11577" lane="9" entrytime="00:07:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:02:01.21" />
                    <SPLIT distance="150" swimtime="00:03:08.96" />
                    <SPLIT distance="200" swimtime="00:04:16.25" />
                    <SPLIT distance="250" swimtime="00:05:20.03" />
                    <SPLIT distance="300" swimtime="00:06:25.47" />
                    <SPLIT distance="350" swimtime="00:07:16.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="6859" heatid="11590" lane="6" entrytime="00:01:58.00" />
                <RESULT eventid="6738" points="349" reactiontime="+124" swimtime="00:06:53.63" resultid="6860" heatid="11632" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:25.89" />
                    <SPLIT distance="200" swimtime="00:03:18.38" />
                    <SPLIT distance="250" swimtime="00:04:12.00" />
                    <SPLIT distance="300" swimtime="00:05:04.77" />
                    <SPLIT distance="350" swimtime="00:06:00.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMT" nation="POL" clubid="7631" name="Toruń Multisport Team">
          <ATHLETES>
            <ATHLETE firstname="Kamil" lastname="Kordowski" birthdate="1997-10-11" gender="M" nation="POL" swrid="5506630" athleteid="7645">
              <RESULTS>
                <RESULT eventid="6077" points="730" reactiontime="+67" swimtime="00:00:25.36" resultid="7646" heatid="11416" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="6306" points="588" reactiontime="+77" swimtime="00:00:57.96" resultid="7647" heatid="11476" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="610" reactiontime="+73" swimtime="00:00:27.94" resultid="7648" heatid="11539" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="6636" points="552" reactiontime="+76" swimtime="00:01:05.73" resultid="7649" heatid="11593" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Gołembiewski" birthdate="1986-10-28" gender="M" nation="POL" athleteid="7632">
              <RESULTS>
                <RESULT eventid="6111" points="577" reactiontime="+82" swimtime="00:02:32.86" resultid="7633" heatid="11430" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:01:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="673" reactiontime="+82" swimtime="00:02:40.37" resultid="7634" heatid="11459" lane="3" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="557" reactiontime="+84" swimtime="00:01:09.01" resultid="7635" heatid="11494" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="717" reactiontime="+81" swimtime="00:01:10.93" resultid="7636" heatid="11520" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="682" swimtime="00:00:32.78" resultid="7637" heatid="11622" lane="0" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Lietz" birthdate="1952-04-24" gender="M" nation="POL" swrid="4754688" athleteid="7638">
              <RESULTS>
                <RESULT eventid="6077" points="543" swimtime="00:00:34.80" resultid="7639" heatid="11407" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="6169" points="529" swimtime="00:14:10.71" resultid="7640" heatid="11647" lane="9" entrytime="00:14:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:38.14" />
                    <SPLIT distance="150" swimtime="00:02:31.50" />
                    <SPLIT distance="200" swimtime="00:03:24.43" />
                    <SPLIT distance="250" swimtime="00:04:17.07" />
                    <SPLIT distance="300" swimtime="00:05:11.03" />
                    <SPLIT distance="350" swimtime="00:06:06.08" />
                    <SPLIT distance="400" swimtime="00:07:01.49" />
                    <SPLIT distance="450" swimtime="00:07:57.19" />
                    <SPLIT distance="500" swimtime="00:08:51.15" />
                    <SPLIT distance="550" swimtime="00:09:45.63" />
                    <SPLIT distance="600" swimtime="00:10:38.94" />
                    <SPLIT distance="650" swimtime="00:11:32.87" />
                    <SPLIT distance="700" swimtime="00:12:27.53" />
                    <SPLIT distance="750" swimtime="00:13:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="575" reactiontime="+80" swimtime="00:01:17.71" resultid="7641" heatid="11470" lane="8" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="501" reactiontime="+82" swimtime="00:00:40.31" resultid="7642" heatid="11533" lane="0" entrytime="00:00:40.40" />
                <RESULT eventid="6535" points="525" swimtime="00:03:03.44" resultid="7643" heatid="11564" lane="8" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:31.28" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="571" reactiontime="+85" swimtime="00:06:35.10" resultid="7644" heatid="11631" lane="5" entrytime="00:06:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:35.90" />
                    <SPLIT distance="150" swimtime="00:02:27.87" />
                    <SPLIT distance="200" swimtime="00:03:19.65" />
                    <SPLIT distance="250" swimtime="00:04:11.27" />
                    <SPLIT distance="300" swimtime="00:05:01.95" />
                    <SPLIT distance="350" swimtime="00:05:51.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7132" name="Mal Wopr Malbork">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Krauze" birthdate="2001-01-01" gender="F" nation="POL" swrid="4732170" athleteid="7131">
              <RESULTS>
                <RESULT eventid="6059" points="748" swimtime="00:00:28.66" resultid="7133" heatid="11400" lane="4" entrytime="00:00:28.56" entrycourse="SCM" />
                <RESULT eventid="6094" points="659" reactiontime="+76" swimtime="00:02:38.65" resultid="7134" heatid="11420" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="820" reactiontime="+74" swimtime="00:01:01.76" resultid="7135" heatid="11461" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="660" reactiontime="+63" swimtime="00:01:12.57" resultid="7136" heatid="11481" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="704" reactiontime="+65" swimtime="00:00:31.31" resultid="7137" heatid="11528" lane="0" entrytime="00:00:31.21" entrycourse="SCM" />
                <RESULT eventid="6518" points="721" reactiontime="+65" swimtime="00:02:17.32" resultid="7138" heatid="11555" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="628" reactiontime="+69" swimtime="00:01:12.57" resultid="7139" heatid="11586" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="692" reactiontime="+64" swimtime="00:04:50.19" resultid="7140" heatid="11624" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:43.20" />
                    <SPLIT distance="200" swimtime="00:02:20.43" />
                    <SPLIT distance="250" swimtime="00:02:57.62" />
                    <SPLIT distance="300" swimtime="00:03:35.69" />
                    <SPLIT distance="350" swimtime="00:04:13.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7264" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Jankowski" birthdate="1968-01-01" gender="M" nation="POL" athleteid="7263">
              <RESULTS>
                <RESULT eventid="6203" points="413" reactiontime="+126" swimtime="00:22:45.56" resultid="7265" heatid="11653" lane="2" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:03.30" />
                    <SPLIT distance="200" swimtime="00:02:48.70" />
                    <SPLIT distance="250" swimtime="00:03:34.30" />
                    <SPLIT distance="300" swimtime="00:04:21.09" />
                    <SPLIT distance="350" swimtime="00:05:07.41" />
                    <SPLIT distance="400" swimtime="00:05:53.46" />
                    <SPLIT distance="450" swimtime="00:06:39.51" />
                    <SPLIT distance="500" swimtime="00:07:25.72" />
                    <SPLIT distance="550" swimtime="00:08:11.89" />
                    <SPLIT distance="600" swimtime="00:08:57.66" />
                    <SPLIT distance="650" swimtime="00:09:43.58" />
                    <SPLIT distance="700" swimtime="00:10:29.64" />
                    <SPLIT distance="750" swimtime="00:11:15.23" />
                    <SPLIT distance="800" swimtime="00:12:01.60" />
                    <SPLIT distance="850" swimtime="00:12:47.57" />
                    <SPLIT distance="900" swimtime="00:13:33.56" />
                    <SPLIT distance="950" swimtime="00:14:20.58" />
                    <SPLIT distance="1000" swimtime="00:15:06.02" />
                    <SPLIT distance="1050" swimtime="00:15:51.85" />
                    <SPLIT distance="1100" swimtime="00:16:37.94" />
                    <SPLIT distance="1150" swimtime="00:17:24.07" />
                    <SPLIT distance="1200" swimtime="00:18:10.25" />
                    <SPLIT distance="1250" swimtime="00:18:56.32" />
                    <SPLIT distance="1300" swimtime="00:19:43.23" />
                    <SPLIT distance="1350" swimtime="00:20:28.74" />
                    <SPLIT distance="1400" swimtime="00:21:14.94" />
                    <SPLIT distance="1450" swimtime="00:22:01.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00905" nation="POL" region="05" clubid="9222" name="MKS Trójka Łódź">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Szwedzki" birthdate="2000-12-12" gender="M" nation="POL" license="100905700604" swrid="4001538" athleteid="9223">
              <RESULTS>
                <RESULT eventid="6111" points="810" reactiontime="+72" swimtime="00:02:16.19" resultid="9224" heatid="11433" lane="5" entrytime="00:02:15.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="655" reactiontime="+69" swimtime="00:18:24.20" resultid="9225" heatid="11652" lane="4" entrytime="00:16:35.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:44.36" />
                    <SPLIT distance="200" swimtime="00:02:21.29" />
                    <SPLIT distance="250" swimtime="00:02:57.47" />
                    <SPLIT distance="300" swimtime="00:03:34.26" />
                    <SPLIT distance="350" swimtime="00:04:11.17" />
                    <SPLIT distance="400" swimtime="00:04:48.55" />
                    <SPLIT distance="450" swimtime="00:05:25.28" />
                    <SPLIT distance="500" swimtime="00:06:02.17" />
                    <SPLIT distance="550" swimtime="00:06:39.08" />
                    <SPLIT distance="600" swimtime="00:07:16.45" />
                    <SPLIT distance="650" swimtime="00:07:53.67" />
                    <SPLIT distance="700" swimtime="00:08:30.86" />
                    <SPLIT distance="750" swimtime="00:09:07.96" />
                    <SPLIT distance="800" swimtime="00:09:45.69" />
                    <SPLIT distance="850" swimtime="00:10:22.85" />
                    <SPLIT distance="900" swimtime="00:11:00.34" />
                    <SPLIT distance="950" swimtime="00:11:37.72" />
                    <SPLIT distance="1000" swimtime="00:12:13.70" />
                    <SPLIT distance="1050" swimtime="00:12:48.25" />
                    <SPLIT distance="1100" swimtime="00:13:26.31" />
                    <SPLIT distance="1150" swimtime="00:14:03.71" />
                    <SPLIT distance="1200" swimtime="00:14:41.42" />
                    <SPLIT distance="1250" swimtime="00:15:18.93" />
                    <SPLIT distance="1300" swimtime="00:15:56.82" />
                    <SPLIT distance="1350" swimtime="00:16:34.06" />
                    <SPLIT distance="1400" swimtime="00:17:11.25" />
                    <SPLIT distance="1450" swimtime="00:17:48.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="716" reactiontime="+76" swimtime="00:02:33.15" resultid="9226" heatid="11460" lane="6" entrytime="00:02:29.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="662" swimtime="00:02:23.19" resultid="9227" heatid="11504" lane="4" entrytime="00:02:17.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="737" reactiontime="+73" swimtime="00:02:01.77" resultid="9228" heatid="11571" lane="3" entrytime="00:01:58.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="621" reactiontime="+74" swimtime="00:05:14.36" resultid="9229" heatid="11579" lane="5" entrytime="00:04:49.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:56.63" />
                    <SPLIT distance="200" swimtime="00:02:35.56" />
                    <SPLIT distance="250" swimtime="00:03:18.66" />
                    <SPLIT distance="300" swimtime="00:04:01.29" />
                    <SPLIT distance="350" swimtime="00:04:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="528" reactiontime="+71" swimtime="00:02:33.24" resultid="9230" heatid="11606" lane="5" entrytime="00:02:18.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:15.76" />
                    <SPLIT distance="150" swimtime="00:01:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="923" reactiontime="+71" swimtime="00:04:10.08" resultid="9231" heatid="11638" lane="3" entrytime="00:04:12.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:31.54" />
                    <SPLIT distance="200" swimtime="00:02:03.53" />
                    <SPLIT distance="250" swimtime="00:02:35.65" />
                    <SPLIT distance="300" swimtime="00:03:07.99" />
                    <SPLIT distance="350" swimtime="00:03:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="9463" name="UKP Unia Oświęcim">
          <ATHLETES>
            <ATHLETE firstname="Barbara" lastname="Lipniarska-Skubis" birthdate="1952-07-01" gender="F" nation="POL" license="501006600377" athleteid="9464">
              <RESULTS>
                <RESULT eventid="6059" points="219" swimtime="00:00:55.27" resultid="9465" heatid="11395" lane="8" />
                <RESULT eventid="6255" points="346" swimtime="00:05:03.46" resultid="9466" heatid="11451" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.68" />
                    <SPLIT distance="100" swimtime="00:02:25.81" />
                    <SPLIT distance="150" swimtime="00:03:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="200" swimtime="00:02:07.60" resultid="9467" heatid="11462" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="245" reactiontime="+120" swimtime="00:04:27.93" resultid="9468" heatid="11554" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.80" />
                    <SPLIT distance="100" swimtime="00:02:08.66" />
                    <SPLIT distance="150" swimtime="00:03:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="266" swimtime="00:01:07.10" resultid="9469" heatid="11609" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9709" name="KU AZS Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Gralewski" birthdate="1994-01-01" gender="M" nation="POL" swrid="4112460" athleteid="9721">
              <RESULTS>
                <RESULT eventid="6077" points="744" reactiontime="+71" swimtime="00:00:25.20" resultid="9722" heatid="11418" lane="0" entrytime="00:00:24.75" entrycourse="SCM" />
                <RESULT eventid="6111" points="629" swimtime="00:02:20.65" resultid="9723" heatid="11432" lane="9" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:05.75" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="686" reactiontime="+68" swimtime="00:00:55.06" resultid="9724" heatid="11478" lane="0" entrytime="00:00:56.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="668" reactiontime="+69" swimtime="00:00:27.11" resultid="9725" heatid="11539" lane="4" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="6535" points="771" reactiontime="+72" swimtime="00:02:01.19" resultid="9726" heatid="11571" lane="1" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="100" swimtime="00:00:59.07" />
                    <SPLIT distance="150" swimtime="00:01:29.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Mordzonek" birthdate="2001-01-01" gender="M" nation="POL" swrid="5337100" athleteid="9717">
              <RESULTS>
                <RESULT eventid="6374" points="534" reactiontime="+73" swimtime="00:02:33.85" resultid="9718" heatid="11504" lane="8" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="570" reactiontime="+75" swimtime="00:02:12.63" resultid="9719" heatid="11570" lane="9" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="150" swimtime="00:01:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="548" reactiontime="+66" swimtime="00:01:06.35" resultid="9720" heatid="11594" lane="4" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8578" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Grochowski" birthdate="1991-01-01" gender="M" nation="POL" swrid="5464090" athleteid="8577">
              <RESULTS>
                <RESULT eventid="6111" points="381" reactiontime="+83" swimtime="00:02:42.84" resultid="8579" heatid="11425" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="401" reactiontime="+71" swimtime="00:00:35.93" resultid="8580" heatid="11443" lane="8" />
                <RESULT eventid="6340" points="404" reactiontime="+85" swimtime="00:01:14.39" resultid="8581" heatid="11488" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="8582" heatid="11530" lane="7" />
                <RESULT eventid="6535" points="391" reactiontime="+84" swimtime="00:02:25.61" resultid="8583" heatid="11562" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="461" reactiontime="+89" swimtime="00:05:10.80" resultid="8584" heatid="11629" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:51.50" />
                    <SPLIT distance="200" swimtime="00:02:30.77" />
                    <SPLIT distance="250" swimtime="00:03:10.27" />
                    <SPLIT distance="300" swimtime="00:03:50.80" />
                    <SPLIT distance="350" swimtime="00:04:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="8930" name="KS AZS AWF Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Korneliusz" lastname="Zapert" birthdate="2000-04-30" gender="M" nation="POL" license="100201700221" swrid="4621914" athleteid="8949">
              <RESULTS>
                <RESULT eventid="6238" points="729" reactiontime="+61" swimtime="00:00:28.25" resultid="8950" heatid="11450" lane="0" entrytime="00:00:27.59" entrycourse="SCM" />
                <RESULT eventid="6306" points="754" reactiontime="+69" swimtime="00:00:55.58" resultid="8951" heatid="11478" lane="1" entrytime="00:00:55.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="762" reactiontime="+63" swimtime="00:00:26.91" resultid="8952" heatid="11541" lane="5" entrytime="00:00:26.41" entrycourse="SCM" />
                <RESULT eventid="6501" points="727" reactiontime="+54" swimtime="00:01:00.94" resultid="8953" heatid="11553" lane="2" entrytime="00:01:00.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="669" reactiontime="+76" swimtime="00:01:02.08" resultid="8954" heatid="11596" lane="9" entrytime="00:01:02.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="730" reactiontime="+65" swimtime="00:02:17.59" resultid="8955" heatid="11605" lane="1" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="150" swimtime="00:01:42.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" swrid="4236079" athleteid="8931">
              <RESULTS>
                <RESULT eventid="6059" points="782" reactiontime="+69" swimtime="00:00:27.44" resultid="8932" heatid="11401" lane="2" entrytime="00:00:27.16" entrycourse="SCM" />
                <RESULT eventid="6094" points="867" reactiontime="+70" swimtime="00:02:27.84" resultid="8933" heatid="11424" lane="5" entrytime="00:02:33.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="822" reactiontime="+68" swimtime="00:00:59.90" resultid="8934" heatid="11466" lane="5" entrytime="00:00:59.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="847" swimtime="00:01:07.41" resultid="8935" heatid="11486" lane="4" entrytime="00:01:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="829" swimtime="00:00:29.37" resultid="8936" heatid="11528" lane="4" entrytime="00:00:28.78" entrycourse="SCM" />
                <RESULT eventid="6518" points="834" swimtime="00:02:12.80" resultid="8937" heatid="11559" lane="4" entrytime="00:02:09.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:03.18" />
                    <SPLIT distance="150" swimtime="00:01:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="828" swimtime="00:01:04.96" resultid="8938" heatid="11588" lane="4" entrytime="00:01:04.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="803" reactiontime="+75" swimtime="00:04:48.14" resultid="8939" heatid="11628" lane="4" entrytime="00:04:45.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:44.30" />
                    <SPLIT distance="200" swimtime="00:02:21.55" />
                    <SPLIT distance="250" swimtime="00:02:58.72" />
                    <SPLIT distance="300" swimtime="00:03:35.96" />
                    <SPLIT distance="350" swimtime="00:04:12.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Pinkosz" birthdate="1998-04-26" gender="M" nation="POL" license="100201700138" swrid="4368915" athleteid="8940">
              <RESULTS>
                <RESULT eventid="6077" points="856" reactiontime="+62" swimtime="00:00:24.16" resultid="8941" heatid="11418" lane="3" entrytime="00:00:24.17" entrycourse="SCM" />
                <RESULT eventid="6169" points="620" reactiontime="+70" swimtime="00:09:52.18" resultid="8942" heatid="11646" lane="4" entrytime="00:10:25.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:04.56" />
                    <SPLIT distance="150" swimtime="00:01:39.85" />
                    <SPLIT distance="200" swimtime="00:02:15.74" />
                    <SPLIT distance="250" swimtime="00:02:52.14" />
                    <SPLIT distance="300" swimtime="00:03:29.43" />
                    <SPLIT distance="350" swimtime="00:04:06.92" />
                    <SPLIT distance="400" swimtime="00:04:44.81" />
                    <SPLIT distance="450" swimtime="00:05:23.09" />
                    <SPLIT distance="500" swimtime="00:06:01.61" />
                    <SPLIT distance="550" swimtime="00:06:40.30" />
                    <SPLIT distance="600" swimtime="00:07:19.72" />
                    <SPLIT distance="650" swimtime="00:07:58.80" />
                    <SPLIT distance="700" swimtime="00:08:38.33" />
                    <SPLIT distance="750" swimtime="00:09:17.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="878" reactiontime="+65" swimtime="00:00:52.83" resultid="8943" heatid="11479" lane="3" entrytime="00:00:52.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="506" swimtime="00:02:36.60" resultid="8944" heatid="11503" lane="4" entrytime="00:02:46.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="852" reactiontime="+59" swimtime="00:00:25.92" resultid="8945" heatid="11541" lane="6" entrytime="00:00:26.53" entrycourse="SCM" />
                <RESULT eventid="6535" points="710" reactiontime="+68" swimtime="00:02:03.33" resultid="8946" heatid="11571" lane="5" entrytime="00:01:57.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:00:59.74" />
                    <SPLIT distance="150" swimtime="00:01:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="734" reactiontime="+61" swimtime="00:01:00.20" resultid="8947" heatid="11596" lane="0" entrytime="00:01:02.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" status="DNS" swimtime="00:00:00.00" resultid="8948" heatid="11637" lane="4" entrytime="00:04:36.08" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7150" name="Rydułtowska Akademia Aktywnego Seniora 60+">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Lippa" birthdate="1946-01-01" gender="F" nation="POL" swrid="5484413" athleteid="7159">
              <RESULTS>
                <RESULT eventid="6059" points="55" swimtime="00:01:30.91" resultid="7160" heatid="11395" lane="3" entrytime="00:01:28.00" entrycourse="SCM" />
                <RESULT eventid="6220" points="88" swimtime="00:01:37.93" resultid="7161" heatid="11439" lane="9" entrytime="00:01:35.00" entrycourse="SCM" />
                <RESULT eventid="6289" points="68" swimtime="00:03:13.31" resultid="7162" heatid="11462" lane="2" entrytime="00:03:09.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="91" reactiontime="+176" swimtime="00:03:28.04" resultid="7163" heatid="11544" lane="6" entrytime="00:03:26.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="90" swimtime="00:06:41.70" resultid="7164" heatid="11555" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.89" />
                    <SPLIT distance="100" swimtime="00:03:13.64" />
                    <SPLIT distance="150" swimtime="00:04:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="109" reactiontime="+184" swimtime="00:07:03.43" resultid="7165" heatid="11599" lane="9" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:39.64" />
                    <SPLIT distance="100" swimtime="00:03:31.07" />
                    <SPLIT distance="150" swimtime="00:05:17.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="140" swimtime="00:13:07.30" resultid="7166" heatid="11624" lane="4" entrytime="00:13:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.14" />
                    <SPLIT distance="100" swimtime="00:03:08.50" />
                    <SPLIT distance="150" swimtime="00:04:47.99" />
                    <SPLIT distance="200" swimtime="00:06:26.42" />
                    <SPLIT distance="250" swimtime="00:08:09.92" />
                    <SPLIT distance="300" swimtime="00:09:50.44" />
                    <SPLIT distance="350" swimtime="00:11:29.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-01-01" gender="M" nation="POL" swrid="4934027" athleteid="7149">
              <RESULTS>
                <RESULT eventid="6111" points="380" reactiontime="+85" swimtime="00:03:38.90" resultid="7151" heatid="11428" lane="7" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:49.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="420" reactiontime="+84" swimtime="00:26:48.57" resultid="7152" heatid="11653" lane="1" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:38.10" />
                    <SPLIT distance="150" swimtime="00:02:31.46" />
                    <SPLIT distance="200" swimtime="00:03:24.20" />
                    <SPLIT distance="250" swimtime="00:04:17.32" />
                    <SPLIT distance="300" swimtime="00:05:10.61" />
                    <SPLIT distance="350" swimtime="00:06:04.18" />
                    <SPLIT distance="400" swimtime="00:06:57.88" />
                    <SPLIT distance="450" swimtime="00:07:51.12" />
                    <SPLIT distance="500" swimtime="00:08:44.46" />
                    <SPLIT distance="550" swimtime="00:09:38.71" />
                    <SPLIT distance="600" swimtime="00:10:32.94" />
                    <SPLIT distance="650" swimtime="00:11:26.92" />
                    <SPLIT distance="700" swimtime="00:12:20.79" />
                    <SPLIT distance="750" swimtime="00:13:15.15" />
                    <SPLIT distance="800" swimtime="00:14:08.36" />
                    <SPLIT distance="850" swimtime="00:15:03.02" />
                    <SPLIT distance="900" swimtime="00:15:57.05" />
                    <SPLIT distance="950" swimtime="00:16:51.57" />
                    <SPLIT distance="1000" swimtime="00:17:46.34" />
                    <SPLIT distance="1050" swimtime="00:18:41.06" />
                    <SPLIT distance="1100" swimtime="00:19:35.51" />
                    <SPLIT distance="1150" swimtime="00:20:31.66" />
                    <SPLIT distance="1200" swimtime="00:21:26.83" />
                    <SPLIT distance="1250" swimtime="00:22:21.42" />
                    <SPLIT distance="1300" swimtime="00:23:15.61" />
                    <SPLIT distance="1350" swimtime="00:24:10.35" />
                    <SPLIT distance="1400" swimtime="00:25:04.92" />
                    <SPLIT distance="1450" swimtime="00:25:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="525" reactiontime="+88" swimtime="00:00:41.29" resultid="7153" heatid="11446" lane="1" entrytime="00:00:41.72" entrycourse="SCM" />
                <RESULT eventid="6374" points="299" reactiontime="+95" swimtime="00:04:10.25" resultid="7154" heatid="11501" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                    <SPLIT distance="100" swimtime="00:01:58.59" />
                    <SPLIT distance="150" swimtime="00:03:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="441" swimtime="00:00:40.12" resultid="7155" heatid="11532" lane="4" entrytime="00:00:41.21" entrycourse="SCM" />
                <RESULT eventid="6569" points="473" reactiontime="+92" swimtime="00:07:52.43" resultid="7156" heatid="11577" lane="0" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.74" />
                    <SPLIT distance="100" swimtime="00:01:57.70" />
                    <SPLIT distance="150" swimtime="00:02:58.46" />
                    <SPLIT distance="200" swimtime="00:03:57.44" />
                    <SPLIT distance="250" swimtime="00:05:04.69" />
                    <SPLIT distance="300" swimtime="00:06:11.00" />
                    <SPLIT distance="350" swimtime="00:07:02.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="286" swimtime="00:01:48.09" resultid="7157" heatid="11591" lane="9" entrytime="00:01:49.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="429" reactiontime="+99" swimtime="00:03:29.00" resultid="7158" heatid="11603" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:39.92" />
                    <SPLIT distance="150" swimtime="00:02:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8390" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Wilk" birthdate="1990-01-01" gender="M" nation="POL" athleteid="8389">
              <RESULTS>
                <RESULT eventid="6077" points="477" reactiontime="+70" swimtime="00:00:28.31" resultid="8391" heatid="11409" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="6306" points="434" reactiontime="+75" swimtime="00:01:04.74" resultid="8392" heatid="11472" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="427" reactiontime="+75" swimtime="00:00:30.37" resultid="8393" heatid="11536" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="6636" points="360" reactiontime="+76" swimtime="00:01:13.98" resultid="8394" heatid="11592" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8433" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Mańczak" birthdate="1971-01-01" gender="M" nation="POL" swrid="4186188" athleteid="8432">
              <RESULTS>
                <RESULT eventid="6306" points="550" reactiontime="+70" swimtime="00:01:04.78" resultid="8434" heatid="11474" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="516" swimtime="00:02:27.17" resultid="8435" heatid="11566" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="626" reactiontime="+82" swimtime="00:00:31.33" resultid="8436" heatid="11537" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="6374" points="466" reactiontime="+74" swimtime="00:02:59.22" resultid="8437" heatid="11502" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:24.31" />
                    <SPLIT distance="150" swimtime="00:02:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="535" swimtime="00:01:13.49" resultid="8438" heatid="11593" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="8956" name="KS Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" swrid="5398297" athleteid="8957">
              <RESULTS>
                <RESULT eventid="6077" points="622" reactiontime="+77" swimtime="00:00:28.68" resultid="8958" heatid="11402" lane="4" />
                <RESULT eventid="6203" points="451" reactiontime="+101" swimtime="00:22:06.90" resultid="8959" heatid="11654" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                    <SPLIT distance="200" swimtime="00:02:45.81" />
                    <SPLIT distance="250" swimtime="00:03:29.68" />
                    <SPLIT distance="300" swimtime="00:04:13.69" />
                    <SPLIT distance="350" swimtime="00:04:57.91" />
                    <SPLIT distance="400" swimtime="00:05:42.09" />
                    <SPLIT distance="450" swimtime="00:06:25.89" />
                    <SPLIT distance="500" swimtime="00:07:10.17" />
                    <SPLIT distance="550" swimtime="00:07:54.47" />
                    <SPLIT distance="600" swimtime="00:08:39.15" />
                    <SPLIT distance="650" swimtime="00:09:23.80" />
                    <SPLIT distance="700" swimtime="00:10:08.66" />
                    <SPLIT distance="750" swimtime="00:10:53.54" />
                    <SPLIT distance="800" swimtime="00:11:38.70" />
                    <SPLIT distance="850" swimtime="00:12:23.95" />
                    <SPLIT distance="900" swimtime="00:13:09.43" />
                    <SPLIT distance="950" swimtime="00:13:54.69" />
                    <SPLIT distance="1000" swimtime="00:14:39.43" />
                    <SPLIT distance="1050" swimtime="00:15:24.35" />
                    <SPLIT distance="1100" swimtime="00:16:09.11" />
                    <SPLIT distance="1150" swimtime="00:16:53.88" />
                    <SPLIT distance="1200" swimtime="00:17:39.03" />
                    <SPLIT distance="1250" swimtime="00:18:24.34" />
                    <SPLIT distance="1300" swimtime="00:19:09.55" />
                    <SPLIT distance="1350" swimtime="00:19:54.41" />
                    <SPLIT distance="1400" swimtime="00:20:39.41" />
                    <SPLIT distance="1450" swimtime="00:21:24.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="510" reactiontime="+75" swimtime="00:00:35.48" resultid="8960" heatid="11447" lane="1" entrytime="00:00:35.57" entrycourse="SCM" />
                <RESULT eventid="6374" points="488" reactiontime="+94" swimtime="00:02:56.43" resultid="8961" heatid="11500" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="574" swimtime="00:00:32.25" resultid="8962" heatid="11536" lane="8" entrytime="00:00:32.19" entrycourse="SCM" />
                <RESULT eventid="6501" points="468" reactiontime="+75" swimtime="00:01:17.90" resultid="8963" heatid="11550" lane="5" entrytime="00:01:18.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="537" reactiontime="+82" swimtime="00:01:13.37" resultid="8964" heatid="11592" lane="4" entrytime="00:01:15.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="499" reactiontime="+82" swimtime="00:02:55.37" resultid="8965" heatid="11604" lane="6" entrytime="00:02:52.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:24.45" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03210" nation="POL" region="10" clubid="9169" name="MKP Gdańsk">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Gorczyca" birthdate="1990-12-24" gender="M" nation="POL" license="103210700105" swrid="4125944" athleteid="9174">
              <RESULTS>
                <RESULT eventid="6433" points="976" reactiontime="+68" swimtime="00:01:01.83" resultid="9175" heatid="11521" lane="6" entrytime="00:01:04.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="968" reactiontime="+69" swimtime="00:00:28.11" resultid="9176" heatid="11623" lane="2" entrytime="00:00:29.53" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Szczepankiewicz" birthdate="1996-01-29" gender="M" nation="POL" license="103210700110" swrid="4264428" athleteid="9170">
              <RESULTS>
                <RESULT eventid="6340" points="700" reactiontime="+68" swimtime="00:01:02.16" resultid="9171" heatid="11496" lane="2" entrytime="00:01:04.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="764" reactiontime="+72" swimtime="00:01:07.85" resultid="9172" heatid="11521" lane="9" entrytime="00:01:09.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="735" reactiontime="+69" swimtime="00:00:31.31" resultid="9173" heatid="11615" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8621" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Skowroński" birthdate="1975-01-01" gender="M" nation="POL" athleteid="8620">
              <RESULTS>
                <RESULT eventid="6535" points="112" swimtime="00:03:57.95" resultid="8622" heatid="11561" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                    <SPLIT distance="100" swimtime="00:01:57.05" />
                    <SPLIT distance="150" swimtime="00:03:00.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7108" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Alina" lastname="Piekarska" birthdate="1947-01-01" gender="F" nation="POL" athleteid="7107">
              <RESULTS>
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="7109" heatid="11607" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8598" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-01-01" gender="M" nation="POL" swrid="4250678" athleteid="8597">
              <RESULTS>
                <RESULT eventid="6077" points="655" reactiontime="+61" swimtime="00:00:25.47" resultid="8599" heatid="11402" lane="6" />
                <RESULT eventid="6111" points="575" reactiontime="+63" swimtime="00:02:22.02" resultid="8600" heatid="11425" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="656" reactiontime="+72" swimtime="00:00:56.43" resultid="8601" heatid="11467" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="630" reactiontime="+67" swimtime="00:01:04.14" resultid="8602" heatid="11488" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="588" swimtime="00:00:27.29" resultid="8603" heatid="11531" lane="8" />
                <RESULT eventid="6569" points="566" reactiontime="+72" swimtime="00:05:22.71" resultid="8604" heatid="11575" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:50.57" />
                    <SPLIT distance="200" swimtime="00:02:33.27" />
                    <SPLIT distance="250" swimtime="00:03:19.51" />
                    <SPLIT distance="300" swimtime="00:04:05.56" />
                    <SPLIT distance="350" swimtime="00:04:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="628" reactiontime="+76" swimtime="00:01:01.45" resultid="8605" heatid="11589" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="587" reactiontime="+79" swimtime="00:00:33.21" resultid="8606" heatid="11613" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="8865" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Marian" lastname="Lasowy" birthdate="1955-07-15" gender="M" nation="POL" license="502016700001" swrid="4967127" athleteid="8912">
              <RESULTS>
                <RESULT eventid="6203" points="408" reactiontime="+117" swimtime="00:27:04.82" resultid="8913" heatid="11654" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="100" swimtime="00:01:38.81" />
                    <SPLIT distance="150" swimtime="00:02:32.80" />
                    <SPLIT distance="200" swimtime="00:03:26.89" />
                    <SPLIT distance="250" swimtime="00:04:21.12" />
                    <SPLIT distance="300" swimtime="00:05:14.45" />
                    <SPLIT distance="350" swimtime="00:06:09.19" />
                    <SPLIT distance="400" swimtime="00:07:03.50" />
                    <SPLIT distance="450" swimtime="00:07:57.85" />
                    <SPLIT distance="500" swimtime="00:08:52.49" />
                    <SPLIT distance="550" swimtime="00:09:46.53" />
                    <SPLIT distance="600" swimtime="00:10:41.31" />
                    <SPLIT distance="650" swimtime="00:11:35.57" />
                    <SPLIT distance="700" swimtime="00:12:30.43" />
                    <SPLIT distance="750" swimtime="00:13:25.04" />
                    <SPLIT distance="800" swimtime="00:14:20.39" />
                    <SPLIT distance="850" swimtime="00:15:15.09" />
                    <SPLIT distance="900" swimtime="00:16:10.30" />
                    <SPLIT distance="950" swimtime="00:17:05.04" />
                    <SPLIT distance="1000" swimtime="00:17:59.90" />
                    <SPLIT distance="1050" swimtime="00:18:54.68" />
                    <SPLIT distance="1100" swimtime="00:19:50.20" />
                    <SPLIT distance="1150" swimtime="00:20:44.79" />
                    <SPLIT distance="1200" swimtime="00:21:40.15" />
                    <SPLIT distance="1250" swimtime="00:22:35.51" />
                    <SPLIT distance="1300" swimtime="00:23:30.21" />
                    <SPLIT distance="1350" swimtime="00:24:25.08" />
                    <SPLIT distance="1400" swimtime="00:25:20.11" />
                    <SPLIT distance="1450" swimtime="00:26:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="298" reactiontime="+112" swimtime="00:01:31.39" resultid="8914" heatid="11467" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="335" reactiontime="+126" swimtime="00:03:20.69" resultid="8915" heatid="11561" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:37.60" />
                    <SPLIT distance="150" swimtime="00:02:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="375" reactiontime="+96" swimtime="00:07:02.87" resultid="8916" heatid="11630" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="150" swimtime="00:02:33.85" />
                    <SPLIT distance="200" swimtime="00:03:28.11" />
                    <SPLIT distance="250" swimtime="00:04:22.64" />
                    <SPLIT distance="300" swimtime="00:05:17.50" />
                    <SPLIT distance="350" swimtime="00:06:12.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Gudaniec" birthdate="1960-01-01" gender="F" nation="POL" athleteid="9916">
              <RESULTS>
                <RESULT eventid="6094" points="547" reactiontime="+82" swimtime="00:03:33.08" resultid="9917" heatid="11421" lane="4" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                    <SPLIT distance="100" swimtime="00:01:43.79" />
                    <SPLIT distance="150" swimtime="00:02:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="623" swimtime="00:25:14.71" resultid="9918" heatid="11650" lane="7" entrytime="00:24:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:33.83" />
                    <SPLIT distance="150" swimtime="00:02:24.42" />
                    <SPLIT distance="200" swimtime="00:03:15.96" />
                    <SPLIT distance="250" swimtime="00:04:06.33" />
                    <SPLIT distance="300" swimtime="00:04:57.07" />
                    <SPLIT distance="350" swimtime="00:05:47.70" />
                    <SPLIT distance="400" swimtime="00:06:38.40" />
                    <SPLIT distance="450" swimtime="00:07:29.23" />
                    <SPLIT distance="500" swimtime="00:08:19.93" />
                    <SPLIT distance="550" swimtime="00:09:11.23" />
                    <SPLIT distance="600" swimtime="00:10:02.11" />
                    <SPLIT distance="650" swimtime="00:10:52.53" />
                    <SPLIT distance="700" swimtime="00:11:43.07" />
                    <SPLIT distance="750" swimtime="00:12:33.71" />
                    <SPLIT distance="800" swimtime="00:13:24.61" />
                    <SPLIT distance="850" swimtime="00:14:15.23" />
                    <SPLIT distance="900" swimtime="00:15:06.17" />
                    <SPLIT distance="950" swimtime="00:15:56.77" />
                    <SPLIT distance="1000" swimtime="00:16:47.66" />
                    <SPLIT distance="1050" swimtime="00:17:38.60" />
                    <SPLIT distance="1100" swimtime="00:18:29.11" />
                    <SPLIT distance="1150" swimtime="00:19:20.28" />
                    <SPLIT distance="1200" swimtime="00:20:11.18" />
                    <SPLIT distance="1250" swimtime="00:21:01.66" />
                    <SPLIT distance="1300" swimtime="00:21:52.42" />
                    <SPLIT distance="1350" swimtime="00:22:43.39" />
                    <SPLIT distance="1400" swimtime="00:23:34.75" />
                    <SPLIT distance="1450" swimtime="00:24:25.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="437" reactiontime="+83" swimtime="00:00:47.83" resultid="9919" heatid="11439" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="6323" points="498" reactiontime="+78" swimtime="00:01:39.75" resultid="9920" heatid="11483" lane="7" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="486" reactiontime="+80" swimtime="00:01:43.16" resultid="9921" heatid="11545" lane="7" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="615" reactiontime="+83" swimtime="00:07:28.22" resultid="9922" heatid="11573" lane="5" entrytime="00:07:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="100" swimtime="00:01:48.77" />
                    <SPLIT distance="150" swimtime="00:02:45.67" />
                    <SPLIT distance="200" swimtime="00:03:42.16" />
                    <SPLIT distance="250" swimtime="00:04:44.98" />
                    <SPLIT distance="300" swimtime="00:05:48.67" />
                    <SPLIT distance="350" swimtime="00:06:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="531" reactiontime="+79" swimtime="00:03:35.28" resultid="9923" heatid="11599" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                    <SPLIT distance="100" swimtime="00:01:46.31" />
                    <SPLIT distance="150" swimtime="00:02:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="514" swimtime="00:06:33.82" resultid="9924" heatid="11626" lane="0" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="150" swimtime="00:02:22.21" />
                    <SPLIT distance="200" swimtime="00:03:13.13" />
                    <SPLIT distance="250" swimtime="00:04:04.05" />
                    <SPLIT distance="300" swimtime="00:04:55.02" />
                    <SPLIT distance="350" swimtime="00:05:45.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Mamrot" birthdate="1972-12-10" gender="M" nation="POL" license="102016700007" swrid="5471728" athleteid="8883">
              <RESULTS>
                <RESULT eventid="6111" points="382" reactiontime="+74" swimtime="00:03:01.87" resultid="8884" heatid="11429" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6169" points="408" reactiontime="+86" swimtime="00:12:04.92" resultid="8885" heatid="11646" lane="0" entrytime="00:11:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                    <SPLIT distance="200" swimtime="00:02:54.06" />
                    <SPLIT distance="250" swimtime="00:03:40.19" />
                    <SPLIT distance="300" swimtime="00:04:26.51" />
                    <SPLIT distance="350" swimtime="00:05:13.42" />
                    <SPLIT distance="400" swimtime="00:06:00.22" />
                    <SPLIT distance="450" swimtime="00:06:46.46" />
                    <SPLIT distance="500" swimtime="00:07:32.98" />
                    <SPLIT distance="550" swimtime="00:08:19.21" />
                    <SPLIT distance="600" swimtime="00:09:05.98" />
                    <SPLIT distance="650" swimtime="00:09:52.32" />
                    <SPLIT distance="700" swimtime="00:10:38.02" />
                    <SPLIT distance="750" swimtime="00:11:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="478" reactiontime="+77" swimtime="00:03:17.85" resultid="8886" heatid="11457" lane="6" entrytime="00:03:25.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                    <SPLIT distance="150" swimtime="00:02:23.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="417" reactiontime="+78" swimtime="00:01:19.40" resultid="8887" heatid="11491" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="448" swimtime="00:01:27.71" resultid="8888" heatid="11518" lane="9" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="484" reactiontime="+68" swimtime="00:00:39.17" resultid="8889" heatid="11618" lane="6" entrytime="00:00:39.77" entrycourse="SCM" />
                <RESULT eventid="6738" points="456" reactiontime="+75" swimtime="00:05:38.21" resultid="8890" heatid="11633" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:02.03" />
                    <SPLIT distance="200" swimtime="00:02:45.08" />
                    <SPLIT distance="250" swimtime="00:03:29.33" />
                    <SPLIT distance="300" swimtime="00:04:14.06" />
                    <SPLIT distance="350" swimtime="00:04:57.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Winiarczyk" birthdate="1972-01-23" gender="M" nation="POL" license="102016700008" athleteid="8866">
              <RESULTS>
                <RESULT eventid="6077" points="677" reactiontime="+67" swimtime="00:00:27.88" resultid="8867" heatid="11414" lane="0" entrytime="00:00:27.80" />
                <RESULT eventid="6169" points="612" reactiontime="+71" swimtime="00:10:33.17" resultid="8868" heatid="11646" lane="3" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:45.85" />
                    <SPLIT distance="200" swimtime="00:02:25.18" />
                    <SPLIT distance="250" swimtime="00:03:05.14" />
                    <SPLIT distance="300" swimtime="00:03:45.27" />
                    <SPLIT distance="350" swimtime="00:04:25.50" />
                    <SPLIT distance="400" swimtime="00:05:06.04" />
                    <SPLIT distance="450" swimtime="00:05:47.24" />
                    <SPLIT distance="500" swimtime="00:06:28.20" />
                    <SPLIT distance="550" swimtime="00:07:09.38" />
                    <SPLIT distance="600" swimtime="00:07:50.83" />
                    <SPLIT distance="650" swimtime="00:08:32.32" />
                    <SPLIT distance="700" swimtime="00:09:13.67" />
                    <SPLIT distance="750" swimtime="00:09:55.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="572" reactiontime="+71" swimtime="00:00:34.16" resultid="8869" heatid="11447" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="6306" points="669" reactiontime="+69" swimtime="00:01:00.70" resultid="8870" heatid="11475" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="629" reactiontime="+66" swimtime="00:02:17.81" resultid="8871" heatid="11568" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="150" swimtime="00:01:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" status="DNS" swimtime="00:00:00.00" resultid="8872" heatid="11577" lane="4" entrytime="00:06:15.00" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8873" heatid="11604" lane="4" entrytime="00:02:50.00" />
                <RESULT eventid="6738" points="650" reactiontime="+67" swimtime="00:05:00.56" resultid="8874" heatid="11635" lane="3" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:10.79" />
                    <SPLIT distance="150" swimtime="00:01:49.37" />
                    <SPLIT distance="200" swimtime="00:02:28.76" />
                    <SPLIT distance="250" swimtime="00:03:07.83" />
                    <SPLIT distance="300" swimtime="00:03:46.75" />
                    <SPLIT distance="350" swimtime="00:04:26.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Gudaniec" birthdate="1988-01-01" gender="F" nation="POL" athleteid="9925">
              <RESULTS>
                <RESULT eventid="6094" points="542" reactiontime="+86" swimtime="00:02:55.27" resultid="9926" heatid="11423" lane="8" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="599" reactiontime="+89" swimtime="00:11:16.48" resultid="9927" heatid="11643" lane="2" entrytime="00:11:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:39.15" />
                    <SPLIT distance="250" swimtime="00:03:21.61" />
                    <SPLIT distance="300" swimtime="00:04:03.97" />
                    <SPLIT distance="350" swimtime="00:04:47.28" />
                    <SPLIT distance="400" swimtime="00:05:30.87" />
                    <SPLIT distance="450" swimtime="00:06:13.73" />
                    <SPLIT distance="500" swimtime="00:06:57.60" />
                    <SPLIT distance="550" swimtime="00:07:40.30" />
                    <SPLIT distance="600" swimtime="00:08:24.02" />
                    <SPLIT distance="650" swimtime="00:09:07.51" />
                    <SPLIT distance="700" swimtime="00:09:50.74" />
                    <SPLIT distance="750" swimtime="00:10:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="497" reactiontime="+82" swimtime="00:01:21.80" resultid="9928" heatid="11485" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="539" reactiontime="+84" swimtime="00:06:06.76" resultid="9929" heatid="11574" lane="8" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:09.98" />
                    <SPLIT distance="200" swimtime="00:02:56.45" />
                    <SPLIT distance="250" swimtime="00:03:49.00" />
                    <SPLIT distance="300" swimtime="00:04:43.21" />
                    <SPLIT distance="350" swimtime="00:05:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="578" reactiontime="+42" swimtime="00:05:23.49" resultid="9930" heatid="11628" lane="9" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:54.02" />
                    <SPLIT distance="200" swimtime="00:02:35.55" />
                    <SPLIT distance="250" swimtime="00:03:17.57" />
                    <SPLIT distance="300" swimtime="00:03:59.94" />
                    <SPLIT distance="350" swimtime="00:04:42.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kielar" birthdate="1974-01-21" gender="M" nation="POL" license="102016700020" swrid="4992896" athleteid="8891">
              <RESULTS>
                <RESULT eventid="6111" points="669" reactiontime="+85" swimtime="00:02:31.32" resultid="8892" heatid="11431" lane="5" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:09.61" />
                    <SPLIT distance="150" swimtime="00:01:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="697" reactiontime="+76" swimtime="00:01:07.64" resultid="8893" heatid="11488" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="518" reactiontime="+89" swimtime="00:02:43.92" resultid="8894" heatid="11504" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:54.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="726" reactiontime="+70" swimtime="00:00:28.57" resultid="8895" heatid="11540" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="6636" points="748" reactiontime="+71" swimtime="00:01:04.49" resultid="8896" heatid="11594" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="708" reactiontime="+76" swimtime="00:00:33.97" resultid="8897" heatid="11620" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Kijanka" birthdate="1982-08-02" gender="F" nation="POL" license="102016600021" athleteid="8875">
              <RESULTS>
                <RESULT eventid="6094" points="459" reactiontime="+76" swimtime="00:03:10.17" resultid="8876" heatid="11422" lane="3" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="447" reactiontime="+80" swimtime="00:12:31.88" resultid="8877" heatid="11644" lane="4" entrytime="00:12:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                    <SPLIT distance="150" swimtime="00:02:13.65" />
                    <SPLIT distance="200" swimtime="00:03:01.69" />
                    <SPLIT distance="250" swimtime="00:03:49.58" />
                    <SPLIT distance="300" swimtime="00:04:37.59" />
                    <SPLIT distance="350" swimtime="00:05:25.55" />
                    <SPLIT distance="400" swimtime="00:06:13.45" />
                    <SPLIT distance="450" swimtime="00:07:00.96" />
                    <SPLIT distance="500" swimtime="00:07:48.51" />
                    <SPLIT distance="550" swimtime="00:08:35.94" />
                    <SPLIT distance="600" swimtime="00:09:23.19" />
                    <SPLIT distance="650" swimtime="00:10:10.65" />
                    <SPLIT distance="700" swimtime="00:10:58.45" />
                    <SPLIT distance="750" swimtime="00:11:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="554" swimtime="00:03:22.25" resultid="8878" heatid="11454" lane="9" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" status="DNS" swimtime="00:00:00.00" resultid="8879" heatid="11483" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="6552" points="492" swimtime="00:06:43.04" resultid="8880" heatid="11574" lane="1" entrytime="00:06:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:34.60" />
                    <SPLIT distance="150" swimtime="00:02:29.96" />
                    <SPLIT distance="200" swimtime="00:03:21.89" />
                    <SPLIT distance="250" swimtime="00:04:17.06" />
                    <SPLIT distance="300" swimtime="00:05:12.03" />
                    <SPLIT distance="350" swimtime="00:05:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="392" reactiontime="+70" swimtime="00:01:28.26" resultid="8881" heatid="11587" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="444" reactiontime="+73" swimtime="00:06:02.93" resultid="8882" heatid="11626" lane="2" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                    <SPLIT distance="150" swimtime="00:02:10.12" />
                    <SPLIT distance="200" swimtime="00:02:57.04" />
                    <SPLIT distance="250" swimtime="00:03:44.16" />
                    <SPLIT distance="300" swimtime="00:04:30.54" />
                    <SPLIT distance="350" swimtime="00:05:17.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kruk" birthdate="1982-01-18" gender="M" nation="POL" license="102016700024" swrid="5506631" athleteid="8898">
              <RESULTS>
                <RESULT eventid="6111" points="391" reactiontime="+91" swimtime="00:02:54.79" resultid="8899" heatid="11430" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                    <SPLIT distance="150" swimtime="00:02:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="431" reactiontime="+86" swimtime="00:21:58.94" resultid="8900" heatid="11653" lane="4" entrytime="00:22:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                    <SPLIT distance="200" swimtime="00:02:37.41" />
                    <SPLIT distance="250" swimtime="00:03:20.73" />
                    <SPLIT distance="300" swimtime="00:04:04.17" />
                    <SPLIT distance="350" swimtime="00:04:47.92" />
                    <SPLIT distance="400" swimtime="00:05:31.91" />
                    <SPLIT distance="450" swimtime="00:06:16.38" />
                    <SPLIT distance="500" swimtime="00:07:01.20" />
                    <SPLIT distance="550" swimtime="00:07:46.09" />
                    <SPLIT distance="600" swimtime="00:08:31.11" />
                    <SPLIT distance="650" swimtime="00:09:16.49" />
                    <SPLIT distance="700" swimtime="00:10:02.02" />
                    <SPLIT distance="750" swimtime="00:10:47.65" />
                    <SPLIT distance="800" swimtime="00:11:32.83" />
                    <SPLIT distance="850" swimtime="00:12:17.63" />
                    <SPLIT distance="900" swimtime="00:13:03.06" />
                    <SPLIT distance="950" swimtime="00:13:48.70" />
                    <SPLIT distance="1000" swimtime="00:14:33.26" />
                    <SPLIT distance="1050" swimtime="00:15:17.74" />
                    <SPLIT distance="1100" swimtime="00:16:02.22" />
                    <SPLIT distance="1150" swimtime="00:16:47.62" />
                    <SPLIT distance="1200" swimtime="00:17:32.81" />
                    <SPLIT distance="1250" swimtime="00:18:17.78" />
                    <SPLIT distance="1300" swimtime="00:19:03.22" />
                    <SPLIT distance="1350" swimtime="00:19:48.23" />
                    <SPLIT distance="1400" swimtime="00:20:33.24" />
                    <SPLIT distance="1450" swimtime="00:21:17.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="469" reactiontime="+81" swimtime="00:01:05.96" resultid="8901" heatid="11473" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="436" reactiontime="+77" swimtime="00:01:18.86" resultid="8902" heatid="11491" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="419" reactiontime="+81" swimtime="00:00:33.58" resultid="8903" heatid="11535" lane="9" entrytime="00:00:34.13" entrycourse="SCM" />
                <RESULT eventid="6535" points="452" reactiontime="+86" swimtime="00:02:27.24" resultid="8904" heatid="11567" lane="2" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:48.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="393" reactiontime="+95" swimtime="00:05:28.37" resultid="8905" heatid="11633" lane="5" entrytime="00:05:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                    <SPLIT distance="200" swimtime="00:02:40.41" />
                    <SPLIT distance="250" swimtime="00:03:23.38" />
                    <SPLIT distance="300" swimtime="00:04:06.11" />
                    <SPLIT distance="350" swimtime="00:04:48.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Ćwikła" birthdate="1974-08-22" gender="M" nation="POL" license="102016700002" swrid="5506628" athleteid="8906">
              <RESULTS>
                <RESULT eventid="6169" points="504" reactiontime="+90" swimtime="00:10:52.88" resultid="8907" heatid="11646" lane="6" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                    <SPLIT distance="200" swimtime="00:02:36.12" />
                    <SPLIT distance="250" swimtime="00:03:16.86" />
                    <SPLIT distance="300" swimtime="00:03:57.51" />
                    <SPLIT distance="350" swimtime="00:04:38.72" />
                    <SPLIT distance="400" swimtime="00:05:19.73" />
                    <SPLIT distance="450" swimtime="00:06:01.34" />
                    <SPLIT distance="500" swimtime="00:06:43.43" />
                    <SPLIT distance="550" swimtime="00:07:25.55" />
                    <SPLIT distance="600" swimtime="00:08:08.03" />
                    <SPLIT distance="650" swimtime="00:08:50.14" />
                    <SPLIT distance="700" swimtime="00:09:31.97" />
                    <SPLIT distance="750" swimtime="00:10:13.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="548" reactiontime="+73" swimtime="00:00:34.05" resultid="8908" heatid="11448" lane="8" entrytime="00:00:33.92" entrycourse="SCM" />
                <RESULT eventid="6501" points="502" reactiontime="+81" swimtime="00:01:14.74" resultid="8909" heatid="11551" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="469" reactiontime="+83" swimtime="00:06:11.92" resultid="8910" heatid="11578" lane="1" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                    <SPLIT distance="150" swimtime="00:02:12.63" />
                    <SPLIT distance="200" swimtime="00:02:58.84" />
                    <SPLIT distance="250" swimtime="00:03:54.98" />
                    <SPLIT distance="300" swimtime="00:04:50.05" />
                    <SPLIT distance="350" swimtime="00:05:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="378" reactiontime="+70" swimtime="00:03:01.87" resultid="8911" heatid="11605" lane="8" entrytime="00:02:44.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:29.28" />
                    <SPLIT distance="150" swimtime="00:02:17.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Wróblewski" birthdate="1990-01-01" gender="M" nation="POL" athleteid="9938">
              <RESULTS>
                <RESULT eventid="6467" points="680" reactiontime="+65" swimtime="00:00:26.00" resultid="9939" heatid="11541" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="6636" points="766" reactiontime="+70" swimtime="00:00:57.50" resultid="9940" heatid="11596" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="723" reactiontime="+72" swimtime="00:04:27.59" resultid="9941" heatid="11636" lane="1" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="150" swimtime="00:01:38.93" />
                    <SPLIT distance="200" swimtime="00:02:12.94" />
                    <SPLIT distance="250" swimtime="00:02:47.05" />
                    <SPLIT distance="300" swimtime="00:03:21.49" />
                    <SPLIT distance="350" swimtime="00:03:55.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Wejnerowska" birthdate="1993-01-01" gender="F" nation="POL" athleteid="9931">
              <RESULTS>
                <RESULT eventid="6059" points="403" swimtime="00:00:34.22" resultid="9932" heatid="11397" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="6094" points="391" swimtime="00:03:12.68" resultid="9933" heatid="11422" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:34.73" />
                    <SPLIT distance="150" swimtime="00:02:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="420" swimtime="00:03:25.15" resultid="9934" heatid="11453" lane="4" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:40.39" />
                    <SPLIT distance="150" swimtime="00:02:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" status="DNS" swimtime="00:00:00.00" resultid="9935" heatid="11556" lane="8" entrytime="00:02:54.00" />
                <RESULT eventid="6552" points="411" reactiontime="+85" swimtime="00:06:43.61" resultid="9936" heatid="11573" lane="4" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:41.47" />
                    <SPLIT distance="150" swimtime="00:02:34.63" />
                    <SPLIT distance="200" swimtime="00:03:26.28" />
                    <SPLIT distance="250" swimtime="00:04:21.50" />
                    <SPLIT distance="300" swimtime="00:05:15.60" />
                    <SPLIT distance="350" swimtime="00:06:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="420" swimtime="00:05:57.60" resultid="9937" heatid="11626" lane="3" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:10.15" />
                    <SPLIT distance="200" swimtime="00:02:57.08" />
                    <SPLIT distance="250" swimtime="00:03:43.77" />
                    <SPLIT distance="300" swimtime="00:04:29.77" />
                    <SPLIT distance="350" swimtime="00:05:15.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+85" swimtime="00:01:47.43" resultid="8918" heatid="11584" lane="7" entrytime="00:01:49.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                    <SPLIT distance="100" swimtime="00:00:55.95" />
                    <SPLIT distance="150" swimtime="00:01:23.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8891" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="8906" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="8866" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="9938" number="4" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" reactiontime="+76" swimtime="00:02:00.51" resultid="8919" heatid="12332" lane="7" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:32.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8906" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="8891" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="9938" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="8866" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6391" reactiontime="+79" swimtime="00:02:29.80" resultid="8917" heatid="11507" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:32.23" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8875" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="9916" number="2" />
                    <RELAYPOSITION athleteid="8891" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="8866" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="9484" name="UKS ,,Trójka&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="9485">
              <RESULTS>
                <RESULT eventid="6374" points="685" reactiontime="+89" swimtime="00:02:29.29" resultid="9486" heatid="11504" lane="2" entrytime="00:02:32.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="644" reactiontime="+89" swimtime="00:05:34.69" resultid="9487" heatid="11576" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:59.78" />
                    <SPLIT distance="200" swimtime="00:02:44.84" />
                    <SPLIT distance="250" swimtime="00:03:31.14" />
                    <SPLIT distance="300" swimtime="00:04:17.52" />
                    <SPLIT distance="350" swimtime="00:04:56.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="644" reactiontime="+95" swimtime="00:01:07.78" resultid="9488" heatid="11589" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8628" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Klimkowski" birthdate="1981-01-01" gender="M" nation="POL" swrid="4629756" athleteid="8627">
              <RESULTS>
                <RESULT eventid="6077" points="14" swimtime="00:01:36.22" resultid="8629" heatid="11404" lane="1" entrytime="00:01:35.59" />
                <RESULT eventid="6238" points="23" swimtime="00:01:34.48" resultid="8630" heatid="11444" lane="0" entrytime="00:01:37.98" />
                <RESULT eventid="6306" points="14" swimtime="00:03:30.65" resultid="8631" heatid="11467" lane="3" entrytime="00:03:11.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="33" swimtime="00:03:02.64" resultid="8632" heatid="11547" lane="0" entrytime="00:03:11.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="16" swimtime="00:07:27.90" resultid="8633" heatid="11560" lane="0" entrytime="00:07:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:42.88" />
                    <SPLIT distance="100" swimtime="00:03:37.12" />
                    <SPLIT distance="150" swimtime="00:05:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="40" swimtime="00:06:18.86" resultid="8634" heatid="11602" lane="8" entrytime="00:06:41.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.89" />
                    <SPLIT distance="100" swimtime="00:03:06.59" />
                    <SPLIT distance="150" swimtime="00:04:46.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="16" swimtime="00:15:51.34" resultid="8635" heatid="11630" lane="2" entrytime="00:14:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.98" />
                    <SPLIT distance="100" swimtime="00:03:48.28" />
                    <SPLIT distance="150" swimtime="00:05:48.15" />
                    <SPLIT distance="200" swimtime="00:07:51.26" />
                    <SPLIT distance="250" swimtime="00:09:51.87" />
                    <SPLIT distance="300" swimtime="00:11:52.64" />
                    <SPLIT distance="350" swimtime="00:13:54.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6942" name="RMKS Rybnik">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" swrid="4992966" athleteid="6943">
              <RESULTS>
                <RESULT eventid="6059" points="760" reactiontime="+77" swimtime="00:00:28.79" resultid="6944" heatid="11401" lane="8" entrytime="00:00:28.20" />
                <RESULT eventid="6094" points="727" swimtime="00:02:43.25" resultid="6945" heatid="11424" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="150" swimtime="00:02:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6289" points="761" swimtime="00:01:04.05" resultid="6946" heatid="11466" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="776" reactiontime="+68" swimtime="00:01:14.13" resultid="6947" heatid="11486" lane="0" entrytime="00:01:13.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="864" reactiontime="+71" swimtime="00:00:30.76" resultid="6948" heatid="11528" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7111" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Rusakiewicz" birthdate="1979-01-01" gender="F" nation="POL" swrid="4050389" athleteid="7110">
              <RESULTS>
                <RESULT eventid="6094" points="776" reactiontime="+83" swimtime="00:02:39.72" resultid="7112" heatid="11420" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:13.78" />
                    <SPLIT distance="150" swimtime="00:02:00.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="634" reactiontime="+80" swimtime="00:02:51.86" resultid="7113" heatid="11498" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="733" reactiontime="+80" swimtime="00:02:23.38" resultid="7114" heatid="11555" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:47.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="113/14" nation="POL" clubid="8347" name="Fundacja HASTEN">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="Bochyńska" birthdate="1990-06-10" gender="F" nation="POL" license="511314600001" swrid="4061587" athleteid="8352" />
            <ATHLETE firstname="Marta" lastname="Piasecka" birthdate="1991-07-19" gender="F" nation="POL" swrid="4072336" athleteid="8357">
              <RESULTS>
                <RESULT eventid="6094" points="806" reactiontime="+92" swimtime="00:02:33.53" resultid="8358" heatid="11424" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="674" reactiontime="+79" swimtime="00:05:40.63" resultid="8359" heatid="11574" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:59.21" />
                    <SPLIT distance="200" swimtime="00:02:40.71" />
                    <SPLIT distance="250" swimtime="00:03:29.36" />
                    <SPLIT distance="300" swimtime="00:04:19.52" />
                    <SPLIT distance="350" swimtime="00:05:00.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Karpińska" birthdate="1991-07-26" gender="F" nation="POL" athleteid="8353">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6186" points="810" reactiontime="+77" swimtime="00:19:42.50" resultid="8354" heatid="11650" lane="4" entrytime="00:19:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:51.80" />
                    <SPLIT distance="200" swimtime="00:02:31.02" />
                    <SPLIT distance="250" swimtime="00:03:10.12" />
                    <SPLIT distance="300" swimtime="00:03:49.24" />
                    <SPLIT distance="350" swimtime="00:04:28.15" />
                    <SPLIT distance="400" swimtime="00:05:07.06" />
                    <SPLIT distance="450" swimtime="00:05:45.55" />
                    <SPLIT distance="500" swimtime="00:06:24.16" />
                    <SPLIT distance="550" swimtime="00:07:02.27" />
                    <SPLIT distance="600" swimtime="00:07:40.61" />
                    <SPLIT distance="650" swimtime="00:08:19.33" />
                    <SPLIT distance="700" swimtime="00:08:57.76" />
                    <SPLIT distance="750" swimtime="00:09:36.08" />
                    <SPLIT distance="800" swimtime="00:10:13.79" />
                    <SPLIT distance="850" swimtime="00:10:54.41" />
                    <SPLIT distance="900" swimtime="00:11:35.70" />
                    <SPLIT distance="950" swimtime="00:12:16.96" />
                    <SPLIT distance="1000" swimtime="00:12:57.71" />
                    <SPLIT distance="1050" swimtime="00:13:38.54" />
                    <SPLIT distance="1100" swimtime="00:14:19.16" />
                    <SPLIT distance="1150" swimtime="00:15:00.01" />
                    <SPLIT distance="1200" swimtime="00:15:41.35" />
                    <SPLIT distance="1250" swimtime="00:16:22.07" />
                    <SPLIT distance="1300" swimtime="00:17:02.80" />
                    <SPLIT distance="1350" swimtime="00:17:43.28" />
                    <SPLIT distance="1400" swimtime="00:18:23.70" />
                    <SPLIT distance="1450" swimtime="00:19:03.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="610" reactiontime="+78" swimtime="00:02:48.28" resultid="8355" heatid="11499" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:57.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="770" reactiontime="+77" swimtime="00:00:30.75" resultid="8356" heatid="11528" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Pawlaczek" birthdate="1993-01-04" gender="F" nation="POL" license="111314600002" swrid="4072670" athleteid="8348">
              <RESULTS>
                <RESULT eventid="6059" points="795" reactiontime="+76" swimtime="00:00:27.30" resultid="8349" heatid="11401" lane="3" entrytime="00:00:26.99" />
                <RESULT eventid="6323" points="828" reactiontime="+78" swimtime="00:01:07.92" resultid="8350" heatid="11486" lane="5" entrytime="00:01:08.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="847" reactiontime="+76" swimtime="00:00:29.16" resultid="8351" heatid="11528" lane="5" entrytime="00:00:29.29" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6586" reactiontime="+78" swimtime="00:01:52.96" resultid="8360" heatid="11581" lane="4" entrytime="00:01:58.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                    <SPLIT distance="100" swimtime="00:00:55.20" />
                    <SPLIT distance="150" swimtime="00:01:25.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8348" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="8357" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="8352" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="8353" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6886" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tobiasz" lastname="Jankowski" birthdate="1983-01-01" gender="M" nation="POL" athleteid="6885">
              <RESULTS>
                <RESULT eventid="6340" points="367" reactiontime="+73" swimtime="00:01:19.31" resultid="6887" heatid="11487" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="6888" heatid="11513" lane="4" />
                <RESULT eventid="6467" points="386" reactiontime="+76" swimtime="00:00:32.45" resultid="6889" heatid="11529" lane="5" />
                <RESULT eventid="6704" points="518" reactiontime="+85" swimtime="00:00:35.92" resultid="6890" heatid="11614" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7168" name="niezrzeszona Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Bołtuć" birthdate="1983-01-01" gender="F" nation="POL" athleteid="7167">
              <RESULTS>
                <RESULT eventid="6186" points="529" swimtime="00:22:41.62" resultid="7169" heatid="11650" lane="2" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                    <SPLIT distance="150" swimtime="00:02:10.26" />
                    <SPLIT distance="200" swimtime="00:02:55.99" />
                    <SPLIT distance="250" swimtime="00:03:41.80" />
                    <SPLIT distance="300" swimtime="00:04:27.26" />
                    <SPLIT distance="350" swimtime="00:05:12.39" />
                    <SPLIT distance="400" swimtime="00:05:57.53" />
                    <SPLIT distance="450" swimtime="00:06:43.00" />
                    <SPLIT distance="500" swimtime="00:07:28.42" />
                    <SPLIT distance="550" swimtime="00:08:13.77" />
                    <SPLIT distance="600" swimtime="00:08:59.23" />
                    <SPLIT distance="650" swimtime="00:09:45.07" />
                    <SPLIT distance="700" swimtime="00:10:31.47" />
                    <SPLIT distance="750" swimtime="00:11:17.41" />
                    <SPLIT distance="800" swimtime="00:12:02.45" />
                    <SPLIT distance="850" swimtime="00:12:47.47" />
                    <SPLIT distance="900" swimtime="00:13:33.44" />
                    <SPLIT distance="950" swimtime="00:14:19.45" />
                    <SPLIT distance="1000" swimtime="00:15:05.84" />
                    <SPLIT distance="1050" swimtime="00:15:52.20" />
                    <SPLIT distance="1100" swimtime="00:16:38.22" />
                    <SPLIT distance="1150" swimtime="00:17:23.71" />
                    <SPLIT distance="1200" swimtime="00:18:09.62" />
                    <SPLIT distance="1250" swimtime="00:18:55.34" />
                    <SPLIT distance="1300" swimtime="00:19:41.38" />
                    <SPLIT distance="1350" swimtime="00:20:27.04" />
                    <SPLIT distance="1400" swimtime="00:21:12.81" />
                    <SPLIT distance="1450" swimtime="00:21:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6289" points="396" reactiontime="+102" swimtime="00:01:18.68" resultid="7170" heatid="11463" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="451" reactiontime="+106" swimtime="00:02:46.99" resultid="7171" heatid="11558" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:02:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="472" reactiontime="+105" swimtime="00:05:50.61" resultid="7172" heatid="11627" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:08.26" />
                    <SPLIT distance="200" swimtime="00:02:53.21" />
                    <SPLIT distance="250" swimtime="00:03:38.16" />
                    <SPLIT distance="300" swimtime="00:04:23.39" />
                    <SPLIT distance="350" swimtime="00:05:08.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="273" reactiontime="+107" swimtime="00:01:38.28" resultid="7173" heatid="11586" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="408" reactiontime="+116" swimtime="00:07:05.31" resultid="7174" heatid="11574" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.17" />
                    <SPLIT distance="100" swimtime="00:01:43.47" />
                    <SPLIT distance="150" swimtime="00:02:39.39" />
                    <SPLIT distance="200" swimtime="00:03:34.60" />
                    <SPLIT distance="250" swimtime="00:04:32.52" />
                    <SPLIT distance="300" swimtime="00:05:31.47" />
                    <SPLIT distance="350" swimtime="00:06:19.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7985" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="8858">
              <RESULTS>
                <RESULT eventid="6272" points="452" swimtime="00:03:30.97" resultid="8859" heatid="11457" lane="1" entrytime="00:03:27.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:40.30" />
                    <SPLIT distance="150" swimtime="00:02:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="221" swimtime="00:03:49.61" resultid="8860" heatid="11501" lane="4" entrytime="00:03:53.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:43.93" />
                    <SPLIT distance="150" swimtime="00:02:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="289" reactiontime="+124" swimtime="00:00:42.40" resultid="8861" heatid="11533" lane="9" entrytime="00:00:40.86" entrycourse="SCM" />
                <RESULT eventid="6569" points="285" reactiontime="+114" swimtime="00:07:41.44" resultid="8862" heatid="11576" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:47.54" />
                    <SPLIT distance="150" swimtime="00:02:52.33" />
                    <SPLIT distance="200" swimtime="00:04:02.07" />
                    <SPLIT distance="250" swimtime="00:04:59.79" />
                    <SPLIT distance="300" swimtime="00:05:57.41" />
                    <SPLIT distance="350" swimtime="00:06:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="266" swimtime="00:01:38.00" resultid="8863" heatid="11591" lane="6" entrytime="00:01:37.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="340" reactiontime="+120" swimtime="00:00:43.67" resultid="8864" heatid="11617" lane="1" entrytime="00:00:43.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Ostapczuk" birthdate="1970-07-13" gender="M" nation="POL" athleteid="8001">
              <RESULTS>
                <RESULT eventid="6272" points="388" reactiontime="+92" swimtime="00:03:32.08" resultid="8002" heatid="11457" lane="0" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:39.92" />
                    <SPLIT distance="150" swimtime="00:02:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="271" reactiontime="+100" swimtime="00:01:31.66" resultid="8003" heatid="11490" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="330" reactiontime="+103" swimtime="00:01:37.16" resultid="8004" heatid="11517" lane="7" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Matusiewicz" birthdate="1998-04-12" gender="M" nation="POL" swrid="5058424" athleteid="7986">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="7987" heatid="11405" lane="1" entrytime="00:00:40.74" />
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7988" heatid="11428" lane="9" entrytime="00:03:44.00" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="7989" heatid="11445" lane="1" entrytime="00:00:45.12" />
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="7990" heatid="11489" lane="3" entrytime="00:01:40.10" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="7991" heatid="11532" lane="1" entrytime="00:00:46.46" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="7992" heatid="11549" lane="6" entrytime="00:01:40.40" />
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="7993" heatid="11591" lane="0" entrytime="00:01:49.78" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7994" heatid="11616" lane="0" entrytime="00:00:51.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Bystry" birthdate="1977-03-14" gender="M" nation="POL" swrid="4754758" athleteid="7995">
              <RESULTS>
                <RESULT eventid="6077" points="599" swimtime="00:00:28.31" resultid="7996" heatid="11413" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="6306" points="605" reactiontime="+76" swimtime="00:01:02.56" resultid="7997" heatid="11476" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="525" reactiontime="+76" swimtime="00:01:14.35" resultid="7998" heatid="11493" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="583" reactiontime="+72" swimtime="00:00:30.74" resultid="7999" heatid="11537" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="8000" heatid="11621" lane="9" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Safrończyk" birthdate="1988-05-30" gender="M" nation="POL" license="510414700001" swrid="4072743" athleteid="8853">
              <RESULTS>
                <RESULT eventid="6272" points="921" swimtime="00:02:24.39" resultid="8854" heatid="11460" lane="4" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="781" reactiontime="+64" swimtime="00:00:59.72" resultid="8855" heatid="11497" lane="3" entrytime="00:00:57.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="816" reactiontime="+64" swimtime="00:01:05.64" resultid="8856" heatid="11521" lane="4" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="845" swimtime="00:00:29.41" resultid="8857" heatid="11623" lane="4" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="8847">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="6077" reactiontime="+66" status="DSQ" swimtime="00:00:00.00" resultid="8848" heatid="11405" lane="2" entrytime="00:00:39.56" entrycourse="SCM" />
                <RESULT eventid="6238" points="237" reactiontime="+80" swimtime="00:00:47.37" resultid="8849" heatid="11444" lane="4" entrytime="00:00:47.88" entrycourse="SCM" />
                <RESULT eventid="6306" points="282" swimtime="00:01:28.39" resultid="8850" heatid="11468" lane="4" entrytime="00:01:37.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="247" reactiontime="+108" swimtime="00:03:21.70" resultid="8851" heatid="11563" lane="1" entrytime="00:03:44.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="100" swimtime="00:01:35.00" />
                    <SPLIT distance="150" swimtime="00:02:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="264" reactiontime="+76" swimtime="00:03:43.01" resultid="8852" heatid="11603" lane="9" entrytime="00:03:53.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                    <SPLIT distance="100" swimtime="00:01:47.86" />
                    <SPLIT distance="150" swimtime="00:02:46.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+193" swimtime="00:02:03.06" resultid="8006" heatid="11583" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="100" swimtime="00:00:51.81" />
                    <SPLIT distance="150" swimtime="00:01:26.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7995" number="1" reactiontime="+193" />
                    <RELAYPOSITION athleteid="8853" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="8001" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="8847" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00612" nation="POL" region="12" clubid="8966" name="KS KSZO Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Sejmicki" birthdate="1961-05-04" gender="M" nation="POL" license="500612700426" swrid="5558380" athleteid="8973">
              <RESULTS>
                <RESULT eventid="6077" points="401" reactiontime="+103" swimtime="00:00:36.38" resultid="8974" heatid="11406" lane="8" entrytime="00:00:36.78" entrycourse="SCM" />
                <RESULT eventid="6272" points="402" reactiontime="+111" swimtime="00:03:44.76" resultid="8975" heatid="11456" lane="2" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:45.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="432" reactiontime="+111" swimtime="00:01:37.69" resultid="8976" heatid="11516" lane="5" entrytime="00:01:41.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="402" reactiontime="+192" swimtime="00:00:44.35" resultid="8977" heatid="11617" lane="0" entrytime="00:00:44.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Żak" birthdate="1959-11-22" gender="M" nation="POL" license="500612700512" swrid="5558381" athleteid="8978">
              <RESULTS>
                <RESULT eventid="6077" points="434" swimtime="00:00:35.45" resultid="8979" heatid="11406" lane="1" entrytime="00:00:36.37" entrycourse="SCM" />
                <RESULT eventid="6238" points="315" reactiontime="+86" swimtime="00:00:46.14" resultid="8980" heatid="11445" lane="9" entrytime="00:00:47.70" entrycourse="SCM" />
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="8981" heatid="11489" lane="6" entrytime="00:01:45.81" entrycourse="SCM" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="8982" heatid="11549" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8983" heatid="11602" lane="3" entrytime="00:04:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Orłowski" birthdate="1960-02-26" gender="M" nation="POL" license="500612700404" athleteid="8967">
              <RESULTS>
                <RESULT eventid="6077" points="314" reactiontime="+73" swimtime="00:00:39.45" resultid="8968" heatid="11406" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="6238" points="209" reactiontime="+82" swimtime="00:00:52.86" resultid="8969" heatid="11445" lane="6" entrytime="00:00:44.00" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="8970" heatid="11469" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="6433" status="DNS" swimtime="00:00:00.00" resultid="8971" heatid="11516" lane="2" entrytime="00:01:43.00" />
                <RESULT eventid="6704" points="270" reactiontime="+93" swimtime="00:00:50.65" resultid="8972" heatid="11617" lane="8" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GBR" clubid="11380" name="Wantage White Horses">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Rybak" birthdate="1980-01-01" gender="M" nation="POL" athleteid="11379">
              <RESULTS>
                <RESULT eventid="6077" points="652" reactiontime="+76" swimtime="00:00:26.76" resultid="11381" heatid="11415" lane="2" entrytime="00:00:26.80" />
                <RESULT eventid="6111" points="555" reactiontime="+88" swimtime="00:02:35.54" resultid="11382" heatid="11431" lane="9" entrytime="00:02:42.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:58.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="665" reactiontime="+80" swimtime="00:01:08.51" resultid="11383" heatid="11492" lane="7" entrytime="00:01:17.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="677" reactiontime="+75" swimtime="00:00:28.62" resultid="11384" heatid="11539" lane="2" entrytime="00:00:28.90" />
                <RESULT eventid="6636" points="656" reactiontime="+78" swimtime="00:01:05.16" resultid="11385" heatid="11595" lane="2" entrytime="00:01:04.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GS&amp;R" nation="POL" clubid="8607" name="Garmin Swimming and Rescue">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Orłowski" birthdate="1982-12-11" gender="M" nation="POL" athleteid="8609">
              <RESULTS>
                <RESULT eventid="6077" points="611" reactiontime="+76" swimtime="00:00:27.35" resultid="8616" heatid="11414" lane="5" entrytime="00:00:27.11" entrycourse="SCM" />
                <RESULT eventid="6306" points="589" reactiontime="+80" swimtime="00:01:01.16" resultid="8617" heatid="11476" lane="8" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="527" reactiontime="+83" swimtime="00:02:19.87" resultid="8618" heatid="11567" lane="5" entrytime="00:02:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="8619" heatid="11593" lane="0" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="6467" points="559" reactiontime="+76" swimtime="00:00:30.49" resultid="11363" heatid="11537" lane="3" entrytime="00:00:30.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Kozanecka" birthdate="2001-06-08" gender="F" nation="POL" swrid="4749880" athleteid="8608">
              <RESULTS>
                <RESULT eventid="6094" points="689" reactiontime="+74" swimtime="00:02:36.33" resultid="8610" heatid="11424" lane="2" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="150" swimtime="00:01:59.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="711" reactiontime="+74" swimtime="00:02:50.09" resultid="8611" heatid="11454" lane="3" entrytime="00:02:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6323" points="658" reactiontime="+72" swimtime="00:01:12.65" resultid="8612" heatid="11486" lane="1" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6415" points="701" reactiontime="+74" swimtime="00:01:19.61" resultid="8613" heatid="11512" lane="3" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="640" reactiontime="+74" swimtime="00:02:22.90" resultid="8614" heatid="11559" lane="6" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" status="DNS" swimtime="00:00:00.00" resultid="8615" heatid="11588" lane="0" entrytime="00:01:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="7852" name="Plavecky klub Havirov">
          <ATHLETES>
            <ATHLETE firstname="Libor" lastname="Hracki" birthdate="1972-08-29" gender="M" nation="CZE" swrid="4934036" athleteid="7853">
              <RESULTS>
                <RESULT eventid="6272" points="681" swimtime="00:02:55.83" resultid="7854" heatid="11458" lane="9" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:23.08" />
                    <SPLIT distance="150" swimtime="00:02:08.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="601" reactiontime="+73" swimtime="00:01:19.57" resultid="7855" heatid="11518" lane="6" entrytime="00:01:25.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="544" reactiontime="+77" swimtime="00:02:24.64" resultid="7856" heatid="11567" lane="1" entrytime="00:02:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="615" swimtime="00:00:36.17" resultid="7857" heatid="11619" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="6738" points="581" reactiontime="+75" swimtime="00:05:12.12" resultid="7858" heatid="11634" lane="1" entrytime="00:05:30.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:52.63" />
                    <SPLIT distance="200" swimtime="00:02:32.70" />
                    <SPLIT distance="250" swimtime="00:03:13.29" />
                    <SPLIT distance="300" swimtime="00:03:53.90" />
                    <SPLIT distance="350" swimtime="00:04:34.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="8697" name="Stowarzyszenie Pływackie Masters Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Kieres" birthdate="1984-06-13" gender="M" nation="POL" license="101713700001" swrid="5282844" athleteid="8756">
              <RESULTS>
                <RESULT eventid="6111" points="413" reactiontime="+76" swimtime="00:02:50.84" resultid="8757" heatid="11426" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:21.93" />
                    <SPLIT distance="150" swimtime="00:02:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6272" points="473" swimtime="00:03:00.38" resultid="8758" heatid="11457" lane="4" entrytime="00:03:10.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:24.80" />
                    <SPLIT distance="150" swimtime="00:02:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="447" reactiontime="+73" swimtime="00:02:45.64" resultid="8759" heatid="11503" lane="6" entrytime="00:02:55.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="464" reactiontime="+69" swimtime="00:01:21.98" resultid="8760" heatid="11518" lane="2" entrytime="00:01:26.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="363" reactiontime="+74" swimtime="00:00:33.11" resultid="8761" heatid="11535" lane="2" entrytime="00:00:33.62" entrycourse="SCM" />
                <RESULT eventid="6636" points="437" reactiontime="+76" swimtime="00:01:12.73" resultid="8762" heatid="11593" lane="8" entrytime="00:01:14.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="445" reactiontime="+73" swimtime="00:00:37.79" resultid="8763" heatid="11618" lane="3" entrytime="00:00:39.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Gregorowicz" birthdate="1974-10-30" gender="M" nation="POL" license="101713700002" swrid="4992729" athleteid="8707">
              <RESULTS>
                <RESULT eventid="6077" points="792" reactiontime="+70" swimtime="00:00:25.79" resultid="8708" heatid="11414" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="6169" points="785" reactiontime="+82" swimtime="00:09:23.36" resultid="8709" heatid="11645" lane="3" entrytime="00:09:26.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="150" swimtime="00:01:42.78" />
                    <SPLIT distance="200" swimtime="00:02:18.57" />
                    <SPLIT distance="250" swimtime="00:02:54.53" />
                    <SPLIT distance="300" swimtime="00:03:30.23" />
                    <SPLIT distance="350" swimtime="00:04:05.88" />
                    <SPLIT distance="400" swimtime="00:04:41.66" />
                    <SPLIT distance="450" swimtime="00:05:17.17" />
                    <SPLIT distance="500" swimtime="00:05:52.57" />
                    <SPLIT distance="550" swimtime="00:06:28.28" />
                    <SPLIT distance="600" swimtime="00:07:03.55" />
                    <SPLIT distance="650" swimtime="00:07:38.69" />
                    <SPLIT distance="700" swimtime="00:08:13.90" />
                    <SPLIT distance="750" swimtime="00:08:48.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="801" reactiontime="+78" swimtime="00:02:21.73" resultid="8710" heatid="11504" lane="5" entrytime="00:02:20.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="769" reactiontime="+74" swimtime="00:00:28.03" resultid="8711" heatid="11537" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="6569" points="824" reactiontime="+73" swimtime="00:05:08.24" resultid="8712" heatid="11579" lane="6" entrytime="00:05:08.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                    <SPLIT distance="200" swimtime="00:02:31.28" />
                    <SPLIT distance="250" swimtime="00:03:15.78" />
                    <SPLIT distance="300" swimtime="00:03:59.26" />
                    <SPLIT distance="350" swimtime="00:04:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="849" reactiontime="+71" swimtime="00:01:01.81" resultid="8713" heatid="11596" lane="1" entrytime="00:01:01.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="742" reactiontime="+78" swimtime="00:04:31.60" resultid="8714" heatid="11638" lane="9" entrytime="00:04:34.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:39.28" />
                    <SPLIT distance="200" swimtime="00:02:13.49" />
                    <SPLIT distance="250" swimtime="00:02:48.14" />
                    <SPLIT distance="300" swimtime="00:03:22.82" />
                    <SPLIT distance="350" swimtime="00:03:57.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Łuczak" birthdate="1978-03-18" gender="M" nation="POL" license="501713700016" swrid="5416815" athleteid="8721">
              <RESULTS>
                <RESULT eventid="6077" points="530" swimtime="00:00:28.67" resultid="8722" heatid="11413" lane="9" entrytime="00:00:28.23" entrycourse="SCM" />
                <RESULT eventid="6272" points="516" swimtime="00:02:58.06" resultid="8723" heatid="11459" lane="9" entrytime="00:02:57.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:09.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="517" reactiontime="+78" swimtime="00:01:19.22" resultid="8724" heatid="11519" lane="7" entrytime="00:01:20.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="587" reactiontime="+65" swimtime="00:00:34.72" resultid="8725" heatid="11621" lane="1" entrytime="00:00:34.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mówiński" birthdate="1969-09-01" gender="M" nation="POL" license="501713700007" swrid="4992726" athleteid="8764">
              <RESULTS>
                <RESULT eventid="6169" points="471" reactiontime="+91" swimtime="00:11:30.90" resultid="8765" heatid="11646" lane="8" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:03.76" />
                    <SPLIT distance="200" swimtime="00:02:47.17" />
                    <SPLIT distance="250" swimtime="00:03:30.94" />
                    <SPLIT distance="300" swimtime="00:04:14.35" />
                    <SPLIT distance="350" swimtime="00:04:57.70" />
                    <SPLIT distance="400" swimtime="00:05:41.22" />
                    <SPLIT distance="450" swimtime="00:06:25.52" />
                    <SPLIT distance="500" swimtime="00:07:09.62" />
                    <SPLIT distance="550" swimtime="00:07:53.68" />
                    <SPLIT distance="600" swimtime="00:08:37.60" />
                    <SPLIT distance="650" swimtime="00:09:21.92" />
                    <SPLIT distance="700" swimtime="00:10:06.18" />
                    <SPLIT distance="750" swimtime="00:10:49.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="431" reactiontime="+87" swimtime="00:03:03.89" resultid="8766" heatid="11503" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="439" reactiontime="+84" swimtime="00:02:35.39" resultid="8767" heatid="11565" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="491" swimtime="00:05:30.16" resultid="8768" heatid="11633" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:18.40" />
                    <SPLIT distance="150" swimtime="00:02:00.65" />
                    <SPLIT distance="200" swimtime="00:02:43.23" />
                    <SPLIT distance="250" swimtime="00:03:26.11" />
                    <SPLIT distance="300" swimtime="00:04:09.14" />
                    <SPLIT distance="350" swimtime="00:04:52.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Grabowski" birthdate="1989-02-10" gender="M" nation="POL" license="501713700028" swrid="5230712" athleteid="8726">
              <RESULTS>
                <RESULT eventid="6077" points="574" swimtime="00:00:26.62" resultid="8727" heatid="11413" lane="4" entrytime="00:00:27.93" entrycourse="SCM" />
                <RESULT eventid="6306" points="532" reactiontime="+75" swimtime="00:01:00.51" resultid="8728" heatid="11474" lane="3" entrytime="00:01:04.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="8729" heatid="11493" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="6467" points="438" swimtime="00:00:30.10" resultid="8730" heatid="11537" lane="8" entrytime="00:00:30.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Matusiak vel Matuszewski" birthdate="1974-06-25" gender="M" nation="POL" license="501713700004" athleteid="8698">
              <RESULTS>
                <RESULT eventid="6077" points="407" swimtime="00:00:32.21" resultid="8699" heatid="11409" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="6238" points="286" reactiontime="+69" swimtime="00:00:42.29" resultid="8701" heatid="11446" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="6306" points="391" reactiontime="+79" swimtime="00:01:12.36" resultid="8702" heatid="11471" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="288" swimtime="00:00:38.88" resultid="8703" heatid="11533" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="6535" points="377" reactiontime="+83" swimtime="00:02:38.78" resultid="8704" heatid="11566" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="8705" heatid="11603" lane="3" entrytime="00:03:15.00" />
                <RESULT eventid="6738" points="403" reactiontime="+83" swimtime="00:05:32.76" resultid="8706" heatid="11634" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:01:58.88" />
                    <SPLIT distance="200" swimtime="00:02:41.10" />
                    <SPLIT distance="250" swimtime="00:03:23.49" />
                    <SPLIT distance="300" swimtime="00:04:06.82" />
                    <SPLIT distance="350" swimtime="00:04:50.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Dąbrowski" birthdate="1974-01-14" gender="M" nation="POL" license="501713700022" swrid="5355776" athleteid="8769">
              <RESULTS>
                <RESULT eventid="6169" points="498" swimtime="00:10:55.54" resultid="8770" heatid="11646" lane="1" entrytime="00:11:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:01:58.77" />
                    <SPLIT distance="200" swimtime="00:02:40.12" />
                    <SPLIT distance="250" swimtime="00:03:21.47" />
                    <SPLIT distance="300" swimtime="00:04:02.70" />
                    <SPLIT distance="350" swimtime="00:04:44.47" />
                    <SPLIT distance="400" swimtime="00:05:26.11" />
                    <SPLIT distance="450" swimtime="00:06:07.85" />
                    <SPLIT distance="500" swimtime="00:06:48.97" />
                    <SPLIT distance="550" swimtime="00:07:30.19" />
                    <SPLIT distance="600" swimtime="00:08:12.60" />
                    <SPLIT distance="650" swimtime="00:08:54.39" />
                    <SPLIT distance="700" swimtime="00:09:36.33" />
                    <SPLIT distance="750" swimtime="00:10:17.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="495" reactiontime="+73" swimtime="00:00:35.22" resultid="8771" heatid="11447" lane="2" entrytime="00:00:34.80" />
                <RESULT eventid="6306" points="499" reactiontime="+81" swimtime="00:01:06.68" resultid="8772" heatid="11474" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6501" points="476" reactiontime="+78" swimtime="00:01:16.04" resultid="8773" heatid="11548" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="492" reactiontime="+80" swimtime="00:02:25.30" resultid="8774" heatid="11567" lane="6" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="483" reactiontime="+79" swimtime="00:02:47.60" resultid="8775" heatid="11601" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:20.60" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="478" reactiontime="+91" swimtime="00:05:14.33" resultid="8776" heatid="11635" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:01:54.56" />
                    <SPLIT distance="200" swimtime="00:02:34.54" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:54.98" />
                    <SPLIT distance="350" swimtime="00:04:35.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gozdan" birthdate="1968-08-16" gender="M" nation="POL" license="501713700009" swrid="5230704" athleteid="8731">
              <RESULTS>
                <RESULT eventid="6077" points="380" reactiontime="+77" swimtime="00:00:33.81" resultid="8732" heatid="11406" lane="4" entrytime="00:00:35.20" entrycourse="SCM" />
                <RESULT eventid="6306" points="282" reactiontime="+84" swimtime="00:01:20.93" resultid="8733" heatid="11470" lane="3" entrytime="00:01:19.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="356" reactiontime="+84" swimtime="00:01:34.68" resultid="8734" heatid="11517" lane="4" entrytime="00:01:32.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="281" reactiontime="+76" swimtime="00:03:00.29" resultid="8735" heatid="11564" lane="5" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6704" points="386" reactiontime="+85" swimtime="00:00:42.24" resultid="8736" heatid="11617" lane="5" entrytime="00:00:42.60" entrycourse="SCM" />
                <RESULT eventid="6738" points="291" swimtime="00:06:32.80" resultid="8737" heatid="11632" lane="8" entrytime="00:06:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:19.95" />
                    <SPLIT distance="200" swimtime="00:03:09.57" />
                    <SPLIT distance="350" swimtime="00:05:44.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Karpisz" birthdate="1993-04-17" gender="M" nation="POL" swrid="4087166" athleteid="7843">
              <RESULTS>
                <RESULT eventid="6077" points="937" reactiontime="+73" swimtime="00:00:23.34" resultid="7844" heatid="11419" lane="6" entrytime="00:00:23.00" />
                <RESULT eventid="6111" points="795" reactiontime="+72" swimtime="00:02:10.10" resultid="7845" heatid="11433" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:01:01.35" />
                    <SPLIT distance="150" swimtime="00:01:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6238" points="836" reactiontime="+61" swimtime="00:00:26.59" resultid="7846" heatid="11450" lane="2" entrytime="00:00:26.02" />
                <RESULT comment="Czas lepszy od Rekordu Polski danej kat. wiek." eventid="6340" points="910" reactiontime="+72" swimtime="00:00:56.95" resultid="7847" heatid="11497" lane="5" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="859" reactiontime="+82" swimtime="00:00:24.93" resultid="7848" heatid="11542" lane="7" entrytime="00:00:24.50" />
                <RESULT eventid="6501" points="882" reactiontime="+64" swimtime="00:00:57.39" resultid="7849" heatid="11553" lane="4" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="7850" heatid="11597" lane="3" entrytime="00:00:54.50" />
                <RESULT eventid="6704" status="DNS" swimtime="00:00:00.00" resultid="7851" heatid="11623" lane="1" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Zembrzuski" birthdate="1992-02-28" gender="M" nation="POL" athleteid="7833">
              <RESULTS>
                <RESULT eventid="6111" status="DNS" swimtime="00:00:00.00" resultid="7834" heatid="11432" lane="5" entrytime="00:02:29.50" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="7835" heatid="11478" lane="9" entrytime="00:00:56.30" />
                <RESULT eventid="6374" reactiontime="+88" status="DNF" swimtime="00:00:00.00" resultid="7836" heatid="11503" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="686" reactiontime="+77" swimtime="00:00:25.93" resultid="7837" heatid="11541" lane="2" entrytime="00:00:26.60" />
                <RESULT eventid="6535" points="598" reactiontime="+82" swimtime="00:02:06.40" resultid="7838" heatid="11569" lane="6" entrytime="00:02:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:03.42" />
                    <SPLIT distance="150" swimtime="00:01:35.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Zaleska" birthdate="1988-01-17" gender="F" nation="POL" license="501713600012" swrid="5355784" athleteid="8738">
              <RESULTS>
                <RESULT eventid="6094" points="566" reactiontime="+81" swimtime="00:02:52.73" resultid="8739" heatid="11422" lane="2" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="580" reactiontime="+70" swimtime="00:22:01.69" resultid="8740" heatid="11650" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:19.07" />
                    <SPLIT distance="150" swimtime="00:02:01.17" />
                    <SPLIT distance="200" swimtime="00:02:43.38" />
                    <SPLIT distance="250" swimtime="00:03:26.00" />
                    <SPLIT distance="300" swimtime="00:04:08.58" />
                    <SPLIT distance="350" swimtime="00:04:51.53" />
                    <SPLIT distance="400" swimtime="00:05:35.37" />
                    <SPLIT distance="450" swimtime="00:06:18.91" />
                    <SPLIT distance="500" swimtime="00:07:03.00" />
                    <SPLIT distance="550" swimtime="00:07:47.11" />
                    <SPLIT distance="600" swimtime="00:08:31.86" />
                    <SPLIT distance="650" swimtime="00:09:16.42" />
                    <SPLIT distance="700" swimtime="00:10:00.73" />
                    <SPLIT distance="750" swimtime="00:10:45.49" />
                    <SPLIT distance="800" swimtime="00:11:30.47" />
                    <SPLIT distance="850" swimtime="00:12:15.34" />
                    <SPLIT distance="900" swimtime="00:12:59.98" />
                    <SPLIT distance="950" swimtime="00:13:44.74" />
                    <SPLIT distance="1000" swimtime="00:14:29.73" />
                    <SPLIT distance="1050" swimtime="00:15:14.76" />
                    <SPLIT distance="1100" swimtime="00:15:59.89" />
                    <SPLIT distance="1150" swimtime="00:16:44.84" />
                    <SPLIT distance="1200" swimtime="00:17:30.22" />
                    <SPLIT distance="1250" swimtime="00:18:15.36" />
                    <SPLIT distance="1300" swimtime="00:19:01.17" />
                    <SPLIT distance="1350" swimtime="00:19:46.83" />
                    <SPLIT distance="1400" swimtime="00:20:31.73" />
                    <SPLIT distance="1450" swimtime="00:21:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6220" points="539" reactiontime="+76" swimtime="00:00:36.64" resultid="8741" heatid="11440" lane="1" entrytime="00:00:38.50" />
                <RESULT eventid="6357" points="618" reactiontime="+76" swimtime="00:02:47.55" resultid="8742" heatid="11499" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:03.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="582" reactiontime="+71" swimtime="00:00:33.75" resultid="8743" heatid="11526" lane="1" entrytime="00:00:35.60" />
                <RESULT eventid="6552" points="519" reactiontime="+86" swimtime="00:06:11.47" resultid="8744" heatid="11574" lane="2" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:22.90" />
                    <SPLIT distance="150" swimtime="00:02:12.12" />
                    <SPLIT distance="200" swimtime="00:03:00.93" />
                    <SPLIT distance="250" swimtime="00:03:53.55" />
                    <SPLIT distance="300" swimtime="00:04:45.72" />
                    <SPLIT distance="350" swimtime="00:05:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="545" reactiontime="+79" swimtime="00:01:16.63" resultid="8745" heatid="11587" lane="5" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="553" reactiontime="+83" swimtime="00:05:28.21" resultid="8746" heatid="11627" lane="8" entrytime="00:05:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:00.27" />
                    <SPLIT distance="200" swimtime="00:02:42.38" />
                    <SPLIT distance="250" swimtime="00:03:24.75" />
                    <SPLIT distance="300" swimtime="00:04:07.46" />
                    <SPLIT distance="350" swimtime="00:04:49.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oriana" lastname="Kowalińska" birthdate="1993-03-19" gender="F" nation="POL" swrid="4086694" athleteid="7826">
              <RESULTS>
                <RESULT eventid="6145" points="798" reactiontime="+84" swimtime="00:09:59.82" resultid="7827" heatid="11643" lane="4" entrytime="00:09:59.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                    <SPLIT distance="200" swimtime="00:02:25.46" />
                    <SPLIT distance="250" swimtime="00:03:02.95" />
                    <SPLIT distance="300" swimtime="00:03:40.56" />
                    <SPLIT distance="350" swimtime="00:04:18.01" />
                    <SPLIT distance="400" swimtime="00:04:55.93" />
                    <SPLIT distance="450" swimtime="00:05:34.02" />
                    <SPLIT distance="500" swimtime="00:06:12.34" />
                    <SPLIT distance="550" swimtime="00:06:50.58" />
                    <SPLIT distance="600" swimtime="00:07:28.84" />
                    <SPLIT distance="650" swimtime="00:08:07.07" />
                    <SPLIT distance="700" swimtime="00:08:45.38" />
                    <SPLIT distance="750" swimtime="00:09:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6357" points="783" swimtime="00:02:29.54" resultid="7828" heatid="11499" lane="4" entrytime="00:02:29.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="678" reactiontime="+81" swimtime="00:00:31.40" resultid="7829" heatid="11528" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="6552" points="791" reactiontime="+83" swimtime="00:05:24.60" resultid="7830" heatid="11574" lane="4" entrytime="00:05:24.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                    <SPLIT distance="200" swimtime="00:02:35.99" />
                    <SPLIT distance="250" swimtime="00:03:23.07" />
                    <SPLIT distance="300" swimtime="00:04:10.83" />
                    <SPLIT distance="350" swimtime="00:04:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6618" points="698" reactiontime="+83" swimtime="00:01:08.74" resultid="7831" heatid="11588" lane="3" entrytime="00:01:08.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="762" reactiontime="+82" swimtime="00:04:53.19" resultid="7832" heatid="11628" lane="5" entrytime="00:04:55.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:48.03" />
                    <SPLIT distance="200" swimtime="00:02:25.32" />
                    <SPLIT distance="250" swimtime="00:03:02.57" />
                    <SPLIT distance="300" swimtime="00:03:40.18" />
                    <SPLIT distance="350" swimtime="00:04:17.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Konopacki" birthdate="1978-04-01" gender="M" nation="POL" license="501713700019" swrid="5282843" athleteid="8747">
              <RESULTS>
                <RESULT eventid="6111" points="543" reactiontime="+72" swimtime="00:02:36.74" resultid="8748" heatid="11425" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6203" points="654" reactiontime="+75" swimtime="00:19:08.31" resultid="8749" heatid="11652" lane="2" entrytime="00:19:03.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                    <SPLIT distance="200" swimtime="00:02:28.87" />
                    <SPLIT distance="250" swimtime="00:03:07.81" />
                    <SPLIT distance="300" swimtime="00:03:46.95" />
                    <SPLIT distance="350" swimtime="00:04:25.33" />
                    <SPLIT distance="400" swimtime="00:05:04.02" />
                    <SPLIT distance="450" swimtime="00:05:42.95" />
                    <SPLIT distance="500" swimtime="00:06:21.75" />
                    <SPLIT distance="550" swimtime="00:07:00.28" />
                    <SPLIT distance="600" swimtime="00:07:38.36" />
                    <SPLIT distance="650" swimtime="00:08:16.93" />
                    <SPLIT distance="700" swimtime="00:08:55.33" />
                    <SPLIT distance="750" swimtime="00:09:33.50" />
                    <SPLIT distance="800" swimtime="00:10:12.05" />
                    <SPLIT distance="850" swimtime="00:10:50.91" />
                    <SPLIT distance="900" swimtime="00:11:29.59" />
                    <SPLIT distance="950" swimtime="00:12:08.45" />
                    <SPLIT distance="1000" swimtime="00:12:47.38" />
                    <SPLIT distance="1050" swimtime="00:13:26.36" />
                    <SPLIT distance="1100" swimtime="00:14:04.97" />
                    <SPLIT distance="1150" swimtime="00:14:43.08" />
                    <SPLIT distance="1200" swimtime="00:15:21.19" />
                    <SPLIT distance="1250" swimtime="00:15:59.98" />
                    <SPLIT distance="1300" swimtime="00:16:38.31" />
                    <SPLIT distance="1350" swimtime="00:17:16.77" />
                    <SPLIT distance="1400" swimtime="00:17:54.95" />
                    <SPLIT distance="1450" swimtime="00:18:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="607" reactiontime="+69" swimtime="00:01:00.53" resultid="8750" heatid="11476" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="413" reactiontime="+72" swimtime="00:02:49.24" resultid="8751" heatid="11503" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:05.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="552" reactiontime="+70" swimtime="00:02:17.76" resultid="8752" heatid="11569" lane="2" entrytime="00:02:14.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="519" reactiontime="+71" swimtime="00:05:37.22" resultid="8753" heatid="11578" lane="4" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:03.26" />
                    <SPLIT distance="200" swimtime="00:02:45.55" />
                    <SPLIT distance="250" swimtime="00:03:34.38" />
                    <SPLIT distance="300" swimtime="00:04:23.67" />
                    <SPLIT distance="350" swimtime="00:05:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="563" reactiontime="+65" swimtime="00:02:37.95" resultid="8754" heatid="11605" lane="2" entrytime="00:02:38.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="572" swimtime="00:04:49.91" resultid="8755" heatid="11637" lane="0" entrytime="00:04:48.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                    <SPLIT distance="200" swimtime="00:02:22.78" />
                    <SPLIT distance="250" swimtime="00:03:00.35" />
                    <SPLIT distance="300" swimtime="00:03:38.25" />
                    <SPLIT distance="350" swimtime="00:04:15.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Lemańczyk" birthdate="1977-10-01" gender="M" nation="POL" license="501713700050" swrid="5537476" athleteid="8715">
              <RESULTS>
                <RESULT eventid="6077" points="331" reactiontime="+80" swimtime="00:00:34.48" resultid="8716" heatid="11406" lane="5" entrytime="00:00:35.97" />
                <RESULT eventid="6272" points="404" reactiontime="+83" swimtime="00:03:19.69" resultid="8717" heatid="11457" lane="2" entrytime="00:03:25.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6433" points="385" reactiontime="+77" swimtime="00:01:30.75" resultid="8718" heatid="11517" lane="6" entrytime="00:01:35.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="270" reactiontime="+91" swimtime="00:02:57.32" resultid="8719" heatid="11564" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="269" swimtime="00:06:20.61" resultid="8720" heatid="11632" lane="0" entrytime="00:06:27.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="200" swimtime="00:03:10.05" />
                    <SPLIT distance="250" swimtime="00:03:58.88" />
                    <SPLIT distance="300" swimtime="00:04:47.61" />
                    <SPLIT distance="350" swimtime="00:05:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Szczuka" birthdate="1992-08-16" gender="M" nation="POL" swrid="4806285" athleteid="7839">
              <RESULTS>
                <RESULT eventid="6111" points="522" reactiontime="+88" swimtime="00:02:26.66" resultid="7840" heatid="11432" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:08.09" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="577" reactiontime="+79" swimtime="00:01:06.06" resultid="7841" heatid="11495" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="587" reactiontime="+94" swimtime="00:05:18.81" resultid="7842" heatid="11578" lane="5" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:52.56" />
                    <SPLIT distance="200" swimtime="00:02:34.63" />
                    <SPLIT distance="250" swimtime="00:03:18.97" />
                    <SPLIT distance="300" swimtime="00:04:04.96" />
                    <SPLIT distance="350" swimtime="00:04:42.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+73" swimtime="00:01:41.09" resultid="8779" heatid="11582" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.59" />
                    <SPLIT distance="100" swimtime="00:00:48.13" />
                    <SPLIT distance="150" swimtime="00:01:14.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7843" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="7833" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="7839" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="8726" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6779" reactiontime="+75" swimtime="00:02:05.01" resultid="8782" heatid="12332" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:37.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8769" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="8721" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="8707" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="8747" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="6610" reactiontime="+85" swimtime="00:01:51.29" resultid="8780" heatid="11582" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:00:57.33" />
                    <SPLIT distance="150" swimtime="00:01:24.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8707" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="8721" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="8769" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="8747" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" reactiontime="+73" swimtime="00:01:52.37" resultid="8777" heatid="11435" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.05" />
                    <SPLIT distance="100" swimtime="00:00:49.03" />
                    <SPLIT distance="150" swimtime="00:01:19.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7843" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="7833" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="7826" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="8738" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6391" reactiontime="+77" swimtime="00:02:03.21" resultid="8778" heatid="11506" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:37.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8738" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="7843" number="2" reactiontime="-14" />
                    <RELAYPOSITION athleteid="7826" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7833" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="7476" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Mikołajczyk" birthdate="1984-01-01" gender="M" nation="POL" athleteid="7475">
              <RESULTS>
                <RESULT comment="O7 - Pływak użył urządzenie lub ubiór zwiększający szybkość, pływalność lub wytrzymałość (np. rękawice, łapki, płetwy, opaski czy substancje klejące)." eventid="6077" reactiontime="+81" status="DSQ" swimtime="00:00:00.00" resultid="7477" heatid="11413" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="6238" points="380" reactiontime="+73" swimtime="00:00:33.78" resultid="7478" heatid="11449" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="6340" status="DNS" swimtime="00:00:00.00" resultid="7479" heatid="11494" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="7480" heatid="11552" lane="2" entrytime="00:01:08.00" />
                <RESULT eventid="6535" points="485" reactiontime="+98" swimtime="00:02:21.85" resultid="7481" heatid="11569" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="471" swimtime="00:05:11.37" resultid="7482" heatid="11638" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                    <SPLIT distance="200" swimtime="00:02:27.53" />
                    <SPLIT distance="250" swimtime="00:03:08.03" />
                    <SPLIT distance="300" swimtime="00:03:49.25" />
                    <SPLIT distance="350" swimtime="00:04:30.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6836" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-01-01" gender="M" nation="POL" athleteid="6835">
              <RESULTS>
                <RESULT eventid="6077" points="323" swimtime="00:00:40.19" resultid="6837" heatid="11405" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="6169" points="363" reactiontime="+93" swimtime="00:14:44.67" resultid="6838" heatid="11648" lane="2" entrytime="00:15:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:44.18" />
                    <SPLIT distance="150" swimtime="00:02:39.34" />
                    <SPLIT distance="200" swimtime="00:03:34.39" />
                    <SPLIT distance="250" swimtime="00:04:29.13" />
                    <SPLIT distance="300" swimtime="00:05:23.82" />
                    <SPLIT distance="350" swimtime="00:06:18.75" />
                    <SPLIT distance="400" swimtime="00:07:14.29" />
                    <SPLIT distance="450" swimtime="00:08:10.11" />
                    <SPLIT distance="500" swimtime="00:09:06.06" />
                    <SPLIT distance="550" swimtime="00:10:02.61" />
                    <SPLIT distance="600" swimtime="00:10:59.70" />
                    <SPLIT distance="650" swimtime="00:11:56.16" />
                    <SPLIT distance="700" swimtime="00:12:52.72" />
                    <SPLIT distance="750" swimtime="00:13:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="277" swimtime="00:01:33.74" resultid="6839" heatid="11468" lane="6" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="222" swimtime="00:00:50.42" resultid="6840" heatid="11532" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="6535" points="287" reactiontime="+97" swimtime="00:03:31.33" resultid="6841" heatid="11563" lane="7" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                    <SPLIT distance="100" swimtime="00:01:43.92" />
                    <SPLIT distance="150" swimtime="00:02:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="322" swimtime="00:07:25.03" resultid="6842" heatid="11631" lane="0" entrytime="00:07:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:48.27" />
                    <SPLIT distance="150" swimtime="00:02:45.21" />
                    <SPLIT distance="200" swimtime="00:03:41.15" />
                    <SPLIT distance="250" swimtime="00:04:37.58" />
                    <SPLIT distance="300" swimtime="00:05:33.87" />
                    <SPLIT distance="350" swimtime="00:06:31.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="7266" name="Individual_Kyiv">
          <ATHLETES>
            <ATHLETE firstname="Serhii" lastname="Chernov" birthdate="1950-07-15" gender="M" nation="UKR" athleteid="7267">
              <RESULTS>
                <RESULT eventid="6077" points="135" reactiontime="+132" swimtime="00:00:55.24" resultid="7268" heatid="11404" lane="6" entrytime="00:00:55.99" entrycourse="LCM" />
                <RESULT eventid="6306" points="131" reactiontime="+131" swimtime="00:02:06.98" resultid="7269" heatid="11467" lane="5" entrytime="00:02:13.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01709" nation="POL" region="09" clubid="8796" name="iSwim Białystok">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Aleksandrowicz" birthdate="1968-08-05" gender="M" nation="POL" license="501709700261" athleteid="8828">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G3" eventid="6111" reactiontime="+77" status="DSQ" swimtime="00:00:00.00" resultid="8829" heatid="11429" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:34.58" />
                    <SPLIT distance="150" swimtime="00:02:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="196" reactiontime="+85" swimtime="00:03:58.95" resultid="8830" heatid="11503" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                    <SPLIT distance="100" swimtime="00:01:46.00" />
                    <SPLIT distance="150" swimtime="00:02:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6569" points="308" reactiontime="+81" swimtime="00:07:23.04" resultid="8831" heatid="11577" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:45.93" />
                    <SPLIT distance="150" swimtime="00:02:47.54" />
                    <SPLIT distance="200" swimtime="00:03:48.23" />
                    <SPLIT distance="250" swimtime="00:04:46.33" />
                    <SPLIT distance="300" swimtime="00:05:45.76" />
                    <SPLIT distance="350" swimtime="00:06:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" status="DNS" swimtime="00:00:00.00" resultid="8832" heatid="11592" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="6738" points="343" swimtime="00:06:11.87" resultid="8833" heatid="11633" lane="0" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                    <SPLIT distance="200" swimtime="00:02:56.38" />
                    <SPLIT distance="250" swimtime="00:03:45.79" />
                    <SPLIT distance="300" swimtime="00:04:34.84" />
                    <SPLIT distance="350" swimtime="00:05:24.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Iłendo" birthdate="1993-02-09" gender="M" nation="POL" license="117/09700014" swrid="4086405" athleteid="8817">
              <RESULTS>
                <RESULT eventid="6077" points="754" reactiontime="+67" swimtime="00:00:25.09" resultid="8818" heatid="11417" lane="9" entrytime="00:00:25.50" />
                <RESULT eventid="6238" points="631" reactiontime="+73" swimtime="00:00:29.20" resultid="8819" heatid="11449" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="8820" heatid="11478" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="6501" points="643" reactiontime="+76" swimtime="00:01:03.75" resultid="8821" heatid="11553" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6670" points="480" reactiontime="+77" swimtime="00:02:28.34" resultid="8822" heatid="11606" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" status="DNS" swimtime="00:00:00.00" resultid="11388" heatid="11571" lane="7" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Humbla" birthdate="1979-01-24" gender="M" nation="POL" license="117/09700001" swrid="4046250" athleteid="8812">
              <RESULTS>
                <RESULT eventid="6077" points="665" reactiontime="+71" swimtime="00:00:26.59" resultid="8813" heatid="11414" lane="6" entrytime="00:00:27.20" />
                <RESULT eventid="6467" status="DNS" swimtime="00:00:00.00" resultid="8815" heatid="11538" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="6704" points="604" reactiontime="+66" swimtime="00:00:34.40" resultid="8816" heatid="11621" lane="8" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Daszuta" birthdate="1973-03-12" gender="M" nation="POL" license="117/09700012" swrid="5421995" athleteid="8808">
              <RESULTS>
                <RESULT eventid="6077" points="619" reactiontime="+74" swimtime="00:00:28.00" resultid="8809" heatid="11414" lane="3" entrytime="00:00:27.19" />
                <RESULT eventid="6467" points="661" reactiontime="+77" swimtime="00:00:29.48" resultid="8810" heatid="11539" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="6704" points="720" reactiontime="+71" swimtime="00:00:33.79" resultid="8811" heatid="11621" lane="4" entrytime="00:00:33.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Stefanowska" birthdate="1974-10-23" gender="F" nation="POL" license="117/09600013" athleteid="8834">
              <RESULTS>
                <RESULT eventid="6145" status="DNS" swimtime="00:00:00.00" resultid="8835" heatid="11644" lane="3" entrytime="00:13:30.00" />
                <RESULT eventid="6289" status="DNS" swimtime="00:00:00.00" resultid="8836" heatid="11462" lane="6" entrytime="00:01:19.00" />
                <RESULT eventid="6450" status="DNS" swimtime="00:00:00.00" resultid="8837" heatid="11525" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="6721" status="DNS" swimtime="00:00:00.00" resultid="8838" heatid="11626" lane="7" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Iwaniuk-Mróz" birthdate="1979-07-17" gender="F" nation="POL" license="117/09600024" swrid="5470495" athleteid="8804">
              <RESULTS>
                <RESULT eventid="6059" points="608" reactiontime="+83" swimtime="00:00:31.01" resultid="8805" heatid="11399" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="6289" points="590" reactiontime="+68" swimtime="00:01:09.70" resultid="8806" heatid="11466" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6450" points="634" reactiontime="+76" swimtime="00:00:34.09" resultid="8807" heatid="11527" lane="0" entrytime="00:00:33.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Perkowski" birthdate="1996-06-10" gender="M" nation="POL" license="117/09700023" swrid="4290969" athleteid="8823">
              <RESULTS>
                <RESULT eventid="6077" points="780" reactiontime="+65" swimtime="00:00:24.81" resultid="8824" heatid="11417" lane="5" entrytime="00:00:24.90" />
                <RESULT eventid="6306" points="684" reactiontime="+64" swimtime="00:00:55.13" resultid="8825" heatid="11479" lane="1" entrytime="00:00:53.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="702" reactiontime="+58" swimtime="00:00:26.66" resultid="8826" heatid="11541" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="6636" points="745" swimtime="00:00:59.49" resultid="8827" heatid="11596" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elżbieta" lastname="Piwowarczyk" birthdate="1966-01-06" gender="F" nation="POL" license="501709600257" swrid="4186247" athleteid="8797">
              <RESULTS>
                <RESULT eventid="6059" points="595" reactiontime="+70" swimtime="00:00:34.15" resultid="8798" heatid="11397" lane="5" entrytime="00:00:35.30" entrycourse="SCM" />
                <RESULT eventid="6220" points="529" reactiontime="+74" swimtime="00:00:41.85" resultid="8799" heatid="11439" lane="4" entrytime="00:00:44.14" />
                <RESULT eventid="6289" points="538" reactiontime="+67" swimtime="00:01:17.09" resultid="8800" heatid="11463" lane="3" entrytime="00:01:19.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6484" points="542" reactiontime="+75" swimtime="00:01:31.22" resultid="8801" heatid="11545" lane="2" entrytime="00:01:33.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="490" reactiontime="+57" swimtime="00:02:54.68" resultid="8802" heatid="11557" lane="8" entrytime="00:02:56.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:23.66" />
                    <SPLIT distance="150" swimtime="00:02:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="511" reactiontime="+76" swimtime="00:03:16.37" resultid="8803" heatid="11599" lane="3" entrytime="00:03:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                    <SPLIT distance="150" swimtime="00:02:25.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Uściłko" birthdate="1995-07-13" gender="M" nation="POL" license="101709700260" swrid="4195032" athleteid="8839">
              <RESULTS>
                <RESULT eventid="6306" points="727" swimtime="00:00:54.01" resultid="8840" heatid="11478" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6535" points="782" swimtime="00:02:00.64" resultid="8841" heatid="11571" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                    <SPLIT distance="100" swimtime="00:00:59.36" />
                    <SPLIT distance="150" swimtime="00:01:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="796" reactiontime="+80" swimtime="00:04:21.34" resultid="8842" heatid="11638" lane="5" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:02.51" />
                    <SPLIT distance="150" swimtime="00:01:35.57" />
                    <SPLIT distance="200" swimtime="00:02:09.19" />
                    <SPLIT distance="250" swimtime="00:02:41.70" />
                    <SPLIT distance="300" swimtime="00:03:14.96" />
                    <SPLIT distance="350" swimtime="00:03:48.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="6610" status="DNS" swimtime="00:00:00.00" resultid="8845" heatid="11584" lane="3" entrytime="00:01:42.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8823" number="1" />
                    <RELAYPOSITION athleteid="8817" number="2" />
                    <RELAYPOSITION athleteid="8812" number="3" />
                    <RELAYPOSITION athleteid="8839" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="6779" reactiontime="+71" swimtime="00:01:55.95" resultid="8846" heatid="12332" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:30.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8817" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8812" number="2" reactiontime="+192" />
                    <RELAYPOSITION athleteid="8823" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="8839" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6128" swimtime="00:02:07.26" resultid="8843" heatid="11436" lane="1" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:00:59.01" />
                    <SPLIT distance="150" swimtime="00:01:33.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8808" number="1" />
                    <RELAYPOSITION athleteid="8804" number="2" />
                    <RELAYPOSITION athleteid="8797" number="3" />
                    <RELAYPOSITION athleteid="8828" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6391" status="DNS" swimtime="00:00:00.00" resultid="8844" heatid="11507" lane="9" entrytime="00:02:24.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8808" number="1" />
                    <RELAYPOSITION athleteid="8804" number="2" />
                    <RELAYPOSITION athleteid="8828" number="3" />
                    <RELAYPOSITION athleteid="8834" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8461" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Chodyna" birthdate="1967-01-01" gender="M" nation="POL" athleteid="8460">
              <RESULTS>
                <RESULT eventid="6077" points="774" reactiontime="+68" swimtime="00:00:28.34" resultid="8462" heatid="11411" lane="5" entrytime="00:00:29.80" />
                <RESULT eventid="6238" points="522" reactiontime="+81" swimtime="00:00:36.43" resultid="8463" heatid="11447" lane="9" entrytime="00:00:37.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02203" nation="POL" region="03" clubid="8920" name="KS AZS AWF Biała Podlaska">
          <ATHLETES>
            <ATHLETE firstname="Nikodem" lastname="Naróg" birthdate="2002-11-22" gender="M" nation="POL" license="102203700140" swrid="5136392" athleteid="8921">
              <RESULTS>
                <RESULT eventid="6077" points="856" reactiontime="+68" swimtime="00:00:24.16" resultid="8922" heatid="11418" lane="6" entrytime="00:00:24.27" entrycourse="SCM" />
                <RESULT eventid="6169" points="761" reactiontime="+67" swimtime="00:09:13.03" resultid="8923" heatid="11648" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:03.67" />
                    <SPLIT distance="150" swimtime="00:01:39.03" />
                    <SPLIT distance="200" swimtime="00:02:15.19" />
                    <SPLIT distance="250" swimtime="00:02:50.93" />
                    <SPLIT distance="300" swimtime="00:03:26.90" />
                    <SPLIT distance="350" swimtime="00:04:03.13" />
                    <SPLIT distance="400" swimtime="00:04:39.16" />
                    <SPLIT distance="450" swimtime="00:05:13.90" />
                    <SPLIT distance="500" swimtime="00:05:49.58" />
                    <SPLIT distance="550" swimtime="00:06:24.18" />
                    <SPLIT distance="600" swimtime="00:06:58.82" />
                    <SPLIT distance="650" swimtime="00:07:32.92" />
                    <SPLIT distance="700" swimtime="00:08:07.73" />
                    <SPLIT distance="750" swimtime="00:08:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6306" points="860" reactiontime="+72" swimtime="00:00:53.19" resultid="8924" heatid="11479" lane="2" entrytime="00:00:53.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6374" points="799" reactiontime="+69" swimtime="00:02:14.52" resultid="8925" heatid="11500" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="964" reactiontime="+69" swimtime="00:00:24.88" resultid="8926" heatid="11542" lane="1" entrytime="00:00:24.61" entrycourse="SCM" />
                <RESULT eventid="6535" points="751" reactiontime="+75" swimtime="00:02:01.05" resultid="8927" heatid="11561" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="100" swimtime="00:00:59.16" />
                    <SPLIT distance="150" swimtime="00:01:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6636" points="876" reactiontime="+70" swimtime="00:00:56.77" resultid="8928" heatid="11597" lane="2" entrytime="00:00:56.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6738" points="795" reactiontime="+83" swimtime="00:04:22.80" resultid="8929" heatid="11629" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:01:01.50" />
                    <SPLIT distance="150" swimtime="00:01:35.49" />
                    <SPLIT distance="200" swimtime="00:02:10.24" />
                    <SPLIT distance="250" swimtime="00:02:45.15" />
                    <SPLIT distance="300" swimtime="00:03:18.51" />
                    <SPLIT distance="350" swimtime="00:03:48.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8554" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Majos" birthdate="1996-01-01" gender="F" nation="POL" swrid="4290447" athleteid="8553">
              <RESULTS>
                <RESULT eventid="6094" points="652" reactiontime="+82" swimtime="00:02:42.52" resultid="8555" heatid="11424" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:02:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6145" points="759" reactiontime="+84" swimtime="00:10:09.88" resultid="8556" heatid="11643" lane="3" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                    <SPLIT distance="200" swimtime="00:02:25.43" />
                    <SPLIT distance="250" swimtime="00:03:03.66" />
                    <SPLIT distance="300" swimtime="00:03:41.93" />
                    <SPLIT distance="350" swimtime="00:04:20.83" />
                    <SPLIT distance="400" swimtime="00:04:59.86" />
                    <SPLIT distance="450" swimtime="00:05:38.70" />
                    <SPLIT distance="500" swimtime="00:06:17.57" />
                    <SPLIT distance="550" swimtime="00:06:56.04" />
                    <SPLIT distance="600" swimtime="00:07:35.13" />
                    <SPLIT distance="650" swimtime="00:08:13.91" />
                    <SPLIT distance="700" swimtime="00:08:52.86" />
                    <SPLIT distance="750" swimtime="00:09:31.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="6862" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Aleksandra" lastname="Sac" birthdate="1999-01-01" gender="F" nation="POL" swrid="4407794" athleteid="6861">
              <RESULTS>
                <RESULT eventid="6094" points="408" swimtime="00:03:06.10" resultid="6863" heatid="11422" lane="6" entrytime="00:03:09.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                    <SPLIT distance="150" swimtime="00:02:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6186" points="450" reactiontime="+90" swimtime="00:22:24.77" resultid="6864" heatid="11650" lane="3" entrytime="00:22:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:07.06" />
                    <SPLIT distance="200" swimtime="00:02:51.83" />
                    <SPLIT distance="250" swimtime="00:03:36.62" />
                    <SPLIT distance="300" swimtime="00:04:21.47" />
                    <SPLIT distance="350" swimtime="00:05:06.50" />
                    <SPLIT distance="400" swimtime="00:05:51.51" />
                    <SPLIT distance="450" swimtime="00:06:36.58" />
                    <SPLIT distance="500" swimtime="00:07:22.00" />
                    <SPLIT distance="550" swimtime="00:08:07.24" />
                    <SPLIT distance="600" swimtime="00:08:52.15" />
                    <SPLIT distance="650" swimtime="00:09:37.15" />
                    <SPLIT distance="700" swimtime="00:10:22.68" />
                    <SPLIT distance="750" swimtime="00:11:07.77" />
                    <SPLIT distance="800" swimtime="00:11:53.26" />
                    <SPLIT distance="850" swimtime="00:12:38.51" />
                    <SPLIT distance="900" swimtime="00:13:24.01" />
                    <SPLIT distance="950" swimtime="00:14:09.21" />
                    <SPLIT distance="1000" swimtime="00:14:54.71" />
                    <SPLIT distance="1050" swimtime="00:15:39.82" />
                    <SPLIT distance="1100" swimtime="00:16:25.44" />
                    <SPLIT distance="1150" swimtime="00:17:10.39" />
                    <SPLIT distance="1200" swimtime="00:17:56.21" />
                    <SPLIT distance="1250" swimtime="00:18:42.12" />
                    <SPLIT distance="1300" swimtime="00:19:27.64" />
                    <SPLIT distance="1350" swimtime="00:20:11.87" />
                    <SPLIT distance="1400" swimtime="00:20:57.50" />
                    <SPLIT distance="1450" swimtime="00:21:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6255" points="364" swimtime="00:03:32.62" resultid="6865" heatid="11453" lane="6" entrytime="00:03:35.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.59" />
                    <SPLIT distance="100" swimtime="00:01:41.89" />
                    <SPLIT distance="150" swimtime="00:02:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6518" points="411" swimtime="00:02:45.52" resultid="6866" heatid="11558" lane="6" entrytime="00:02:40.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6552" points="431" reactiontime="+80" swimtime="00:06:39.21" resultid="6867" heatid="11574" lane="7" entrytime="00:06:22.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:26.32" />
                    <SPLIT distance="200" swimtime="00:03:16.77" />
                    <SPLIT distance="250" swimtime="00:04:13.84" />
                    <SPLIT distance="300" swimtime="00:05:10.35" />
                    <SPLIT distance="350" swimtime="00:05:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6653" points="339" reactiontime="+84" swimtime="00:03:08.85" resultid="6868" heatid="11599" lane="4" entrytime="00:03:05.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:31.42" />
                    <SPLIT distance="150" swimtime="00:02:21.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6721" points="449" reactiontime="+70" swimtime="00:05:35.10" resultid="6869" heatid="11627" lane="5" entrytime="00:05:35.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:02:00.81" />
                    <SPLIT distance="200" swimtime="00:02:43.51" />
                    <SPLIT distance="250" swimtime="00:03:26.29" />
                    <SPLIT distance="300" swimtime="00:04:09.74" />
                    <SPLIT distance="350" swimtime="00:04:53.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" clubid="9678" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Kamil" lastname="Bernaś" birthdate="1984-02-13" gender="M" nation="POL" athleteid="9679">
              <RESULTS>
                <RESULT eventid="6306" points="485" reactiontime="+68" swimtime="00:01:02.83" resultid="9680" heatid="11467" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="425" reactiontime="+71" swimtime="00:00:31.41" resultid="9681" heatid="11531" lane="6" />
                <RESULT eventid="6535" points="419" reactiontime="+71" swimtime="00:02:28.95" resultid="9682" heatid="11561" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:48.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kaczmarek" birthdate="1983-07-27" gender="M" nation="POL" swrid="5537972" athleteid="9689">
              <RESULTS>
                <RESULT eventid="6077" status="DNS" swimtime="00:00:00.00" resultid="9690" heatid="11413" lane="8" entrytime="00:00:28.10" entrycourse="SCM" />
                <RESULT eventid="6238" status="DNS" swimtime="00:00:00.00" resultid="9691" heatid="11448" lane="7" entrytime="00:00:33.11" entrycourse="SCM" />
                <RESULT eventid="6306" status="DNS" swimtime="00:00:00.00" resultid="9692" heatid="11475" lane="2" entrytime="00:01:02.80" entrycourse="SCM" />
                <RESULT eventid="6501" status="DNS" swimtime="00:00:00.00" resultid="9693" heatid="11548" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Thiem" birthdate="1963-01-01" gender="M" nation="POL" athleteid="9914">
              <RESULTS>
                <RESULT eventid="6535" points="210" swimtime="00:03:33.15" resultid="9915" heatid="11561" lane="9" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                    <SPLIT distance="100" swimtime="00:01:47.31" />
                    <SPLIT distance="150" swimtime="00:02:41.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Juszkiewicz" birthdate="1974-05-10" gender="M" nation="POL" swrid="5537971" athleteid="9694">
              <RESULTS>
                <RESULT eventid="6306" points="461" reactiontime="+76" swimtime="00:01:08.46" resultid="9695" heatid="11473" lane="0" entrytime="00:01:09.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="340" reactiontime="+81" swimtime="00:00:36.76" resultid="9696" heatid="11531" lane="1" />
                <RESULT eventid="6670" status="DNS" swimtime="00:00:00.00" resultid="9697" heatid="11602" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Jankowiak" birthdate="1981-12-27" gender="M" nation="POL" athleteid="9683">
              <RESULTS>
                <RESULT eventid="6077" points="492" reactiontime="+69" swimtime="00:00:29.40" resultid="9684" heatid="11402" lane="5" />
                <RESULT eventid="6169" points="420" reactiontime="+77" swimtime="00:11:22.89" resultid="9685" heatid="11648" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                    <SPLIT distance="200" swimtime="00:02:45.54" />
                    <SPLIT distance="250" swimtime="00:03:29.47" />
                    <SPLIT distance="300" swimtime="00:04:13.07" />
                    <SPLIT distance="350" swimtime="00:04:56.98" />
                    <SPLIT distance="400" swimtime="00:05:40.10" />
                    <SPLIT distance="450" swimtime="00:06:23.54" />
                    <SPLIT distance="500" swimtime="00:07:06.81" />
                    <SPLIT distance="550" swimtime="00:07:50.43" />
                    <SPLIT distance="600" swimtime="00:08:33.51" />
                    <SPLIT distance="650" swimtime="00:10:00.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6340" points="426" reactiontime="+72" swimtime="00:01:19.50" resultid="9686" heatid="11487" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6467" points="403" reactiontime="+76" swimtime="00:00:34.02" resultid="9687" heatid="11529" lane="3" />
                <RESULT eventid="6535" points="389" reactiontime="+74" swimtime="00:02:34.77" resultid="9688" heatid="11560" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:53.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="MKP BOBRY DEBICA" version="Build 23153">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Dębica" name="Otwarte Mistrzostwa Masters Polski w pływaniu" course="LCM" deadline="2013-05-30" nation="POL" organizer="MKP BOBRY DĘBICA" organizer.url="http://bobrydebica.com" timing="AUTOMATIC">
      <AGEDATE value="2013-12-31" type="YEAR" />
      <POOL lanemin="1" lanemax="8" />
      <POINTTABLE pointtableid="1008" name="DSV Master Performance Table" version="2004" />
      <SESSIONS>
        <SESSION date="2013-06-14" daytime="15:30" name="I Blok" number="1" warmupfrom="13:50" warmupuntil="14:50">
          <EVENTS>
            <EVENT eventid="1061" daytime="15:30" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1062" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2314" />
                    <RANKING order="2" place="2" resultid="5741" />
                    <RANKING order="3" place="3" resultid="5748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2516" />
                    <RANKING order="2" place="2" resultid="4420" />
                    <RANKING order="3" place="3" resultid="6704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                    <RANKING order="2" place="2" resultid="6733" />
                    <RANKING order="3" place="3" resultid="4532" />
                    <RANKING order="4" place="4" resultid="5638" />
                    <RANKING order="5" place="-1" resultid="4497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2510" />
                    <RANKING order="2" place="2" resultid="4559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3133" />
                    <RANKING order="2" place="2" resultid="5733" />
                    <RANKING order="3" place="3" resultid="4538" />
                    <RANKING order="4" place="4" resultid="5857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5831" />
                    <RANKING order="2" place="2" resultid="6018" />
                    <RANKING order="3" place="3" resultid="3784" />
                    <RANKING order="4" place="4" resultid="5031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3107" />
                    <RANKING order="2" place="2" resultid="5786" />
                    <RANKING order="3" place="3" resultid="3840" />
                    <RANKING order="4" place="4" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5777" />
                    <RANKING order="2" place="2" resultid="3102" />
                    <RANKING order="3" place="3" resultid="4609" />
                    <RANKING order="4" place="4" resultid="9030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2694" />
                    <RANKING order="2" place="2" resultid="2683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5804" />
                    <RANKING order="2" place="-1" resultid="2715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1075" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1076" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1063" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10095" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10096" daytime="15:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10097" daytime="15:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10098" daytime="15:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10099" daytime="15:35" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="15:35" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1719" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2336" />
                    <RANKING order="2" place="2" resultid="5620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1720" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4645" />
                    <RANKING order="2" place="2" resultid="2354" />
                    <RANKING order="3" place="3" resultid="5771" />
                    <RANKING order="4" place="4" resultid="4512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1721" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2258" />
                    <RANKING order="2" place="2" resultid="9036" />
                    <RANKING order="3" place="3" resultid="4398" />
                    <RANKING order="4" place="4" resultid="4270" />
                    <RANKING order="5" place="5" resultid="4289" />
                    <RANKING order="6" place="6" resultid="7962" />
                    <RANKING order="7" place="7" resultid="4517" />
                    <RANKING order="8" place="-1" resultid="4554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1722" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4362" />
                    <RANKING order="2" place="2" resultid="5645" />
                    <RANKING order="3" place="3" resultid="3807" />
                    <RANKING order="4" place="4" resultid="8182" />
                    <RANKING order="5" place="5" resultid="2248" />
                    <RANKING order="6" place="6" resultid="4688" />
                    <RANKING order="7" place="-1" resultid="4507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1723" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3745" />
                    <RANKING order="2" place="2" resultid="2600" />
                    <RANKING order="3" place="3" resultid="2688" />
                    <RANKING order="4" place="4" resultid="5993" />
                    <RANKING order="5" place="5" resultid="5938" />
                    <RANKING order="6" place="6" resultid="3761" />
                    <RANKING order="7" place="7" resultid="5859" />
                    <RANKING order="8" place="8" resultid="5864" />
                    <RANKING order="9" place="9" resultid="9046" />
                    <RANKING order="10" place="-1" resultid="2636" />
                    <RANKING order="11" place="-1" resultid="3824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1724" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2207" />
                    <RANKING order="2" place="2" resultid="2502" />
                    <RANKING order="3" place="3" resultid="7695" />
                    <RANKING order="4" place="4" resultid="7679" />
                    <RANKING order="5" place="5" resultid="3793" />
                    <RANKING order="6" place="6" resultid="6695" />
                    <RANKING order="7" place="7" resultid="3555" />
                    <RANKING order="8" place="8" resultid="6011" />
                    <RANKING order="9" place="9" resultid="3172" />
                    <RANKING order="10" place="-1" resultid="5722" />
                    <RANKING order="11" place="-1" resultid="6752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1725" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2378" />
                    <RANKING order="2" place="2" resultid="5820" />
                    <RANKING order="3" place="3" resultid="4489" />
                    <RANKING order="4" place="4" resultid="2498" />
                    <RANKING order="5" place="5" resultid="3163" />
                    <RANKING order="6" place="6" resultid="2706" />
                    <RANKING order="7" place="7" resultid="9052" />
                    <RANKING order="8" place="-1" resultid="5668" />
                    <RANKING order="9" place="-1" resultid="6006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1726" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5630" />
                    <RANKING order="2" place="2" resultid="4654" />
                    <RANKING order="3" place="3" resultid="3124" />
                    <RANKING order="4" place="4" resultid="5999" />
                    <RANKING order="5" place="5" resultid="3778" />
                    <RANKING order="6" place="6" resultid="3858" />
                    <RANKING order="7" place="7" resultid="5684" />
                    <RANKING order="8" place="8" resultid="8171" />
                    <RANKING order="9" place="9" resultid="3195" />
                    <RANKING order="10" place="-1" resultid="2776" />
                    <RANKING order="11" place="-1" resultid="3180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1727" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4630" />
                    <RANKING order="2" place="2" resultid="8161" />
                    <RANKING order="3" place="3" resultid="4412" />
                    <RANKING order="4" place="4" resultid="3565" />
                    <RANKING order="5" place="5" resultid="2646" />
                    <RANKING order="6" place="6" resultid="5036" />
                    <RANKING order="7" place="7" resultid="4353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1728" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2263" />
                    <RANKING order="2" place="2" resultid="6684" />
                    <RANKING order="3" place="3" resultid="2700" />
                    <RANKING order="4" place="4" resultid="2710" />
                    <RANKING order="5" place="5" resultid="3078" />
                    <RANKING order="6" place="6" resultid="2591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1729" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2661" />
                    <RANKING order="2" place="2" resultid="2641" />
                    <RANKING order="3" place="3" resultid="5021" />
                    <RANKING order="4" place="4" resultid="3215" />
                    <RANKING order="5" place="5" resultid="3245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1730" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2195" />
                    <RANKING order="2" place="2" resultid="6725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1731" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1732" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1733" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10100" daytime="15:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10101" daytime="15:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10102" daytime="15:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10103" daytime="15:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10104" daytime="15:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10105" daytime="15:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10106" daytime="15:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10107" daytime="15:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10108" daytime="15:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10109" daytime="15:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10110" daytime="15:50" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="15:50" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1734" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2315" />
                    <RANKING order="2" place="2" resultid="5849" />
                    <RANKING order="3" place="3" resultid="2763" />
                    <RANKING order="4" place="4" resultid="2489" />
                    <RANKING order="5" place="5" resultid="4371" />
                    <RANKING order="6" place="6" resultid="7713" />
                    <RANKING order="7" place="7" resultid="5742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1735" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4421" />
                    <RANKING order="2" place="2" resultid="5813" />
                    <RANKING order="3" place="3" resultid="5766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1737" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2676" />
                    <RANKING order="2" place="2" resultid="3134" />
                    <RANKING order="3" place="3" resultid="5734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6744" />
                    <RANKING order="2" place="2" resultid="3785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1740" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5970" />
                    <RANKING order="2" place="2" resultid="3112" />
                    <RANKING order="3" place="3" resultid="9024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1741" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4996" />
                    <RANKING order="2" place="2" resultid="5778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1742" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1743" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1744" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1745" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1746" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1747" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1748" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10111" daytime="15:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10112" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10113" daytime="16:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="16:05" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1749" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2631" />
                    <RANKING order="2" place="2" resultid="2559" />
                    <RANKING order="3" place="3" resultid="5621" />
                    <RANKING order="4" place="4" resultid="7956" />
                    <RANKING order="5" place="-1" resultid="5866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1750" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4399" />
                    <RANKING order="2" place="2" resultid="4294" />
                    <RANKING order="3" place="3" resultid="5659" />
                    <RANKING order="4" place="4" resultid="4381" />
                    <RANKING order="5" place="5" resultid="4518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3262" />
                    <RANKING order="2" place="2" resultid="4363" />
                    <RANKING order="3" place="3" resultid="3801" />
                    <RANKING order="4" place="4" resultid="3738" />
                    <RANKING order="5" place="5" resultid="5646" />
                    <RANKING order="6" place="6" resultid="7946" />
                    <RANKING order="7" place="7" resultid="4274" />
                    <RANKING order="8" place="-1" resultid="6762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3746" />
                    <RANKING order="2" place="2" resultid="2689" />
                    <RANKING order="3" place="3" resultid="3255" />
                    <RANKING order="4" place="4" resultid="3231" />
                    <RANKING order="5" place="5" resultid="3762" />
                    <RANKING order="6" place="-1" resultid="3825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2208" />
                    <RANKING order="2" place="2" resultid="6696" />
                    <RANKING order="3" place="3" resultid="3556" />
                    <RANKING order="4" place="4" resultid="6689" />
                    <RANKING order="5" place="-1" resultid="2832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4490" />
                    <RANKING order="2" place="2" resultid="6666" />
                    <RANKING order="3" place="3" resultid="2379" />
                    <RANKING order="4" place="4" resultid="3770" />
                    <RANKING order="5" place="5" resultid="4625" />
                    <RANKING order="6" place="6" resultid="3164" />
                    <RANKING order="7" place="7" resultid="5669" />
                    <RANKING order="8" place="8" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2328" />
                    <RANKING order="2" place="2" resultid="5014" />
                    <RANKING order="3" place="3" resultid="3181" />
                    <RANKING order="4" place="-1" resultid="2758" />
                    <RANKING order="5" place="-1" resultid="2777" />
                    <RANKING order="6" place="-1" resultid="3125" />
                    <RANKING order="7" place="-1" resultid="4699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6712" />
                    <RANKING order="2" place="2" resultid="5953" />
                    <RANKING order="3" place="3" resultid="2478" />
                    <RANKING order="4" place="4" resultid="3566" />
                    <RANKING order="5" place="5" resultid="4413" />
                    <RANKING order="6" place="6" resultid="3753" />
                    <RANKING order="7" place="7" resultid="3224" />
                    <RANKING order="8" place="8" resultid="4354" />
                    <RANKING order="9" place="9" resultid="3187" />
                    <RANKING order="10" place="10" resultid="3581" />
                    <RANKING order="11" place="-1" resultid="4407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1758" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2264" />
                    <RANKING order="2" place="2" resultid="4596" />
                    <RANKING order="3" place="3" resultid="7717" />
                    <RANKING order="4" place="4" resultid="3079" />
                    <RANKING order="5" place="5" resultid="2592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3216" />
                    <RANKING order="2" place="2" resultid="3246" />
                    <RANKING order="3" place="3" resultid="5753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1760" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1761" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1762" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1763" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10114" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10115" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10116" daytime="16:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10117" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10118" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10119" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10120" daytime="16:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10121" daytime="16:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10122" daytime="16:40" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1125" daytime="16:40" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10304" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1157" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4427" />
                    <RANKING order="2" place="2" resultid="4567" />
                    <RANKING order="3" place="3" resultid="4329" />
                    <RANKING order="4" place="4" resultid="8140" />
                    <RANKING order="5" place="-1" resultid="7725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5665" />
                    <RANKING order="2" place="2" resultid="5892" />
                    <RANKING order="3" place="3" resultid="6770" />
                    <RANKING order="4" place="4" resultid="4331" />
                    <RANKING order="5" place="-1" resultid="9051" />
                    <RANKING order="6" place="-1" resultid="4570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5894" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="3872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2721" />
                    <RANKING order="2" place="2" resultid="2722" />
                    <RANKING order="3" place="3" resultid="9476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2719" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10123" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10124" daytime="16:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10125" daytime="16:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="16:50" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1764" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5871" />
                    <RANKING order="2" place="2" resultid="4372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1765" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2243" />
                    <RANKING order="2" place="2" resultid="6705" />
                    <RANKING order="3" place="3" resultid="7690" />
                    <RANKING order="4" place="4" resultid="8178" />
                    <RANKING order="5" place="5" resultid="4526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1766" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1767" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1768" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4539" />
                    <RANKING order="2" place="2" resultid="3866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1769" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2364" />
                    <RANKING order="2" place="2" resultid="5652" />
                    <RANKING order="3" place="3" resultid="2784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1770" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5971" />
                    <RANKING order="2" place="2" resultid="5787" />
                    <RANKING order="3" place="3" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1771" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1772" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1773" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1774" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1775" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1776" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1777" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1778" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10293" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10294" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10295" daytime="17:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1711" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1162" daytime="17:45" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1779" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1780" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2348" />
                    <RANKING order="2" place="2" resultid="4646" />
                    <RANKING order="3" place="3" resultid="2355" />
                    <RANKING order="4" place="4" resultid="4316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1781" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4295" />
                    <RANKING order="2" place="2" resultid="2770" />
                    <RANKING order="3" place="3" resultid="6677" />
                    <RANKING order="4" place="4" resultid="6703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1782" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2369" />
                    <RANKING order="2" place="2" resultid="8183" />
                    <RANKING order="3" place="3" resultid="5727" />
                    <RANKING order="4" place="4" resultid="4310" />
                    <RANKING order="5" place="-1" resultid="6763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1783" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5860" />
                    <RANKING order="2" place="2" resultid="3232" />
                    <RANKING order="3" place="3" resultid="2637" />
                    <RANKING order="4" place="4" resultid="2483" />
                    <RANKING order="5" place="5" resultid="5929" />
                    <RANKING order="6" place="6" resultid="4279" />
                    <RANKING order="7" place="7" resultid="6741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1784" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4637" />
                    <RANKING order="2" place="2" resultid="7684" />
                    <RANKING order="3" place="3" resultid="5674" />
                    <RANKING order="4" place="4" resultid="5709" />
                    <RANKING order="5" place="5" resultid="5837" />
                    <RANKING order="6" place="6" resultid="6012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1785" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2499" />
                    <RANKING order="2" place="2" resultid="2792" />
                    <RANKING order="3" place="3" resultid="6717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1786" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5631" />
                    <RANKING order="2" place="2" resultid="5980" />
                    <RANKING order="3" place="3" resultid="3850" />
                    <RANKING order="4" place="4" resultid="3238" />
                    <RANKING order="5" place="-1" resultid="2187" />
                    <RANKING order="6" place="-1" resultid="4700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1787" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3092" />
                    <RANKING order="2" place="2" resultid="5037" />
                    <RANKING order="3" place="3" resultid="2745" />
                    <RANKING order="4" place="4" resultid="3582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1788" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1789" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2662" />
                    <RANKING order="2" place="2" resultid="5022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1790" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1791" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1792" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1793" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10296" daytime="17:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10297" daytime="18:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10298" daytime="18:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10299" daytime="18:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10300" daytime="19:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10301" daytime="19:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1709" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2013-06-15" daytime="09:00" name="2 Blok" number="2" warmupfrom="07:40" warmupuntil="08:40">
          <EVENTS>
            <EVENT eventid="1178" daytime="09:00" gender="F" number="8" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1794" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2730" />
                    <RANKING order="2" place="2" resultid="5844" />
                    <RANKING order="3" place="3" resultid="2764" />
                    <RANKING order="4" place="4" resultid="5850" />
                    <RANKING order="5" place="5" resultid="2490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1795" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8153" />
                    <RANKING order="2" place="2" resultid="2517" />
                    <RANKING order="3" place="3" resultid="5814" />
                    <RANKING order="4" place="4" resultid="7969" />
                    <RANKING order="5" place="5" resultid="4422" />
                    <RANKING order="6" place="6" resultid="2572" />
                    <RANKING order="7" place="7" resultid="8179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1796" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4392" />
                    <RANKING order="2" place="2" resultid="3270" />
                    <RANKING order="3" place="3" resultid="4267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1797" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1798" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3135" />
                    <RANKING order="2" place="2" resultid="5735" />
                    <RANKING order="3" place="3" resultid="4540" />
                    <RANKING order="4" place="4" resultid="5882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1799" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5761" />
                    <RANKING order="2" place="2" resultid="6019" />
                    <RANKING order="3" place="3" resultid="2785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1800" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5972" />
                    <RANKING order="2" place="2" resultid="3204" />
                    <RANKING order="3" place="-1" resultid="3108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1801" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4997" />
                    <RANKING order="2" place="2" resultid="5779" />
                    <RANKING order="3" place="3" resultid="3103" />
                    <RANKING order="4" place="4" resultid="7703" />
                    <RANKING order="5" place="5" resultid="2606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1802" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2695" />
                    <RANKING order="2" place="2" resultid="2613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1803" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4588" />
                    <RANKING order="2" place="2" resultid="2716" />
                    <RANKING order="3" place="3" resultid="4502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1804" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1805" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6738" />
                    <RANKING order="2" place="2" resultid="4666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1806" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1807" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1808" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10126" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10127" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10128" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10129" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10130" daytime="09:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="09:05" gender="M" number="9" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1809" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4477" />
                    <RANKING order="2" place="2" resultid="7957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1810" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4647" />
                    <RANKING order="2" place="2" resultid="2555" />
                    <RANKING order="3" place="3" resultid="4484" />
                    <RANKING order="4" place="4" resultid="2357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1811" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4296" />
                    <RANKING order="2" place="2" resultid="5660" />
                    <RANKING order="3" place="3" resultid="6678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1812" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3739" />
                    <RANKING order="2" place="2" resultid="2249" />
                    <RANKING order="3" place="3" resultid="3815" />
                    <RANKING order="4" place="4" resultid="4301" />
                    <RANKING order="5" place="5" resultid="4275" />
                    <RANKING order="6" place="6" resultid="5828" />
                    <RANKING order="7" place="-1" resultid="6764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1813" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2690" />
                    <RANKING order="2" place="2" resultid="3826" />
                    <RANKING order="3" place="3" resultid="5994" />
                    <RANKING order="4" place="4" resultid="2253" />
                    <RANKING order="5" place="5" resultid="5939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1814" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6697" />
                    <RANKING order="2" place="2" resultid="2337" />
                    <RANKING order="3" place="3" resultid="2798" />
                    <RANKING order="4" place="4" resultid="4638" />
                    <RANKING order="5" place="5" resultid="5675" />
                    <RANKING order="6" place="6" resultid="6013" />
                    <RANKING order="7" place="-1" resultid="6753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1815" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4491" />
                    <RANKING order="2" place="2" resultid="2380" />
                    <RANKING order="3" place="3" resultid="5821" />
                    <RANKING order="4" place="4" resultid="3165" />
                    <RANKING order="5" place="5" resultid="2812" />
                    <RANKING order="6" place="6" resultid="2707" />
                    <RANKING order="7" place="7" resultid="7953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1816" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5632" />
                    <RANKING order="2" place="2" resultid="3126" />
                    <RANKING order="3" place="3" resultid="6000" />
                    <RANKING order="4" place="4" resultid="10302" />
                    <RANKING order="5" place="5" resultid="3182" />
                    <RANKING order="6" place="6" resultid="3859" />
                    <RANKING order="7" place="7" resultid="3196" />
                    <RANKING order="8" place="8" resultid="2587" />
                    <RANKING order="9" place="-1" resultid="2188" />
                    <RANKING order="10" place="-1" resultid="2759" />
                    <RANKING order="11" place="-1" resultid="4547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1817" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8162" />
                    <RANKING order="2" place="2" resultid="5038" />
                    <RANKING order="3" place="3" resultid="3093" />
                    <RANKING order="4" place="4" resultid="3832" />
                    <RANKING order="5" place="5" resultid="3754" />
                    <RANKING order="6" place="6" resultid="3567" />
                    <RANKING order="7" place="7" resultid="4355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1818" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4597" />
                    <RANKING order="2" place="2" resultid="2657" />
                    <RANKING order="3" place="3" resultid="3080" />
                    <RANKING order="4" place="4" resultid="2711" />
                    <RANKING order="5" place="5" resultid="6685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1819" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2663" />
                    <RANKING order="2" place="2" resultid="3217" />
                    <RANKING order="3" place="3" resultid="5023" />
                    <RANKING order="4" place="4" resultid="5946" />
                    <RANKING order="5" place="5" resultid="3247" />
                    <RANKING order="6" place="6" resultid="2623" />
                    <RANKING order="7" place="7" resultid="5754" />
                    <RANKING order="8" place="8" resultid="3574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1820" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3210" />
                    <RANKING order="2" place="2" resultid="5046" />
                    <RANKING order="3" place="3" resultid="6727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1821" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8145" />
                    <RANKING order="2" place="2" resultid="2565" />
                    <RANKING order="3" place="3" resultid="5706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1822" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1823" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10131" daytime="09:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10132" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10133" daytime="09:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10134" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10135" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10136" daytime="09:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10137" daytime="09:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10138" daytime="09:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10139" daytime="09:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10140" daytime="09:20" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="09:20" gender="F" number="10" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1824" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2316" />
                    <RANKING order="2" place="2" resultid="2731" />
                    <RANKING order="3" place="3" resultid="5749" />
                    <RANKING order="4" place="4" resultid="5845" />
                    <RANKING order="5" place="5" resultid="5872" />
                    <RANKING order="6" place="6" resultid="5851" />
                    <RANKING order="7" place="7" resultid="4373" />
                    <RANKING order="8" place="8" resultid="5743" />
                    <RANKING order="9" place="-1" resultid="5879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1825" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2518" />
                    <RANKING order="2" place="2" resultid="5815" />
                    <RANKING order="3" place="3" resultid="8154" />
                    <RANKING order="4" place="4" resultid="6671" />
                    <RANKING order="5" place="5" resultid="2573" />
                    <RANKING order="6" place="6" resultid="4471" />
                    <RANKING order="7" place="7" resultid="6706" />
                    <RANKING order="8" place="8" resultid="7691" />
                    <RANKING order="9" place="9" resultid="4527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1826" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6029" />
                    <RANKING order="2" place="2" resultid="4393" />
                    <RANKING order="3" place="3" resultid="5640" />
                    <RANKING order="4" place="4" resultid="4533" />
                    <RANKING order="5" place="5" resultid="6734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1827" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4562" />
                    <RANKING order="2" place="2" resultid="6721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1828" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="4541" />
                    <RANKING order="3" place="3" resultid="3867" />
                    <RANKING order="4" place="4" resultid="4284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1829" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2365" />
                    <RANKING order="2" place="2" resultid="5762" />
                    <RANKING order="3" place="3" resultid="6020" />
                    <RANKING order="4" place="4" resultid="5653" />
                    <RANKING order="5" place="5" resultid="2786" />
                    <RANKING order="6" place="-1" resultid="3786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1830" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3113" />
                    <RANKING order="2" place="2" resultid="5973" />
                    <RANKING order="3" place="3" resultid="3205" />
                    <RANKING order="4" place="4" resultid="6025" />
                    <RANKING order="5" place="5" resultid="3841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1831" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1832" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5004" />
                    <RANKING order="2" place="2" resultid="2684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1833" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4503" />
                    <RANKING order="2" place="2" resultid="5806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1834" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1835" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1836" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1837" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1838" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10141" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10142" daytime="09:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10143" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10144" daytime="09:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10145" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10146" daytime="09:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="09:35" gender="M" number="11" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1839" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4478" />
                    <RANKING order="2" place="2" resultid="2560" />
                    <RANKING order="3" place="3" resultid="5622" />
                    <RANKING order="4" place="4" resultid="3846" />
                    <RANKING order="5" place="-1" resultid="4431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1840" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4648" />
                    <RANKING order="2" place="2" resultid="5772" />
                    <RANKING order="3" place="3" resultid="2578" />
                    <RANKING order="4" place="4" resultid="4317" />
                    <RANKING order="5" place="5" resultid="4474" />
                    <RANKING order="6" place="6" resultid="4513" />
                    <RANKING order="7" place="7" resultid="4693" />
                    <RANKING order="8" place="-1" resultid="6758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1841" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9037" />
                    <RANKING order="2" place="2" resultid="2259" />
                    <RANKING order="3" place="3" resultid="4400" />
                    <RANKING order="4" place="4" resultid="2772" />
                    <RANKING order="5" place="5" resultid="2826" />
                    <RANKING order="6" place="6" resultid="4290" />
                    <RANKING order="7" place="7" resultid="6679" />
                    <RANKING order="8" place="8" resultid="4519" />
                    <RANKING order="9" place="-1" resultid="2703" />
                    <RANKING order="10" place="-1" resultid="4555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1842" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3263" />
                    <RANKING order="2" place="2" resultid="4364" />
                    <RANKING order="3" place="3" resultid="4388" />
                    <RANKING order="4" place="4" resultid="5647" />
                    <RANKING order="5" place="5" resultid="3740" />
                    <RANKING order="6" place="6" resultid="3808" />
                    <RANKING order="7" place="7" resultid="2370" />
                    <RANKING order="8" place="8" resultid="2821" />
                    <RANKING order="9" place="9" resultid="8053" />
                    <RANKING order="10" place="10" resultid="5728" />
                    <RANKING order="11" place="11" resultid="4689" />
                    <RANKING order="12" place="-1" resultid="4508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1843" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2601" />
                    <RANKING order="2" place="2" resultid="5987" />
                    <RANKING order="3" place="3" resultid="3233" />
                    <RANKING order="4" place="4" resultid="5930" />
                    <RANKING order="5" place="5" resultid="5940" />
                    <RANKING order="6" place="6" resultid="3763" />
                    <RANKING order="7" place="7" resultid="9047" />
                    <RANKING order="8" place="-1" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1844" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2503" />
                    <RANKING order="2" place="2" resultid="2833" />
                    <RANKING order="3" place="3" resultid="6698" />
                    <RANKING order="4" place="4" resultid="7696" />
                    <RANKING order="5" place="5" resultid="3794" />
                    <RANKING order="6" place="6" resultid="2799" />
                    <RANKING order="7" place="7" resultid="7685" />
                    <RANKING order="8" place="8" resultid="4639" />
                    <RANKING order="9" place="9" resultid="3557" />
                    <RANKING order="10" place="10" resultid="5710" />
                    <RANKING order="11" place="11" resultid="5838" />
                    <RANKING order="12" place="12" resultid="3173" />
                    <RANKING order="13" place="13" resultid="6690" />
                    <RANKING order="14" place="-1" resultid="6754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1845" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6667" />
                    <RANKING order="2" place="2" resultid="2807" />
                    <RANKING order="3" place="3" resultid="2381" />
                    <RANKING order="4" place="4" resultid="3771" />
                    <RANKING order="5" place="5" resultid="9040" />
                    <RANKING order="6" place="6" resultid="3166" />
                    <RANKING order="7" place="7" resultid="3139" />
                    <RANKING order="8" place="8" resultid="6718" />
                    <RANKING order="9" place="-1" resultid="5715" />
                    <RANKING order="10" place="-1" resultid="5822" />
                    <RANKING order="11" place="-1" resultid="6007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1846" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2778" />
                    <RANKING order="2" place="2" resultid="8172" />
                    <RANKING order="3" place="3" resultid="3239" />
                    <RANKING order="4" place="4" resultid="3851" />
                    <RANKING order="5" place="-1" resultid="2189" />
                    <RANKING order="6" place="-1" resultid="4548" />
                    <RANKING order="7" place="-1" resultid="4701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1847" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6713" />
                    <RANKING order="2" place="2" resultid="8166" />
                    <RANKING order="3" place="3" resultid="4414" />
                    <RANKING order="4" place="4" resultid="5039" />
                    <RANKING order="5" place="5" resultid="4631" />
                    <RANKING order="6" place="6" resultid="3568" />
                    <RANKING order="7" place="7" resultid="2647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1848" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2265" />
                    <RANKING order="2" place="2" resultid="4598" />
                    <RANKING order="3" place="3" resultid="7719" />
                    <RANKING order="4" place="4" resultid="6686" />
                    <RANKING order="5" place="5" resultid="2593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1849" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2664" />
                    <RANKING order="2" place="2" resultid="5024" />
                    <RANKING order="3" place="3" resultid="2624" />
                    <RANKING order="4" place="4" resultid="5755" />
                    <RANKING order="5" place="5" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1850" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1851" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2756" />
                    <RANKING order="2" place="2" resultid="8146" />
                    <RANKING order="3" place="3" resultid="2566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1852" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1853" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10147" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10148" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10149" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10150" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10151" daytime="09:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10152" daytime="09:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10153" daytime="09:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10154" daytime="09:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10155" daytime="09:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10156" daytime="09:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10157" daytime="09:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10158" daytime="09:55" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1244" daytime="09:55" gender="F" number="12" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1340" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1341" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6771" />
                    <RANKING order="2" place="2" resultid="4323" />
                    <RANKING order="3" place="-1" resultid="4573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10159" daytime="09:55" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="10:00" gender="M" number="13" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1346" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1347" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4324" />
                    <RANKING order="2" place="-1" resultid="4571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3819" />
                    <RANKING order="2" place="2" resultid="4428" />
                    <RANKING order="3" place="3" resultid="6772" />
                    <RANKING order="4" place="4" resultid="5897" />
                    <RANKING order="5" place="5" resultid="4326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5899" />
                    <RANKING order="2" place="2" resultid="4677" />
                    <RANKING order="3" place="3" resultid="3820" />
                    <RANKING order="4" place="4" resultid="3147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2724" />
                    <RANKING order="2" place="2" resultid="2725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10160" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10161" daytime="10:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1276" daytime="10:05" gender="F" number="14" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1854" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1855" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1856" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1857" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1858" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1859" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1860" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1861" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5780" />
                    <RANKING order="2" place="2" resultid="9031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1862" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1863" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1864" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1865" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1866" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1867" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1868" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10162" daytime="10:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1292" daytime="10:10" gender="M" number="15" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1869" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1870" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2349" />
                    <RANKING order="2" place="2" resultid="2356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1871" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1872" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1873" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3747" />
                    <RANKING order="2" place="2" resultid="5861" />
                    <RANKING order="3" place="3" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1874" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2209" />
                    <RANKING order="2" place="2" resultid="5723" />
                    <RANKING order="3" place="3" resultid="6014" />
                    <RANKING order="4" place="-1" resultid="3795" />
                    <RANKING order="5" place="-1" resultid="7680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1875" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2793" />
                    <RANKING order="2" place="2" resultid="3772" />
                    <RANKING order="3" place="3" resultid="3120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1876" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5633" />
                    <RANKING order="2" place="2" resultid="2329" />
                    <RANKING order="3" place="3" resultid="4655" />
                    <RANKING order="4" place="4" resultid="5981" />
                    <RANKING order="5" place="5" resultid="3197" />
                    <RANKING order="6" place="-1" resultid="3127" />
                    <RANKING order="7" place="-1" resultid="8173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1877" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4632" />
                    <RANKING order="2" place="2" resultid="3188" />
                    <RANKING order="3" place="3" resultid="3583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1878" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2266" />
                    <RANKING order="2" place="2" resultid="3081" />
                    <RANKING order="3" place="-1" resultid="7720" />
                    <RANKING order="4" place="-1" resultid="4599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1879" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1880" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1881" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1882" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1883" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10163" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10164" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10165" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10166" daytime="10:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1308" daytime="10:30" gender="F" number="16" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1884" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2317" />
                    <RANKING order="2" place="2" resultid="2491" />
                    <RANKING order="3" place="3" resultid="4374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1885" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5767" />
                    <RANKING order="2" place="2" resultid="6672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1886" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4498" />
                    <RANKING order="2" place="2" resultid="4303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1887" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1888" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2678" />
                    <RANKING order="2" place="2" resultid="3868" />
                    <RANKING order="3" place="3" resultid="5883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1889" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6745" />
                    <RANKING order="2" place="2" resultid="5654" />
                    <RANKING order="3" place="3" resultid="3787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1890" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5833" />
                    <RANKING order="2" place="2" resultid="3114" />
                    <RANKING order="3" place="3" resultid="9025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1891" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4998" />
                    <RANKING order="2" place="2" resultid="2607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1892" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1893" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1894" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1895" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1896" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1897" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1898" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10167" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10168" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10169" daytime="10:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="10:45" gender="M" number="17" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1899" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2632" />
                    <RANKING order="2" place="2" resultid="4432" />
                    <RANKING order="3" place="3" resultid="7958" />
                    <RANKING order="4" place="-1" resultid="5867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1900" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6749" />
                    <RANKING order="2" place="2" resultid="2579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1901" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4401" />
                    <RANKING order="2" place="2" resultid="5661" />
                    <RANKING order="3" place="3" resultid="4520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1902" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4365" />
                    <RANKING order="2" place="2" resultid="3802" />
                    <RANKING order="3" place="3" resultid="3809" />
                    <RANKING order="4" place="4" resultid="5959" />
                    <RANKING order="5" place="5" resultid="4311" />
                    <RANKING order="6" place="-1" resultid="3816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1903" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3256" />
                    <RANKING order="2" place="2" resultid="5988" />
                    <RANKING order="3" place="3" resultid="5931" />
                    <RANKING order="4" place="4" resultid="5995" />
                    <RANKING order="5" place="5" resultid="3159" />
                    <RANKING order="6" place="6" resultid="2484" />
                    <RANKING order="7" place="7" resultid="3764" />
                    <RANKING order="8" place="8" resultid="4280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1904" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2504" />
                    <RANKING order="2" place="2" resultid="7697" />
                    <RANKING order="3" place="3" resultid="5677" />
                    <RANKING order="4" place="4" resultid="7686" />
                    <RANKING order="5" place="5" resultid="6691" />
                    <RANKING order="6" place="6" resultid="3558" />
                    <RANKING order="7" place="7" resultid="3174" />
                    <RANKING order="8" place="8" resultid="5839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1905" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4626" />
                    <RANKING order="2" place="2" resultid="2813" />
                    <RANKING order="3" place="3" resultid="9041" />
                    <RANKING order="4" place="-1" resultid="5716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1906" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                    <RANKING order="2" place="2" resultid="2330" />
                    <RANKING order="3" place="3" resultid="3779" />
                    <RANKING order="4" place="4" resultid="6001" />
                    <RANKING order="5" place="5" resultid="3860" />
                    <RANKING order="6" place="6" resultid="3852" />
                    <RANKING order="7" place="7" resultid="5686" />
                    <RANKING order="8" place="-1" resultid="4702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1907" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5954" />
                    <RANKING order="2" place="2" resultid="2479" />
                    <RANKING order="3" place="3" resultid="4408" />
                    <RANKING order="4" place="4" resultid="3225" />
                    <RANKING order="5" place="5" resultid="3755" />
                    <RANKING order="6" place="6" resultid="3189" />
                    <RANKING order="7" place="7" resultid="3584" />
                    <RANKING order="8" place="8" resultid="4356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1908" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3088" />
                    <RANKING order="2" place="2" resultid="2594" />
                    <RANKING order="3" place="-1" resultid="4600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1909" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2642" />
                    <RANKING order="2" place="2" resultid="3218" />
                    <RANKING order="3" place="3" resultid="2625" />
                    <RANKING order="4" place="4" resultid="5947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1910" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3211" />
                    <RANKING order="2" place="2" resultid="6728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1911" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1912" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1913" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10170" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10171" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10172" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10173" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10174" daytime="11:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10175" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10176" daytime="11:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10177" daytime="11:15" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2013-06-15" daytime="16:00" name="3 Blok" number="3" warmupfrom="14:40" warmupuntil="15:40">
          <EVENTS>
            <EVENT eventid="1352" daytime="16:00" gender="F" number="18" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1914" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2318" />
                    <RANKING order="2" place="2" resultid="2492" />
                    <RANKING order="3" place="3" resultid="7714" />
                    <RANKING order="4" place="4" resultid="5744" />
                    <RANKING order="5" place="5" resultid="5874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1915" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4423" />
                    <RANKING order="2" place="2" resultid="8155" />
                    <RANKING order="3" place="3" resultid="5768" />
                    <RANKING order="4" place="4" resultid="6673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1916" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4499" />
                    <RANKING order="2" place="2" resultid="4304" />
                    <RANKING order="3" place="3" resultid="3271" />
                    <RANKING order="4" place="4" resultid="4534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1917" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1918" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1919" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6746" />
                    <RANKING order="2" place="2" resultid="5763" />
                    <RANKING order="3" place="3" resultid="3788" />
                    <RANKING order="4" place="4" resultid="5032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1920" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3115" />
                    <RANKING order="2" place="2" resultid="9026" />
                    <RANKING order="3" place="-1" resultid="5834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1921" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4999" />
                    <RANKING order="2" place="2" resultid="9032" />
                    <RANKING order="3" place="3" resultid="4610" />
                    <RANKING order="4" place="4" resultid="4307" />
                    <RANKING order="5" place="5" resultid="7705" />
                    <RANKING order="6" place="-1" resultid="2608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1922" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5005" />
                    <RANKING order="2" place="2" resultid="2614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1923" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1924" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1925" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1926" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1927" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1928" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10178" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10179" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10180" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10181" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10182" daytime="16:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1369" daytime="16:10" gender="M" number="19" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1929" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2633" />
                    <RANKING order="2" place="2" resultid="7959" />
                    <RANKING order="3" place="3" resultid="4433" />
                    <RANKING order="4" place="-1" resultid="5868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1930" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6750" />
                    <RANKING order="2" place="2" resultid="2324" />
                    <RANKING order="3" place="3" resultid="2580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1931" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5662" />
                    <RANKING order="2" place="2" resultid="9471" />
                    <RANKING order="3" place="3" resultid="4521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1932" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3810" />
                    <RANKING order="2" place="2" resultid="3803" />
                    <RANKING order="3" place="3" resultid="7947" />
                    <RANKING order="4" place="4" resultid="5648" />
                    <RANKING order="5" place="5" resultid="3817" />
                    <RANKING order="6" place="6" resultid="4674" />
                    <RANKING order="7" place="7" resultid="4312" />
                    <RANKING order="8" place="8" resultid="4366" />
                    <RANKING order="9" place="-1" resultid="6766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1933" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3257" />
                    <RANKING order="2" place="2" resultid="5996" />
                    <RANKING order="3" place="3" resultid="3748" />
                    <RANKING order="4" place="4" resultid="5932" />
                    <RANKING order="5" place="5" resultid="5989" />
                    <RANKING order="6" place="6" resultid="3160" />
                    <RANKING order="7" place="7" resultid="9048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1934" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2505" />
                    <RANKING order="2" place="2" resultid="7698" />
                    <RANKING order="3" place="3" resultid="5678" />
                    <RANKING order="4" place="4" resultid="5711" />
                    <RANKING order="5" place="5" resultid="6692" />
                    <RANKING order="6" place="6" resultid="3559" />
                    <RANKING order="7" place="7" resultid="3175" />
                    <RANKING order="8" place="-1" resultid="6755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1935" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2382" />
                    <RANKING order="2" place="2" resultid="4627" />
                    <RANKING order="3" place="3" resultid="2814" />
                    <RANKING order="4" place="4" resultid="5823" />
                    <RANKING order="5" place="5" resultid="3140" />
                    <RANKING order="6" place="6" resultid="5717" />
                    <RANKING order="7" place="7" resultid="2804" />
                    <RANKING order="8" place="-1" resultid="4492" />
                    <RANKING order="9" place="-1" resultid="6008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1936" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6002" />
                    <RANKING order="2" place="2" resultid="2331" />
                    <RANKING order="3" place="3" resultid="3780" />
                    <RANKING order="4" place="4" resultid="3099" />
                    <RANKING order="5" place="5" resultid="3861" />
                    <RANKING order="6" place="6" resultid="3853" />
                    <RANKING order="7" place="7" resultid="2588" />
                    <RANKING order="8" place="8" resultid="5685" />
                    <RANKING order="9" place="9" resultid="3198" />
                    <RANKING order="10" place="-1" resultid="4549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1937" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5955" />
                    <RANKING order="2" place="2" resultid="2480" />
                    <RANKING order="3" place="3" resultid="4409" />
                    <RANKING order="4" place="4" resultid="4415" />
                    <RANKING order="5" place="5" resultid="3226" />
                    <RANKING order="6" place="6" resultid="4357" />
                    <RANKING order="7" place="-1" resultid="2768" />
                    <RANKING order="8" place="-1" resultid="8163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1938" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3089" />
                    <RANKING order="2" place="2" resultid="2267" />
                    <RANKING order="3" place="3" resultid="6687" />
                    <RANKING order="4" place="-1" resultid="4601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1939" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3219" />
                    <RANKING order="2" place="2" resultid="5948" />
                    <RANKING order="3" place="3" resultid="2626" />
                    <RANKING order="4" place="4" resultid="2643" />
                    <RANKING order="5" place="5" resultid="3576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1940" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3212" />
                    <RANKING order="2" place="2" resultid="6729" />
                    <RANKING order="3" place="3" resultid="5048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1941" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1942" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1943" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10183" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10184" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10185" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10186" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10187" daytime="16:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10188" daytime="16:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10189" daytime="16:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10190" daytime="16:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10191" daytime="16:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10192" daytime="16:20" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1385" daytime="16:20" gender="F" number="20" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1944" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2732" />
                    <RANKING order="2" place="2" resultid="2765" />
                    <RANKING order="3" place="3" resultid="5846" />
                    <RANKING order="4" place="4" resultid="5852" />
                    <RANKING order="5" place="5" resultid="2493" />
                    <RANKING order="6" place="6" resultid="4375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1945" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8156" />
                    <RANKING order="2" place="2" resultid="5816" />
                    <RANKING order="3" place="3" resultid="7970" />
                    <RANKING order="4" place="4" resultid="8180" />
                    <RANKING order="5" place="-1" resultid="2574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1946" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4394" />
                    <RANKING order="2" place="2" resultid="3272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1947" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6722" />
                    <RANKING order="2" place="2" resultid="4563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1948" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3136" />
                    <RANKING order="2" place="2" resultid="5736" />
                    <RANKING order="3" place="3" resultid="4542" />
                    <RANKING order="4" place="4" resultid="5885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1949" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6021" />
                    <RANKING order="2" place="2" resultid="2787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1950" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5974" />
                    <RANKING order="2" place="2" resultid="3109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1951" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5000" />
                    <RANKING order="2" place="2" resultid="2374" />
                    <RANKING order="3" place="3" resultid="5781" />
                    <RANKING order="4" place="4" resultid="3104" />
                    <RANKING order="5" place="5" resultid="4614" />
                    <RANKING order="6" place="6" resultid="2609" />
                    <RANKING order="7" place="7" resultid="7706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1952" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2696" />
                    <RANKING order="2" place="2" resultid="2615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1953" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4504" />
                    <RANKING order="2" place="2" resultid="4589" />
                    <RANKING order="3" place="3" resultid="5808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1954" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1955" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6739" />
                    <RANKING order="2" place="2" resultid="4669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1956" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1957" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1958" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10193" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10194" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10195" daytime="16:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10196" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10197" daytime="16:30" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1401" daytime="16:30" gender="M" number="21" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1959" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1960" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2556" />
                    <RANKING order="2" place="2" resultid="4649" />
                    <RANKING order="3" place="3" resultid="4485" />
                    <RANKING order="4" place="4" resultid="6759" />
                    <RANKING order="5" place="5" resultid="2358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1961" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4402" />
                    <RANKING order="2" place="2" resultid="5663" />
                    <RANKING order="3" place="3" resultid="6680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1962" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3741" />
                    <RANKING order="2" place="2" resultid="4389" />
                    <RANKING order="3" place="3" resultid="2250" />
                    <RANKING order="4" place="4" resultid="4276" />
                    <RANKING order="5" place="5" resultid="5829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1963" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="3828" />
                    <RANKING order="3" place="3" resultid="2602" />
                    <RANKING order="4" place="4" resultid="2254" />
                    <RANKING order="5" place="5" resultid="5941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1964" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6699" />
                    <RANKING order="2" place="2" resultid="2338" />
                    <RANKING order="3" place="3" resultid="2800" />
                    <RANKING order="4" place="4" resultid="5724" />
                    <RANKING order="5" place="5" resultid="3796" />
                    <RANKING order="6" place="6" resultid="5679" />
                    <RANKING order="7" place="7" resultid="4640" />
                    <RANKING order="8" place="8" resultid="6015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1965" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4493" />
                    <RANKING order="2" place="2" resultid="2383" />
                    <RANKING order="3" place="3" resultid="5824" />
                    <RANKING order="4" place="4" resultid="9042" />
                    <RANKING order="5" place="5" resultid="3167" />
                    <RANKING order="6" place="-1" resultid="7954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1966" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5634" />
                    <RANKING order="2" place="2" resultid="4619" />
                    <RANKING order="3" place="3" resultid="10303" />
                    <RANKING order="4" place="4" resultid="3183" />
                    <RANKING order="5" place="5" resultid="8174" />
                    <RANKING order="6" place="-1" resultid="2760" />
                    <RANKING order="7" place="-1" resultid="3128" />
                    <RANKING order="8" place="-1" resultid="4550" />
                    <RANKING order="9" place="-1" resultid="4703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1967" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6714" />
                    <RANKING order="2" place="2" resultid="8165" />
                    <RANKING order="3" place="3" resultid="5040" />
                    <RANKING order="4" place="4" resultid="3094" />
                    <RANKING order="5" place="5" resultid="3756" />
                    <RANKING order="6" place="6" resultid="3569" />
                    <RANKING order="7" place="7" resultid="4358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1968" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4602" />
                    <RANKING order="2" place="2" resultid="2658" />
                    <RANKING order="3" place="3" resultid="3082" />
                    <RANKING order="4" place="4" resultid="2712" />
                    <RANKING order="5" place="5" resultid="2595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1969" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2665" />
                    <RANKING order="2" place="2" resultid="5025" />
                    <RANKING order="3" place="3" resultid="3249" />
                    <RANKING order="4" place="4" resultid="5756" />
                    <RANKING order="5" place="5" resultid="3577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1970" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5049" />
                    <RANKING order="2" place="2" resultid="6730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1971" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8147" />
                    <RANKING order="2" place="2" resultid="2567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1972" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1973" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10198" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10199" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10200" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10201" daytime="16:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10202" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10203" daytime="16:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10204" daytime="16:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10205" daytime="16:50" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1417" daytime="16:50" gender="F" number="22" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1513" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1514" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6773" />
                    <RANKING order="2" place="-1" resultid="4574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5904" />
                    <RANKING order="2" place="2" resultid="4322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10206" daytime="16:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1433" daytime="16:55" gender="M" number="23" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1519" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1520" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4325" />
                    <RANKING order="2" place="2" resultid="6774" />
                    <RANKING order="3" place="-1" resultid="4572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3821" />
                    <RANKING order="2" place="2" resultid="4429" />
                    <RANKING order="3" place="3" resultid="5898" />
                    <RANKING order="4" place="4" resultid="4327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4678" />
                    <RANKING order="2" place="2" resultid="3822" />
                    <RANKING order="3" place="3" resultid="5900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1524" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10207" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10208" daytime="16:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1449" daytime="17:00" gender="F" number="24" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1975" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5875" />
                    <RANKING order="2" place="2" resultid="5853" />
                    <RANKING order="3" place="3" resultid="5750" />
                    <RANKING order="4" place="4" resultid="4376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1976" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                    <RANKING order="2" place="2" resultid="2519" />
                    <RANKING order="3" place="3" resultid="2747" />
                    <RANKING order="4" place="4" resultid="6674" />
                    <RANKING order="5" place="5" resultid="2575" />
                    <RANKING order="6" place="6" resultid="6708" />
                    <RANKING order="7" place="7" resultid="7692" />
                    <RANKING order="8" place="8" resultid="4528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1977" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6030" />
                    <RANKING order="2" place="2" resultid="4395" />
                    <RANKING order="3" place="3" resultid="5641" />
                    <RANKING order="4" place="4" resultid="6735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1978" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6723" />
                    <RANKING order="2" place="2" resultid="4564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1979" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4543" />
                    <RANKING order="2" place="2" resultid="3869" />
                    <RANKING order="3" place="3" resultid="4285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1980" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2366" />
                    <RANKING order="2" place="2" resultid="6747" />
                    <RANKING order="3" place="3" resultid="6022" />
                    <RANKING order="4" place="4" resultid="2788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1981" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3206" />
                    <RANKING order="2" place="2" resultid="6026" />
                    <RANKING order="3" place="3" resultid="3842" />
                    <RANKING order="4" place="4" resultid="9027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1982" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9033" />
                    <RANKING order="2" place="2" resultid="4615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1983" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1984" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1985" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1986" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1987" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1988" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1989" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10209" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10210" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10211" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10212" daytime="17:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10213" daytime="17:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1465" daytime="17:20" gender="M" number="25" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1990" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5624" />
                    <RANKING order="2" place="2" resultid="4479" />
                    <RANKING order="3" place="3" resultid="3847" />
                    <RANKING order="4" place="4" resultid="4434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1991" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4650" />
                    <RANKING order="2" place="2" resultid="2350" />
                    <RANKING order="3" place="3" resultid="5773" />
                    <RANKING order="4" place="-1" resultid="4694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1992" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2771" />
                    <RANKING order="2" place="2" resultid="2827" />
                    <RANKING order="3" place="3" resultid="4556" />
                    <RANKING order="4" place="4" resultid="4291" />
                    <RANKING order="5" place="5" resultid="4383" />
                    <RANKING order="6" place="6" resultid="6681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1993" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3264" />
                    <RANKING order="2" place="2" resultid="2371" />
                    <RANKING order="3" place="3" resultid="3811" />
                    <RANKING order="4" place="4" resultid="2822" />
                    <RANKING order="5" place="5" resultid="5729" />
                    <RANKING order="6" place="6" resultid="8054" />
                    <RANKING order="7" place="-1" resultid="4509" />
                    <RANKING order="8" place="-1" resultid="4690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1994" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5990" />
                    <RANKING order="2" place="2" resultid="3234" />
                    <RANKING order="3" place="3" resultid="5933" />
                    <RANKING order="4" place="4" resultid="3765" />
                    <RANKING order="5" place="5" resultid="5942" />
                    <RANKING order="6" place="6" resultid="6742" />
                    <RANKING order="7" place="-1" resultid="3829" />
                    <RANKING order="8" place="-1" resultid="4281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1995" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2506" />
                    <RANKING order="2" place="2" resultid="7681" />
                    <RANKING order="3" place="3" resultid="2834" />
                    <RANKING order="4" place="4" resultid="7687" />
                    <RANKING order="5" place="5" resultid="6700" />
                    <RANKING order="6" place="6" resultid="3797" />
                    <RANKING order="7" place="7" resultid="4641" />
                    <RANKING order="8" place="8" resultid="5840" />
                    <RANKING order="9" place="9" resultid="3560" />
                    <RANKING order="10" place="10" resultid="3176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1996" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6668" />
                    <RANKING order="2" place="2" resultid="2808" />
                    <RANKING order="3" place="3" resultid="3773" />
                    <RANKING order="4" place="4" resultid="2794" />
                    <RANKING order="5" place="5" resultid="9043" />
                    <RANKING order="6" place="6" resultid="5718" />
                    <RANKING order="7" place="7" resultid="6719" />
                    <RANKING order="8" place="-1" resultid="3168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1997" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3129" />
                    <RANKING order="2" place="2" resultid="6003" />
                    <RANKING order="3" place="3" resultid="2779" />
                    <RANKING order="4" place="4" resultid="5982" />
                    <RANKING order="5" place="5" resultid="3240" />
                    <RANKING order="6" place="6" resultid="3862" />
                    <RANKING order="7" place="-1" resultid="2190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1998" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6715" />
                    <RANKING order="2" place="2" resultid="8167" />
                    <RANKING order="3" place="3" resultid="5041" />
                    <RANKING order="4" place="4" resultid="4633" />
                    <RANKING order="5" place="5" resultid="3190" />
                    <RANKING order="6" place="6" resultid="3585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1999" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4603" />
                    <RANKING order="2" place="2" resultid="7721" />
                    <RANKING order="3" place="3" resultid="2596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2000" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2666" />
                    <RANKING order="2" place="2" resultid="3220" />
                    <RANKING order="3" place="3" resultid="5026" />
                    <RANKING order="4" place="4" resultid="5757" />
                    <RANKING order="5" place="5" resultid="5949" />
                    <RANKING order="6" place="6" resultid="2627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2001" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2002" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8148" />
                    <RANKING order="2" place="2" resultid="2568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2003" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2004" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10214" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10215" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10216" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10217" daytime="17:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10218" daytime="17:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10219" daytime="17:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10220" daytime="17:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10221" daytime="17:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10222" daytime="17:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10223" daytime="17:55" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1481" daytime="17:55" gender="F" number="26" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2005" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2006" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2007" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="2008" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="2009" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2679" />
                    <RANKING order="2" place="2" resultid="5737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2010" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5655" />
                    <RANKING order="2" place="2" resultid="3789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2011" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2012" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2013" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                    <RANKING order="2" place="2" resultid="5006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2014" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="2015" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="2016" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="2017" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2018" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2019" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10224" daytime="17:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10225" daytime="18:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1497" daytime="18:15" gender="M" number="27" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2020" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2021" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2351" />
                    <RANKING order="2" place="2" resultid="4318" />
                    <RANKING order="3" place="3" resultid="2359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2022" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4403" />
                    <RANKING order="2" place="2" resultid="4297" />
                    <RANKING order="3" place="3" resultid="4384" />
                    <RANKING order="4" place="4" resultid="4522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2023" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3804" />
                    <RANKING order="2" place="2" resultid="3818" />
                    <RANKING order="3" place="-1" resultid="4367" />
                    <RANKING order="4" place="-1" resultid="6767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2024" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3749" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="5862" />
                    <RANKING order="4" place="4" resultid="3766" />
                    <RANKING order="5" place="5" resultid="9054" />
                    <RANKING order="6" place="-1" resultid="2485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2025" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="2211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2026" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3774" />
                    <RANKING order="2" place="2" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2027" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4620" />
                    <RANKING order="2" place="2" resultid="2332" />
                    <RANKING order="3" place="3" resultid="5017" />
                    <RANKING order="4" place="4" resultid="3854" />
                    <RANKING order="5" place="-1" resultid="4704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2028" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5956" />
                    <RANKING order="2" place="2" resultid="3570" />
                    <RANKING order="3" place="3" resultid="3757" />
                    <RANKING order="4" place="4" resultid="4416" />
                    <RANKING order="5" place="5" resultid="3095" />
                    <RANKING order="6" place="6" resultid="3227" />
                    <RANKING order="7" place="7" resultid="3191" />
                    <RANKING order="8" place="8" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2029" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2268" />
                    <RANKING order="2" place="2" resultid="7722" />
                    <RANKING order="3" place="3" resultid="3083" />
                    <RANKING order="4" place="-1" resultid="4604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2030" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2031" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="2032" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2033" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2034" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10226" daytime="18:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10227" daytime="18:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10228" daytime="18:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10229" daytime="18:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10230" daytime="18:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10231" daytime="18:55" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2013-06-16" daytime="09:00" name="4 Blok" number="4" warmupfrom="07:40" warmupuntil="08:40">
          <EVENTS>
            <EVENT eventid="1525" daytime="09:00" gender="F" number="28" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2035" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5745" />
                    <RANKING order="2" place="2" resultid="5876" />
                    <RANKING order="3" place="-1" resultid="5880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2036" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6675" />
                    <RANKING order="2" place="2" resultid="6710" />
                    <RANKING order="3" place="3" resultid="4529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2037" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3273" />
                    <RANKING order="2" place="2" resultid="5642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2038" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2039" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2040" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2041" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2042" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2043" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="2044" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="2045" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2046" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="2047" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2048" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2049" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10232" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10233" daytime="09:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1542" daytime="09:05" gender="M" number="29" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2050" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4480" />
                    <RANKING order="2" place="2" resultid="5626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2051" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4651" />
                    <RANKING order="2" place="2" resultid="2360" />
                    <RANKING order="3" place="3" resultid="8142" />
                    <RANKING order="4" place="4" resultid="4514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2052" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9038" />
                    <RANKING order="2" place="2" resultid="4271" />
                    <RANKING order="3" place="3" resultid="2828" />
                    <RANKING order="4" place="4" resultid="4292" />
                    <RANKING order="5" place="5" resultid="4385" />
                    <RANKING order="6" place="6" resultid="4523" />
                    <RANKING order="7" place="-1" resultid="4557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2053" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2251" />
                    <RANKING order="2" place="2" resultid="2823" />
                    <RANKING order="3" place="-1" resultid="4368" />
                    <RANKING order="4" place="-1" resultid="6768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2054" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3750" />
                    <RANKING order="2" place="2" resultid="2603" />
                    <RANKING order="3" place="3" resultid="2639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2055" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2212" />
                    <RANKING order="2" place="2" resultid="7682" />
                    <RANKING order="3" place="3" resultid="5725" />
                    <RANKING order="4" place="4" resultid="3561" />
                    <RANKING order="5" place="-1" resultid="6016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2056" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2795" />
                    <RANKING order="2" place="2" resultid="5670" />
                    <RANKING order="3" place="3" resultid="3122" />
                    <RANKING order="4" place="-1" resultid="5825" />
                    <RANKING order="5" place="-1" resultid="6009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2057" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5635" />
                    <RANKING order="2" place="2" resultid="4656" />
                    <RANKING order="3" place="3" resultid="2333" />
                    <RANKING order="4" place="4" resultid="5983" />
                    <RANKING order="5" place="5" resultid="3184" />
                    <RANKING order="6" place="6" resultid="3855" />
                    <RANKING order="7" place="-1" resultid="3130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2058" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4417" />
                    <RANKING order="2" place="2" resultid="4634" />
                    <RANKING order="3" place="3" resultid="3571" />
                    <RANKING order="4" place="4" resultid="3587" />
                    <RANKING order="5" place="-1" resultid="4359" />
                    <RANKING order="6" place="-1" resultid="8168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2059" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2269" />
                    <RANKING order="2" place="2" resultid="7723" />
                    <RANKING order="3" place="3" resultid="3084" />
                    <RANKING order="4" place="4" resultid="2597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2060" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2061" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2198" />
                    <RANKING order="2" place="2" resultid="6731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2062" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2063" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2064" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10234" daytime="09:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10235" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10236" daytime="09:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10237" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10238" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10239" daytime="09:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10240" daytime="09:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1558" daytime="09:20" gender="F" number="30" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2065" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2320" />
                    <RANKING order="2" place="2" resultid="5847" />
                    <RANKING order="3" place="3" resultid="5751" />
                    <RANKING order="4" place="4" resultid="2494" />
                    <RANKING order="5" place="5" resultid="5746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2066" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4424" />
                    <RANKING order="2" place="2" resultid="8157" />
                    <RANKING order="3" place="3" resultid="4472" />
                    <RANKING order="4" place="-1" resultid="2520" />
                    <RANKING order="5" place="-1" resultid="2576" />
                    <RANKING order="6" place="-1" resultid="7693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2067" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9053" />
                    <RANKING order="2" place="2" resultid="4268" />
                    <RANKING order="3" place="3" resultid="4535" />
                    <RANKING order="4" place="4" resultid="6736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2068" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2069" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3870" />
                    <RANKING order="2" place="2" resultid="4286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2070" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5764" />
                    <RANKING order="2" place="2" resultid="6023" />
                    <RANKING order="3" place="3" resultid="5656" />
                    <RANKING order="4" place="4" resultid="5033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2071" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3116" />
                    <RANKING order="2" place="2" resultid="3207" />
                    <RANKING order="3" place="3" resultid="3843" />
                    <RANKING order="4" place="4" resultid="6027" />
                    <RANKING order="5" place="5" resultid="9028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2072" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5783" />
                    <RANKING order="2" place="2" resultid="3105" />
                    <RANKING order="3" place="3" resultid="4611" />
                    <RANKING order="4" place="4" resultid="4308" />
                    <RANKING order="5" place="5" resultid="7707" />
                    <RANKING order="6" place="6" resultid="2610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2073" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5007" />
                    <RANKING order="2" place="2" resultid="2686" />
                    <RANKING order="3" place="3" resultid="2616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2074" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2718" />
                    <RANKING order="2" place="2" resultid="4505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2075" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2076" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="2077" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2078" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2079" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10241" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10242" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10243" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10244" daytime="09:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10245" daytime="09:25" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1574" daytime="09:25" gender="M" number="31" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2080" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5627" />
                    <RANKING order="2" place="2" resultid="4481" />
                    <RANKING order="3" place="3" resultid="4435" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="-1" resultid="7960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2081" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5774" />
                    <RANKING order="2" place="2" resultid="6760" />
                    <RANKING order="3" place="3" resultid="2325" />
                    <RANKING order="4" place="4" resultid="2581" />
                    <RANKING order="5" place="5" resultid="4475" />
                    <RANKING order="6" place="6" resultid="4515" />
                    <RANKING order="7" place="7" resultid="4695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2082" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2260" />
                    <RANKING order="2" place="2" resultid="9039" />
                    <RANKING order="3" place="3" resultid="2773" />
                    <RANKING order="4" place="4" resultid="6682" />
                    <RANKING order="5" place="5" resultid="2704" />
                    <RANKING order="6" place="-1" resultid="2829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2083" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3742" />
                    <RANKING order="2" place="2" resultid="5649" />
                    <RANKING order="3" place="3" resultid="3265" />
                    <RANKING order="4" place="4" resultid="8185" />
                    <RANKING order="5" place="5" resultid="8055" />
                    <RANKING order="6" place="6" resultid="7948" />
                    <RANKING order="7" place="7" resultid="2824" />
                    <RANKING order="8" place="8" resultid="5730" />
                    <RANKING order="9" place="9" resultid="4691" />
                    <RANKING order="10" place="10" resultid="4675" />
                    <RANKING order="11" place="-1" resultid="4510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2084" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5991" />
                    <RANKING order="2" place="2" resultid="3235" />
                    <RANKING order="3" place="3" resultid="3830" />
                    <RANKING order="4" place="4" resultid="5997" />
                    <RANKING order="5" place="5" resultid="2604" />
                    <RANKING order="6" place="6" resultid="5934" />
                    <RANKING order="7" place="7" resultid="5943" />
                    <RANKING order="8" place="8" resultid="9049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2085" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="2507" />
                    <RANKING order="3" place="3" resultid="7700" />
                    <RANKING order="4" place="4" resultid="3798" />
                    <RANKING order="5" place="5" resultid="6701" />
                    <RANKING order="6" place="6" resultid="2801" />
                    <RANKING order="7" place="7" resultid="4642" />
                    <RANKING order="8" place="8" resultid="7688" />
                    <RANKING order="9" place="9" resultid="5712" />
                    <RANKING order="10" place="10" resultid="5841" />
                    <RANKING order="11" place="11" resultid="3177" />
                    <RANKING order="12" place="12" resultid="6693" />
                    <RANKING order="13" place="-1" resultid="6756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2086" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6669" />
                    <RANKING order="2" place="2" resultid="2384" />
                    <RANKING order="3" place="3" resultid="2809" />
                    <RANKING order="4" place="4" resultid="9044" />
                    <RANKING order="5" place="5" resultid="2708" />
                    <RANKING order="6" place="6" resultid="3141" />
                    <RANKING order="7" place="7" resultid="2815" />
                    <RANKING order="8" place="8" resultid="3169" />
                    <RANKING order="9" place="9" resultid="4321" />
                    <RANKING order="10" place="10" resultid="2805" />
                    <RANKING order="11" place="-1" resultid="6010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2087" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4657" />
                    <RANKING order="2" place="2" resultid="2191" />
                    <RANKING order="3" place="3" resultid="3781" />
                    <RANKING order="4" place="4" resultid="3863" />
                    <RANKING order="5" place="5" resultid="8175" />
                    <RANKING order="6" place="6" resultid="3241" />
                    <RANKING order="7" place="7" resultid="5687" />
                    <RANKING order="8" place="-1" resultid="2780" />
                    <RANKING order="9" place="-1" resultid="4551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2088" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4418" />
                    <RANKING order="2" place="2" resultid="5042" />
                    <RANKING order="3" place="3" resultid="4635" />
                    <RANKING order="4" place="-1" resultid="8164" />
                    <RANKING order="5" place="-1" resultid="2648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2089" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2701" />
                    <RANKING order="2" place="1" resultid="4605" />
                    <RANKING order="3" place="3" resultid="2270" />
                    <RANKING order="4" place="4" resultid="6688" />
                    <RANKING order="5" place="5" resultid="2713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2090" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2667" />
                    <RANKING order="2" place="2" resultid="3221" />
                    <RANKING order="3" place="3" resultid="5950" />
                    <RANKING order="4" place="4" resultid="5027" />
                    <RANKING order="5" place="5" resultid="5758" />
                    <RANKING order="6" place="6" resultid="3578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2091" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2092" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2754" />
                    <RANKING order="2" place="2" resultid="2569" />
                    <RANKING order="3" place="3" resultid="5707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2093" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2094" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10246" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10247" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10248" daytime="09:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10249" daytime="09:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10250" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10251" daytime="09:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10252" daytime="09:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10253" daytime="09:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10254" daytime="09:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10255" daytime="09:35" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10256" daytime="09:35" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10257" daytime="09:40" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1590" daytime="09:40" gender="F" number="32" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2095" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2766" />
                    <RANKING order="2" place="2" resultid="5854" />
                    <RANKING order="3" place="3" resultid="2495" />
                    <RANKING order="4" place="4" resultid="4377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2096" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5817" />
                    <RANKING order="2" place="2" resultid="7971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2097" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4396" />
                    <RANKING order="2" place="2" resultid="3274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2098" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2099" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5738" />
                    <RANKING order="2" place="2" resultid="4544" />
                    <RANKING order="3" place="3" resultid="5886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2100" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6024" />
                    <RANKING order="2" place="2" resultid="2789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2101" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5976" />
                    <RANKING order="2" place="2" resultid="9029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2102" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5001" />
                    <RANKING order="2" place="2" resultid="2375" />
                    <RANKING order="3" place="3" resultid="4616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2103" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2104" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2105" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="2106" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2107" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2108" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2109" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10258" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10259" daytime="09:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10260" daytime="09:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1606" daytime="09:55" gender="M" number="33" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2110" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2111" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4486" />
                    <RANKING order="2" place="2" resultid="2361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2112" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2113" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3743" />
                    <RANKING order="2" place="2" resultid="4390" />
                    <RANKING order="3" place="3" resultid="4277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2114" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="3767" />
                    <RANKING order="3" place="3" resultid="2255" />
                    <RANKING order="4" place="-1" resultid="3831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2115" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2339" />
                    <RANKING order="2" place="2" resultid="6702" />
                    <RANKING order="3" place="3" resultid="2802" />
                    <RANKING order="4" place="4" resultid="7701" />
                    <RANKING order="5" place="5" resultid="3799" />
                    <RANKING order="6" place="6" resultid="4643" />
                    <RANKING order="7" place="7" resultid="5681" />
                    <RANKING order="8" place="8" resultid="6017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2116" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4494" />
                    <RANKING order="2" place="2" resultid="3775" />
                    <RANKING order="3" place="3" resultid="3170" />
                    <RANKING order="4" place="-1" resultid="5826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2117" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4621" />
                    <RANKING order="2" place="2" resultid="3131" />
                    <RANKING order="3" place="3" resultid="5018" />
                    <RANKING order="4" place="4" resultid="3185" />
                    <RANKING order="5" place="-1" resultid="2761" />
                    <RANKING order="6" place="-1" resultid="4705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2118" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6716" />
                    <RANKING order="2" place="2" resultid="3758" />
                    <RANKING order="3" place="3" resultid="3096" />
                    <RANKING order="4" place="4" resultid="3192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2119" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4606" />
                    <RANKING order="2" place="2" resultid="2659" />
                    <RANKING order="3" place="3" resultid="3085" />
                    <RANKING order="4" place="4" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2120" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5028" />
                    <RANKING order="2" place="2" resultid="3252" />
                    <RANKING order="3" place="3" resultid="10310" />
                    <RANKING order="4" place="4" resultid="5759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2121" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2122" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8149" />
                    <RANKING order="2" place="2" resultid="2570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2123" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2124" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10261" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10262" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10263" daytime="10:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10264" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10265" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10266" daytime="10:15" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1622" daytime="10:20" gender="X" number="34" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1702" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2584" />
                    <RANKING order="2" place="-1" resultid="5890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4426" />
                    <RANKING order="2" place="2" resultid="4328" />
                    <RANKING order="3" place="3" resultid="6775" />
                    <RANKING order="4" place="4" resultid="5889" />
                    <RANKING order="5" place="5" resultid="8141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5893" />
                    <RANKING order="2" place="2" resultid="5666" />
                    <RANKING order="3" place="3" resultid="9050" />
                    <RANKING order="4" place="4" resultid="4330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5895" />
                    <RANKING order="2" place="2" resultid="3144" />
                    <RANKING order="3" place="3" resultid="3873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2728" />
                    <RANKING order="2" place="2" resultid="9475" />
                    <RANKING order="3" place="3" resultid="5896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2720" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10267" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10268" daytime="10:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10269" daytime="10:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1638" daytime="10:30" gender="F" number="35" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2125" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2126" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4425" />
                    <RANKING order="2" place="2" resultid="8158" />
                    <RANKING order="3" place="3" resultid="5769" />
                    <RANKING order="4" place="4" resultid="6676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2127" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4500" />
                    <RANKING order="2" place="2" resultid="4305" />
                    <RANKING order="3" place="-1" resultid="4536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2128" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2129" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2681" />
                    <RANKING order="2" place="2" resultid="5887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2130" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6748" />
                    <RANKING order="2" place="2" resultid="3791" />
                    <RANKING order="3" place="-1" resultid="5034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2131" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3117" />
                    <RANKING order="2" place="2" resultid="5835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2132" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5002" />
                    <RANKING order="2" place="2" resultid="9035" />
                    <RANKING order="3" place="3" resultid="2611" />
                    <RANKING order="4" place="4" resultid="7708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2133" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5008" />
                    <RANKING order="2" place="2" resultid="2617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2134" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2135" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2136" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2137" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="2138" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2139" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10270" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10271" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10272" daytime="10:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10273" daytime="10:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1654" daytime="10:40" gender="M" number="36" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2140" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7961" />
                    <RANKING order="2" place="2" resultid="4436" />
                    <RANKING order="3" place="-1" resultid="5869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2141" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6751" />
                    <RANKING order="2" place="2" resultid="2582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2142" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5664" />
                    <RANKING order="2" place="2" resultid="4524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2143" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3805" />
                    <RANKING order="2" place="2" resultid="3812" />
                    <RANKING order="3" place="3" resultid="7949" />
                    <RANKING order="4" place="-1" resultid="4676" />
                    <RANKING order="5" place="-1" resultid="4313" />
                    <RANKING order="6" place="-1" resultid="4369" />
                    <RANKING order="7" place="-1" resultid="6769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2144" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3751" />
                    <RANKING order="2" place="2" resultid="3259" />
                    <RANKING order="3" place="3" resultid="5935" />
                    <RANKING order="4" place="4" resultid="5998" />
                    <RANKING order="5" place="5" resultid="3161" />
                    <RANKING order="6" place="-1" resultid="2486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2145" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2508" />
                    <RANKING order="2" place="2" resultid="5688" />
                    <RANKING order="3" place="3" resultid="5713" />
                    <RANKING order="4" place="4" resultid="6694" />
                    <RANKING order="5" place="5" resultid="3178" />
                    <RANKING order="6" place="-1" resultid="6757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2146" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2385" />
                    <RANKING order="2" place="2" resultid="4495" />
                    <RANKING order="3" place="3" resultid="4628" />
                    <RANKING order="4" place="4" resultid="2816" />
                    <RANKING order="5" place="5" resultid="9045" />
                    <RANKING order="6" place="6" resultid="5719" />
                    <RANKING order="7" place="7" resultid="5671" />
                    <RANKING order="8" place="8" resultid="3142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2147" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6004" />
                    <RANKING order="2" place="2" resultid="4622" />
                    <RANKING order="3" place="3" resultid="2334" />
                    <RANKING order="4" place="4" resultid="3782" />
                    <RANKING order="5" place="5" resultid="3100" />
                    <RANKING order="6" place="6" resultid="3864" />
                    <RANKING order="7" place="7" resultid="3199" />
                    <RANKING order="8" place="8" resultid="2589" />
                    <RANKING order="9" place="-1" resultid="4552" />
                    <RANKING order="10" place="-1" resultid="4706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2148" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5957" />
                    <RANKING order="2" place="2" resultid="2481" />
                    <RANKING order="3" place="3" resultid="4410" />
                    <RANKING order="4" place="4" resultid="3228" />
                    <RANKING order="5" place="5" resultid="4360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2149" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2150" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2644" />
                    <RANKING order="2" place="2" resultid="3222" />
                    <RANKING order="3" place="3" resultid="2628" />
                    <RANKING order="4" place="4" resultid="5951" />
                    <RANKING order="5" place="5" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2151" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6732" />
                    <RANKING order="2" place="-1" resultid="3213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2152" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2153" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2154" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10274" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10275" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10276" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10277" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10278" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10279" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10280" daytime="10:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10281" daytime="11:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1670" daytime="11:00" gender="F" number="37" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2155" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5877" />
                    <RANKING order="2" place="2" resultid="5855" />
                    <RANKING order="3" place="3" resultid="4378" />
                    <RANKING order="4" place="4" resultid="7715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2156" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2245" />
                    <RANKING order="2" place="2" resultid="5818" />
                    <RANKING order="3" place="3" resultid="7694" />
                    <RANKING order="4" place="4" resultid="6711" />
                    <RANKING order="5" place="5" resultid="4530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2157" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6031" />
                    <RANKING order="2" place="2" resultid="5643" />
                    <RANKING order="3" place="3" resultid="6737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2158" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2204" />
                    <RANKING order="2" place="2" resultid="4566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2159" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3137" />
                    <RANKING order="2" place="2" resultid="5739" />
                    <RANKING order="3" place="3" resultid="4545" />
                    <RANKING order="4" place="4" resultid="3871" />
                    <RANKING order="5" place="5" resultid="4287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2160" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2367" />
                    <RANKING order="2" place="2" resultid="5657" />
                    <RANKING order="3" place="3" resultid="2790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2161" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5977" />
                    <RANKING order="2" place="2" resultid="3208" />
                    <RANKING order="3" place="3" resultid="6028" />
                    <RANKING order="4" place="4" resultid="3844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2162" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5784" />
                    <RANKING order="2" place="2" resultid="4617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2163" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="2164" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4591" />
                    <RANKING order="2" place="2" resultid="5811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2165" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="2166" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="2167" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2168" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2169" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10282" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10283" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10284" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10285" daytime="11:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1686" daytime="11:35" gender="M" number="38" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2170" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="2171" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2352" />
                    <RANKING order="2" place="2" resultid="4652" />
                    <RANKING order="3" place="3" resultid="6761" />
                    <RANKING order="4" place="4" resultid="5775" />
                    <RANKING order="5" place="5" resultid="4319" />
                    <RANKING order="6" place="6" resultid="4696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2172" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4405" />
                    <RANKING order="2" place="2" resultid="4298" />
                    <RANKING order="3" place="3" resultid="6683" />
                    <RANKING order="4" place="-1" resultid="4386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2173" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3266" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="5650" />
                    <RANKING order="4" place="4" resultid="8186" />
                    <RANKING order="5" place="5" resultid="5731" />
                    <RANKING order="6" place="-1" resultid="3813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2174" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3260" />
                    <RANKING order="2" place="2" resultid="5992" />
                    <RANKING order="3" place="3" resultid="3236" />
                    <RANKING order="4" place="4" resultid="3768" />
                    <RANKING order="5" place="5" resultid="5944" />
                    <RANKING order="6" place="6" resultid="4282" />
                    <RANKING order="7" place="7" resultid="6743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2175" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7683" />
                    <RANKING order="2" place="2" resultid="2837" />
                    <RANKING order="3" place="3" resultid="7689" />
                    <RANKING order="4" place="4" resultid="5842" />
                    <RANKING order="5" place="5" resultid="3563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2176" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6670" />
                    <RANKING order="2" place="2" resultid="2810" />
                    <RANKING order="3" place="3" resultid="3776" />
                    <RANKING order="4" place="4" resultid="2796" />
                    <RANKING order="5" place="5" resultid="5720" />
                    <RANKING order="6" place="-1" resultid="6720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2177" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5636" />
                    <RANKING order="2" place="2" resultid="5984" />
                    <RANKING order="3" place="3" resultid="2781" />
                    <RANKING order="4" place="4" resultid="6005" />
                    <RANKING order="5" place="5" resultid="3856" />
                    <RANKING order="6" place="6" resultid="3242" />
                    <RANKING order="7" place="7" resultid="8176" />
                    <RANKING order="8" place="-1" resultid="2192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2178" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3572" />
                    <RANKING order="2" place="2" resultid="3759" />
                    <RANKING order="3" place="3" resultid="5043" />
                    <RANKING order="4" place="4" resultid="3552" />
                    <RANKING order="5" place="5" resultid="3588" />
                    <RANKING order="6" place="6" resultid="3193" />
                    <RANKING order="7" place="-1" resultid="5012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2179" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4607" />
                    <RANKING order="2" place="2" resultid="7724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2180" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2181" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2182" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2183" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="2184" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10286" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10287" daytime="11:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10288" daytime="11:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10289" daytime="11:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10290" daytime="12:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10291" daytime="12:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10292" daytime="12:15" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="SPCHR" name="UKS SP 8 Chrzanów" nation="POL" region="MAL" shortname="SP 8 Chrzanów">
          <CONTACT email="abalp@poczta.onet.pl" name="Zabrzański" phone="692076808" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2186">
              <RESULTS>
                <RESULT eventid="1162" status="DNS" swimtime="00:00:00.00" resultid="2187" heatid="10298" lane="8" entrytime="00:24:07.00" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="2188" heatid="10136" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1228" status="DSQ" swimtime="00:01:12.96" resultid="2189" heatid="10151" lane="5" entrytime="00:01:10.50" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="2190" heatid="10218" lane="2" entrytime="00:02:45.00" />
                <RESULT eventid="1574" points="597" swimtime="00:00:31.00" resultid="2191" heatid="10251" lane="5" entrytime="00:00:30.70" />
                <RESULT eventid="1686" status="DNS" swimtime="00:00:00.00" resultid="2192" heatid="10288" lane="4" entrytime="00:06:05.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEINO" name="KP Delfin Inowrocław" nation="POL" region="KUJ" shortname="Delfin Inowrocław">
          <CONTACT city="INOWROCŁAW" name="KP DELFIN INOWROCŁAW" phone="604667374" state="KUJ-P" street="WIERZBIŃSKIEGO" zip="88-100" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="ZYGMUNT" gender="M" lastname="LEWANDOWSKI" nation="POL" athleteid="2194">
              <RESULTS>
                <RESULT eventid="1077" points="325" swimtime="00:00:52.31" resultid="2195" heatid="10101" lane="1" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1162" points="645" swimtime="00:29:33.96" resultid="2196" heatid="10301" lane="5" entrytime="00:30:00.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="538" swimtime="00:03:28.51" resultid="2197" heatid="10216" lane="8" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="415" swimtime="00:02:03.41" resultid="2198" heatid="10235" lane="2" entrytime="00:02:00.00" entrycourse="LCM" />
                <RESULT eventid="1686" points="511" swimtime="00:07:33.50" resultid="2199" heatid="10286" lane="3" entrytime="00:07:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.15" />
                    <SPLIT distance="200" swimtime="00:03:48.21" />
                    <SPLIT distance="300" swimtime="00:05:44.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZALM" name="AZS Almamer" nation="POL">
          <CONTACT city="warszawa" email="udyta.judi@vp.pl" name="soltyk" phone="504 412 418j" street="bagatela" zip="00-585" />
          <ATHLETES>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="2202">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1141" points="642" swimtime="00:10:49.38" resultid="2203" heatid="10293" lane="3" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="200" swimtime="00:02:35.01" />
                    <SPLIT distance="300" swimtime="00:03:57.37" />
                    <SPLIT distance="400" swimtime="00:05:20.06" />
                    <SPLIT distance="500" swimtime="00:06:42.84" />
                    <SPLIT distance="600" swimtime="00:08:05.62" />
                    <SPLIT distance="700" swimtime="00:09:28.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1670" points="604" swimtime="00:05:16.79" resultid="2204" heatid="10285" lane="3" entrytime="00:05:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="200" swimtime="00:02:34.08" />
                    <SPLIT distance="300" swimtime="00:03:55.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMTS" name="Swimming Masters Team Szczecin" nation="POL" shortname="Masters Team Szczecin">
          <CONTACT email="milosz@smts.pl" name="Kaczanowski Miłosz" phone="888 18 1234" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-22" firstname="MIŁOSZ" gender="M" lastname="KACZANOWSKI" nation="POL" athleteid="2206">
              <RESULTS>
                <RESULT eventid="1077" points="879" swimtime="00:00:28.59" resultid="2207" heatid="10100" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1109" points="818" swimtime="00:02:29.48" resultid="2208" heatid="10122" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="592" swimtime="00:02:48.87" resultid="2209" heatid="10166" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="747" swimtime="00:05:34.67" resultid="2211" heatid="10231" lane="2" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.88" />
                    <SPLIT distance="200" swimtime="00:02:46.57" />
                    <SPLIT distance="300" swimtime="00:04:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="854" swimtime="00:01:04.65" resultid="2212" heatid="10236" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="1195" points="692" swimtime="00:00:32.62" resultid="2337" heatid="10132" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1401" points="755" reactiontime="+71" swimtime="00:01:11.46" resultid="2338" heatid="10198" lane="4" entrytime="00:02:00.00" />
                <RESULT eventid="1606" points="735" reactiontime="+69" swimtime="00:02:36.16" resultid="2339" heatid="10266" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02111" name="KS Górnik Sosnowiec" nation="POL" region="SLA" shortname="Górnik Sosnowiec">
          <CONTACT city="Sosnowiec" email="gosos@wp.pl" internet="http://plywanie.sosnowiec.pl/" name="KS Górnik Sosnowiec" phone="531309751" state="SLA" street="ul. Hubala-Dobrzańskiego 99" zip="41-200" />
        </CLUB>
        <CLUB type="CLUB" code="SATCZ" name="Sambor Tczew" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1986-11-14" firstname="Kamila" gender="F" lastname="Ormianin" nation="POL" athleteid="2242">
              <RESULTS>
                <RESULT eventid="1141" points="497" swimtime="00:11:41.01" resultid="2243" heatid="10293" lane="6" entrytime="00:10:56.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="200" swimtime="00:02:44.82" />
                    <SPLIT distance="300" swimtime="00:04:12.48" />
                    <SPLIT distance="400" swimtime="00:05:41.55" />
                    <SPLIT distance="500" swimtime="00:07:12.29" />
                    <SPLIT distance="600" swimtime="00:08:43.74" />
                    <SPLIT distance="700" swimtime="00:10:12.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="597" swimtime="00:02:25.92" resultid="2244" heatid="10213" lane="4" entrytime="00:02:22.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1670" points="588" swimtime="00:05:17.50" resultid="2245" heatid="10285" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="200" swimtime="00:02:36.97" />
                    <SPLIT distance="300" swimtime="00:03:58.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="2322">
              <RESULTS>
                <RESULT eventid="1369" points="732" swimtime="00:00:31.38" resultid="2324" heatid="10192" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1574" points="612" swimtime="00:00:26.77" resultid="2325" heatid="10257" lane="1" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra " gender="F" lastname="Hebel" nation="POL" athleteid="2571">
              <RESULTS>
                <RESULT eventid="1178" points="348" swimtime="00:00:43.25" resultid="2572" heatid="10128" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1212" points="410" swimtime="00:01:17.29" resultid="2573" heatid="10144" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1385" status="DNS" swimtime="00:00:00.00" resultid="2574" heatid="10195" lane="2" entrytime="00:01:37.00" />
                <RESULT eventid="1449" points="347" swimtime="00:02:54.82" resultid="2575" heatid="10212" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DSQ" swimtime="00:00:34.14" resultid="2576" heatid="10244" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="2577">
              <RESULTS>
                <RESULT eventid="1228" points="485" swimtime="00:01:04.35" resultid="2578" heatid="10154" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="1324" points="491" swimtime="00:02:59.86" resultid="2579" heatid="10176" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="551" swimtime="00:00:34.50" resultid="2580" heatid="10192" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1574" points="499" swimtime="00:00:28.67" resultid="2581" heatid="10253" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1654" points="461" swimtime="00:01:21.77" resultid="2582" heatid="10280" lane="2" entrytime="00:01:19.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1125" swimtime="00:01:59.02" resultid="2583" heatid="10125" lane="7" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2242" number="1" />
                    <RELAYPOSITION athleteid="2577" number="2" />
                    <RELAYPOSITION athleteid="2571" number="3" />
                    <RELAYPOSITION athleteid="2322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+103" swimtime="00:02:18.36" resultid="2584" heatid="10269" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2242" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="2577" number="2" />
                    <RELAYPOSITION athleteid="2571" number="3" />
                    <RELAYPOSITION athleteid="2322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NIEZRZ" name="Niezrzeszony" nation="POL">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK PIOTR" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1977-02-01" firstname="Mariusz" gender="M" lastname="Wójcicki" nation="POL" athleteid="2246">
              <RESULTS>
                <RESULT eventid="1077" points="494" swimtime="00:00:31.80" resultid="2248" heatid="10107" lane="3" entrytime="00:00:31.15" />
                <RESULT eventid="1195" points="541" swimtime="00:00:33.72" resultid="2249" heatid="10139" lane="6" entrytime="00:00:33.25" />
                <RESULT eventid="1401" points="408" reactiontime="+75" swimtime="00:01:19.29" resultid="2250" heatid="10203" lane="3" entrytime="00:01:15.51" />
                <RESULT eventid="1542" points="464" swimtime="00:01:13.71" resultid="2251" heatid="10239" lane="2" entrytime="00:01:10.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-08-25" firstname="Krzysztof" gender="M" lastname="Micorek" nation="POL" athleteid="2335">
              <RESULTS>
                <RESULT eventid="1077" points="743" swimtime="00:00:27.39" resultid="2336" heatid="10110" lane="6" entrytime="00:00:27.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" athleteid="2346">
              <RESULTS>
                <RESULT eventid="1542" points="674" swimtime="00:01:03.34" resultid="8142" heatid="10239" lane="4" entrytime="00:01:04.55" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1162" points="675" swimtime="00:18:21.99" resultid="2348" heatid="10296" lane="4" entrytime="00:18:29.55" />
                <RESULT eventid="1292" points="770" swimtime="00:02:17.29" resultid="2349" heatid="10166" lane="4" entrytime="00:02:16.35">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="518" swimtime="00:02:17.79" resultid="2350" heatid="10223" lane="3" entrytime="00:02:08.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="516" swimtime="00:05:38.82" resultid="2351" heatid="10231" lane="5" entrytime="00:05:09.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="200" swimtime="00:02:47.26" />
                    <SPLIT distance="300" swimtime="00:04:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="672" swimtime="00:04:35.65" resultid="2352" heatid="10292" lane="3" entrytime="00:04:37.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="200" swimtime="00:02:18.31" />
                    <SPLIT distance="300" swimtime="00:03:28.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Sebastian" gender="M" lastname="Pikusa" nation="POL" athleteid="2353">
              <RESULTS>
                <RESULT eventid="1077" points="719" swimtime="00:00:28.30" resultid="2354" heatid="10110" lane="8" entrytime="00:00:28.15" />
                <RESULT eventid="1162" points="493" swimtime="00:20:23.47" resultid="2355" heatid="10296" lane="5" entrytime="00:18:35.98" />
                <RESULT eventid="1292" points="474" swimtime="00:02:41.43" resultid="2356" heatid="10166" lane="5" entrytime="00:02:19.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="553" swimtime="00:00:31.85" resultid="2357" heatid="10139" lane="4" entrytime="00:00:31.99" />
                <RESULT eventid="1401" points="409" reactiontime="+83" swimtime="00:01:15.70" resultid="2358" heatid="10205" lane="7" entrytime="00:01:07.88" />
                <RESULT eventid="1497" points="407" swimtime="00:06:06.82" resultid="2359" heatid="10231" lane="6" entrytime="00:05:15.91">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="200" swimtime="00:02:58.55" />
                    <SPLIT distance="300" swimtime="00:04:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="677" swimtime="00:01:03.24" resultid="2360" heatid="10240" lane="7" entrytime="00:01:02.55" />
                <RESULT eventid="1606" points="372" reactiontime="+80" swimtime="00:02:53.72" resultid="2361" heatid="10266" lane="4" entrytime="00:02:24.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="2373">
              <RESULTS>
                <RESULT eventid="1385" points="677" reactiontime="+96" swimtime="00:01:33.36" resultid="2374" heatid="10194" lane="3" entrytime="00:01:44.13" />
                <RESULT eventid="1590" points="808" reactiontime="+108" swimtime="00:03:19.14" resultid="2375" heatid="10259" lane="8" entrytime="00:03:36.48">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-07-31" firstname="Tomasz" gender="M" lastname="Jaron " nation="POL" athleteid="2482">
              <RESULTS>
                <RESULT eventid="1162" points="373" swimtime="00:23:37.68" resultid="2483" heatid="10298" lane="6" entrytime="00:23:30.00" />
                <RESULT eventid="1324" points="431" swimtime="00:03:18.90" resultid="2484" heatid="10175" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="2485" heatid="10229" lane="8" entrytime="00:06:45.00" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="2486" heatid="10278" lane="8" entrytime="00:01:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-16" firstname="PIOTR" gender="M" lastname="URBAŃCZYK" nation="POL" athleteid="2554">
              <RESULTS>
                <RESULT eventid="1195" points="695" swimtime="00:00:29.52" resultid="2555" heatid="10140" lane="4" entrytime="00:00:29.99" />
                <RESULT eventid="1401" points="694" reactiontime="+76" swimtime="00:01:03.49" resultid="2556" heatid="10205" lane="4" entrytime="00:01:03.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-12-09" firstname="Natalia" gender="F" lastname="Borek" nation="POL" athleteid="2729">
              <RESULTS>
                <RESULT eventid="1178" points="803" swimtime="00:00:32.04" resultid="2730" heatid="10130" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1212" points="657" swimtime="00:01:04.20" resultid="2731" heatid="10146" lane="5" entrytime="00:01:04.00" />
                <RESULT eventid="1385" points="765" reactiontime="+74" swimtime="00:01:10.05" resultid="2732" heatid="10197" lane="4" entrytime="00:01:07.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="Zielezinski" nation="POL" athleteid="2744">
              <RESULTS>
                <RESULT eventid="1162" points="364" swimtime="00:28:29.67" resultid="2745" heatid="10299" lane="1" entrytime="00:26:00.00" />
                <RESULT eventid="1686" points="380" swimtime="00:06:47.09" resultid="3552" heatid="10287" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="200" swimtime="00:03:07.47" />
                    <SPLIT distance="300" swimtime="00:04:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="537" swimtime="00:00:41.12" resultid="3832" heatid="10136" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-02" firstname="DOROTA" gender="F" lastname="MORTKA" nation="POL" athleteid="2746">
              <RESULTS>
                <RESULT eventid="1449" points="448" swimtime="00:02:40.60" resultid="2747" heatid="10213" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="F" lastname="Kotusińska" nation="POL" athleteid="4470">
              <RESULTS>
                <RESULT eventid="1212" points="383" swimtime="00:01:19.11" resultid="4471" heatid="10144" lane="1" entrytime="00:01:18.00" />
                <RESULT eventid="1558" points="427" swimtime="00:00:35.05" resultid="4472" heatid="10244" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-12" firstname="Marcin" gender="M" lastname="Garbacki" nation="POL" athleteid="4473">
              <RESULTS>
                <RESULT eventid="1228" points="448" swimtime="00:01:06.07" resultid="4474" heatid="10153" lane="2" entrytime="00:01:06.00" />
                <RESULT eventid="1574" points="488" swimtime="00:00:28.88" resultid="4475" heatid="10254" lane="6" entrytime="00:00:28.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="Jąkalski" nation="POL" athleteid="4483">
              <RESULTS>
                <RESULT eventid="1195" points="629" swimtime="00:00:30.51" resultid="4484" heatid="10140" lane="3" entrytime="00:00:30.01" />
                <RESULT eventid="1401" points="555" reactiontime="+68" swimtime="00:01:08.38" resultid="4485" heatid="10205" lane="2" entrytime="00:01:07.50" />
                <RESULT eventid="1606" points="485" reactiontime="+81" swimtime="00:02:38.94" resultid="4486" heatid="10266" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="Dziekoński  " nation="POL" athleteid="5020">
              <RESULTS>
                <RESULT eventid="1077" points="423" swimtime="00:00:45.42" resultid="5021" heatid="10101" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="1162" points="378" swimtime="00:30:43.24" resultid="5022" heatid="10300" lane="8" entrytime="00:29:35.00" />
                <RESULT eventid="1195" points="411" swimtime="00:00:51.37" resultid="5023" heatid="10134" lane="3" entrytime="00:00:47.00" />
                <RESULT eventid="1228" points="336" swimtime="00:01:36.44" resultid="5024" heatid="10148" lane="1" entrytime="00:01:35.00" />
                <RESULT eventid="1401" points="338" reactiontime="+82" swimtime="00:02:01.30" resultid="5025" heatid="10199" lane="2" entrytime="00:01:54.00" />
                <RESULT eventid="1465" points="347" swimtime="00:03:40.02" resultid="5026" heatid="10215" lane="5" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="391" swimtime="00:00:41.20" resultid="5027" heatid="10247" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1606" points="342" reactiontime="+98" swimtime="00:04:24.87" resultid="5028" heatid="10262" lane="6" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:11.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="5035">
              <RESULTS>
                <RESULT eventid="1077" points="535" swimtime="00:00:37.39" resultid="5036" heatid="10103" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1162" points="430" swimtime="00:26:57.68" resultid="5037" heatid="10300" lane="3" entrytime="00:28:30.00" />
                <RESULT eventid="1195" points="625" swimtime="00:00:39.10" resultid="5038" heatid="10137" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1228" points="570" swimtime="00:01:15.20" resultid="5039" heatid="10150" lane="2" entrytime="00:01:14.00" />
                <RESULT eventid="1401" points="529" reactiontime="+89" swimtime="00:01:30.97" resultid="5040" heatid="10201" lane="3" entrytime="00:01:29.00" />
                <RESULT eventid="1465" points="508" swimtime="00:02:56.94" resultid="5041" heatid="10218" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="581" swimtime="00:00:32.69" resultid="5042" heatid="10251" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1686" points="419" swimtime="00:06:34.13" resultid="5043" heatid="10288" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.18" />
                    <SPLIT distance="200" swimtime="00:03:09.73" />
                    <SPLIT distance="300" swimtime="00:04:54.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Witold" gender="M" lastname="SZCZECHLA" nation="POL" athleteid="5667">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="5668" heatid="10104" lane="7" entrytime="00:00:37.50" />
                <RESULT eventid="1109" points="352" swimtime="00:03:30.34" resultid="5669" heatid="10117" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="226" swimtime="00:01:43.57" resultid="5670" heatid="10236" lane="3" entrytime="00:01:33.00" />
                <RESULT eventid="1654" points="381" swimtime="00:01:40.32" resultid="5671" heatid="10277" lane="6" entrytime="00:01:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-10" firstname="Emil" gender="M" lastname="Paciorkowski" nation="POL" athleteid="8170">
              <RESULTS>
                <RESULT eventid="1077" points="229" swimtime="00:00:45.84" resultid="8171" heatid="10101" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1228" points="348" swimtime="00:01:23.42" resultid="8172" heatid="10149" lane="1" entrytime="00:01:24.00" />
                <RESULT eventid="1292" status="DNF" swimtime="00:00:00.00" resultid="8173" heatid="10163" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="164" reactiontime="+107" swimtime="00:02:03.44" resultid="8174" heatid="10199" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="1574" points="437" swimtime="00:00:34.39" resultid="8175" heatid="10249" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1686" points="244" swimtime="00:07:37.70" resultid="8176" heatid="10288" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.95" />
                    <SPLIT distance="200" swimtime="00:03:42.08" />
                    <SPLIT distance="300" swimtime="00:05:42.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03001" name="MUKP Just Swim Jelenia Góra" nation="POL" region="WR" shortname="Just Swim">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz Marcin" phone="509071929" zip="58-506" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="WASZKEWICZ" nation="POL" license="M0300120009" athleteid="2257">
              <RESULTS>
                <RESULT eventid="1077" points="831" swimtime="00:00:26.86" resultid="2258" heatid="10110" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1228" points="667" swimtime="00:00:57.95" resultid="2259" heatid="10158" lane="4" entrytime="00:00:54.00" />
                <RESULT eventid="1574" points="756" swimtime="00:00:25.32" resultid="2260" heatid="10257" lane="4" entrytime="00:00:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" name="MOSiR Ostrowiec" nation="POL">
          <CONTACT name="Różalski" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="M01012200001" athleteid="2262">
              <RESULTS>
                <RESULT eventid="1077" points="803" swimtime="00:00:34.26" resultid="2263" heatid="10105" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1109" points="640" swimtime="00:03:20.63" resultid="2264" heatid="10116" lane="5" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="680" swimtime="00:01:15.09" resultid="2265" heatid="10150" lane="3" entrytime="00:01:14.00" />
                <RESULT eventid="1292" points="410" swimtime="00:04:06.96" resultid="2266" heatid="10164" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="541" swimtime="00:00:44.41" resultid="2267" heatid="10187" lane="2" entrytime="00:00:42.50" />
                <RESULT eventid="1497" points="463" swimtime="00:08:03.44" resultid="2268" heatid="10228" lane="8" entrytime="00:07:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.46" />
                    <SPLIT distance="200" swimtime="00:04:06.72" />
                    <SPLIT distance="300" swimtime="00:06:18.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="417" swimtime="00:01:41.80" resultid="2269" heatid="10236" lane="2" entrytime="00:01:40.00" />
                <RESULT eventid="1574" points="581" swimtime="00:00:33.87" resultid="2270" heatid="10250" lane="2" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSKRA" name="AZS UJ CM Kraków " nation="POL" shortname="AZS UJ  Kraków ">
          <ATHLETES>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="2312">
              <RESULTS>
                <RESULT eventid="1061" points="603" swimtime="00:00:32.66" resultid="2314" heatid="10099" lane="5" entrytime="00:00:32.23" />
                <RESULT eventid="1093" points="709" swimtime="00:02:35.74" resultid="2315" heatid="10113" lane="4" entrytime="00:02:32.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="703" swimtime="00:01:02.75" resultid="2316" heatid="10146" lane="4" entrytime="00:01:02.60" />
                <RESULT eventid="1308" points="606" swimtime="00:02:59.53" resultid="2317" heatid="10169" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="701" swimtime="00:00:36.92" resultid="2318" heatid="10182" lane="5" entrytime="00:00:36.21" />
                <RESULT eventid="1481" points="626" swimtime="00:05:39.59" resultid="2319" heatid="10225" lane="4" entrytime="00:05:19.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                    <SPLIT distance="200" swimtime="00:02:44.46" />
                    <SPLIT distance="300" swimtime="00:04:19.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="669" swimtime="00:00:29.28" resultid="2320" heatid="10245" lane="4" entrytime="00:00:28.99" />
                <RESULT eventid="1638" points="628" swimtime="00:01:22.38" resultid="2321" heatid="10273" lane="5" entrytime="00:01:20.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RACIB" name="AZS PWSZ Racibórz" nation="POL" region="ŚLĄSK" shortname="AZS Racibórz">
          <CONTACT city="Racibórz" email="m,kunicki@" name="Marcin Kunicki" phone="504 233 267" state="ŚLĄSK" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="2327">
              <RESULTS>
                <RESULT eventid="1109" points="635" swimtime="00:02:59.99" resultid="2328" heatid="10118" lane="5" entrytime="00:03:02.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="502" swimtime="00:03:11.47" resultid="2329" heatid="10165" lane="2" entrytime="00:03:06.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="563" swimtime="00:03:19.51" resultid="2330" heatid="10175" lane="7" entrytime="00:03:14.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="649" swimtime="00:00:38.34" resultid="2331" heatid="10189" lane="7" entrytime="00:00:38.24" entrycourse="SCM" />
                <RESULT eventid="1497" points="617" swimtime="00:06:36.97" resultid="2332" heatid="10230" lane="1" entrytime="00:06:17.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="200" swimtime="00:03:12.81" />
                    <SPLIT distance="300" swimtime="00:05:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="404" swimtime="00:01:27.01" resultid="2333" heatid="10238" lane="8" entrytime="00:01:19.65" entrycourse="SCM" />
                <RESULT eventid="1654" points="588" swimtime="00:01:28.67" resultid="2334" heatid="10279" lane="5" entrytime="00:01:24.53" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SZCZC" name="MKP Szczecin" nation="POL" region="ZAC">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" name="Kowalczyk" phone="509758055" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="2363">
              <RESULTS>
                <RESULT eventid="1141" points="869" swimtime="00:10:45.92" resultid="2364" heatid="10293" lane="4" entrytime="00:10:29.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="200" swimtime="00:02:34.13" />
                    <SPLIT distance="300" swimtime="00:03:55.87" />
                    <SPLIT distance="400" swimtime="00:05:17.42" />
                    <SPLIT distance="500" swimtime="00:06:39.39" />
                    <SPLIT distance="600" swimtime="00:08:01.85" />
                    <SPLIT distance="700" swimtime="00:09:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="760" swimtime="00:01:09.61" resultid="2365" heatid="10146" lane="8" entrytime="00:01:08.25" />
                <RESULT eventid="1449" points="804" swimtime="00:02:28.35" resultid="2366" heatid="10213" lane="5" entrytime="00:02:23.65">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="793" swimtime="00:05:16.50" resultid="2367" heatid="10285" lane="5" entrytime="00:05:07.29">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="200" swimtime="00:02:33.76" />
                    <SPLIT distance="300" swimtime="00:03:55.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="2368">
              <RESULTS>
                <RESULT eventid="1162" points="544" swimtime="00:20:05.34" resultid="2369" heatid="10296" lane="1" entrytime="00:20:15.00" />
                <RESULT eventid="1228" points="554" swimtime="00:01:02.62" resultid="2370" heatid="10156" lane="3" entrytime="00:01:01.50" />
                <RESULT eventid="1465" points="608" swimtime="00:02:17.11" resultid="2371" heatid="10222" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="565" swimtime="00:04:56.73" resultid="2372" heatid="10291" lane="5" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="200" swimtime="00:02:27.12" />
                    <SPLIT distance="300" swimtime="00:03:43.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ŹILINA" name="PSK Žilina" nation="SVK">
          <ATHLETES>
            <ATHLETE birthdate="1960-11-14" firstname="Rastislav" gender="M" lastname="Pavlik" nation="SVK" athleteid="2376">
              <RESULTS>
                <RESULT eventid="1077" points="797" swimtime="00:00:29.90" resultid="2378" heatid="10108" lane="6" entrytime="00:00:30.40" />
                <RESULT eventid="1109" points="827" swimtime="00:02:38.25" resultid="2379" heatid="10121" lane="6" entrytime="00:02:34.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="824" swimtime="00:00:32.66" resultid="2380" heatid="10140" lane="8" entrytime="00:00:31.90" />
                <RESULT eventid="1228" points="732" swimtime="00:01:03.12" resultid="2381" heatid="10156" lane="1" entrytime="00:01:01.70" />
                <RESULT eventid="1369" points="787" swimtime="00:00:34.87" resultid="2382" heatid="10191" lane="5" entrytime="00:00:34.10" />
                <RESULT eventid="1401" points="815" reactiontime="+75" swimtime="00:01:11.92" resultid="2383" heatid="10204" lane="4" entrytime="00:01:09.30" />
                <RESULT eventid="1574" points="682" swimtime="00:00:28.82" resultid="2384" heatid="10256" lane="1" entrytime="00:00:27.40" />
                <RESULT eventid="1654" points="753" swimtime="00:01:19.98" resultid="2385" heatid="10280" lane="4" entrytime="00:01:17.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGRY" name="Marlin Gryfino" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski " nation="POL" athleteid="2476">
              <RESULTS>
                <RESULT eventid="1109" points="548" swimtime="00:03:16.86" resultid="2478" heatid="10117" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="576" swimtime="00:03:32.15" resultid="2479" heatid="10173" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="539" swimtime="00:00:42.09" resultid="2480" heatid="10187" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1654" points="548" swimtime="00:01:36.49" resultid="2481" heatid="10277" lane="3" entrytime="00:01:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSWAR" name="AZS SGGW Warszawa" nation="POL" shortname="AZS Warszawa">
          <CONTACT name="Nawrocka Manuela" phone="+48606704926" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="2488">
              <RESULTS>
                <RESULT eventid="1093" points="520" swimtime="00:02:52.72" resultid="2489" heatid="10113" lane="8" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="468" swimtime="00:00:38.37" resultid="2490" heatid="10130" lane="1" entrytime="00:00:36.10" />
                <RESULT eventid="1308" points="452" swimtime="00:03:17.87" resultid="2491" heatid="10169" lane="1" entrytime="00:03:15.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="457" swimtime="00:00:42.57" resultid="2492" heatid="10182" lane="1" entrytime="00:00:41.60" />
                <RESULT eventid="1385" points="452" reactiontime="+78" swimtime="00:01:23.46" resultid="2493" heatid="10197" lane="2" entrytime="00:01:17.50" />
                <RESULT eventid="1558" points="589" swimtime="00:00:30.54" resultid="2494" heatid="10245" lane="7" entrytime="00:00:30.99" />
                <RESULT eventid="1590" points="424" reactiontime="+80" swimtime="00:03:00.47" resultid="2495" heatid="10260" lane="2" entrytime="00:02:50.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOSIE" name="Wodnik Siemianowice Śląskie" nation="POL" shortname="Wodnik Siemianowice">
          <CONTACT name="Szymik" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="2497">
              <RESULTS>
                <RESULT eventid="1077" points="490" swimtime="00:00:35.17" resultid="2498" heatid="10105" lane="7" entrytime="00:00:35.80" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1162" points="578" swimtime="00:21:54.93" resultid="2499" heatid="10297" lane="1" entrytime="00:22:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIWAR" name="Sinnet Warszawa" nation="POL">
          <CONTACT city="Warszawa" email="piotrbarski@uw.edu.pl" name="Barski" street="Polinezyjska" zip="02-777" />
          <ATHLETES>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="2501">
              <RESULTS>
                <RESULT eventid="1077" points="834" swimtime="00:00:29.09" resultid="2502" heatid="10109" lane="5" entrytime="00:00:29.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1228" points="813" swimtime="00:00:58.66" resultid="2503" heatid="10153" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1324" points="761" swimtime="00:02:48.66" resultid="2504" heatid="10177" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="702" swimtime="00:00:34.55" resultid="2505" heatid="10192" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1465" points="750" swimtime="00:02:14.85" resultid="2506" heatid="10223" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="710" swimtime="00:00:27.49" resultid="2507" heatid="10257" lane="2" entrytime="00:00:26.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1654" points="754" swimtime="00:01:15.51" resultid="2508" heatid="10281" lane="3" entrytime="00:01:14.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-25" firstname="Agnieszka" gender="F" lastname="Besler" nation="POL" athleteid="2509">
              <RESULTS>
                <RESULT eventid="1061" points="456" swimtime="00:00:37.98" resultid="2510" heatid="10098" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="1308" points="452" swimtime="00:03:28.95" resultid="2511" heatid="10168" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="475" swimtime="00:00:42.88" resultid="2512" heatid="10181" lane="3" entrytime="00:00:42.50" />
                <RESULT eventid="1558" points="562" swimtime="00:00:32.47" resultid="2513" heatid="10243" lane="7" entrytime="00:00:36.50" />
                <RESULT eventid="1638" points="468" swimtime="00:01:35.54" resultid="2514" heatid="10272" lane="6" entrytime="00:01:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-18" firstname="Joanna" gender="F" lastname="Janicka" nation="POL" athleteid="2515">
              <RESULTS>
                <RESULT eventid="1061" points="655" swimtime="00:00:33.55" resultid="2516" heatid="10099" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1178" points="637" swimtime="00:00:35.38" resultid="2517" heatid="10126" lane="1" />
                <RESULT eventid="1212" points="683" swimtime="00:01:05.22" resultid="2518" heatid="10146" lane="6" entrytime="00:01:07.00" />
                <RESULT eventid="1449" points="569" swimtime="00:02:28.28" resultid="2519" heatid="10212" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DSQ" swimtime="00:00:29.32" resultid="2520" heatid="10245" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIGLI" name="Sikret Gliwice" nation="POL">
          <CONTACT city="GLIWICE" email="JOANNAECO@WP.PL" name="ZAGAŁA JOANNA" phone="601427257" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="2522">
              <RESULTS>
                <RESULT eventid="1093" points="335" swimtime="00:03:54.87" resultid="9024" heatid="10111" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="361" swimtime="00:04:10.58" resultid="9025" heatid="10167" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="428" swimtime="00:00:50.30" resultid="9026" heatid="10179" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1449" points="314" swimtime="00:03:30.70" resultid="9027" heatid="10210" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="383" swimtime="00:00:40.10" resultid="9028" heatid="10242" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1590" points="369" reactiontime="+87" swimtime="00:03:58.43" resultid="9029" heatid="10258" lane="5" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="2529">
              <RESULTS>
                <RESULT eventid="1061" points="280" swimtime="00:00:51.28" resultid="9030" heatid="10097" lane="1" entrytime="00:00:47.00" />
                <RESULT eventid="1276" points="285" swimtime="00:04:42.32" resultid="9031" heatid="10162" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="420" swimtime="00:00:51.33" resultid="9032" heatid="10180" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1449" points="306" swimtime="00:03:43.08" resultid="9033" heatid="10210" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" status="DSQ" swimtime="00:02:19.12" resultid="9034" heatid="10232" lane="2" entrytime="00:02:00.00" />
                <RESULT eventid="1638" points="386" swimtime="00:01:59.81" resultid="9035" heatid="10271" lane="4" entrytime="00:01:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-28" firstname="Łukasz" gender="M" lastname="Stolarczyk" nation="POL" athleteid="2536">
              <RESULTS>
                <RESULT eventid="1077" points="690" swimtime="00:00:28.58" resultid="9036" heatid="10110" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1228" points="703" swimtime="00:00:56.96" resultid="9037" heatid="10158" lane="8" entrytime="00:00:59.00" />
                <RESULT eventid="1542" points="699" swimtime="00:01:02.78" resultid="9038" heatid="10240" lane="2" entrytime="00:01:02.00" />
                <RESULT eventid="1574" points="675" swimtime="00:00:26.29" resultid="9039" heatid="10257" lane="6" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-15" firstname="Mieczysław" gender="M" lastname="Mydłowski" nation="POL" athleteid="2540">
              <RESULTS>
                <RESULT eventid="1228" points="546" swimtime="00:01:09.57" resultid="9040" heatid="10152" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="1324" points="524" swimtime="00:03:19.96" resultid="9041" heatid="10174" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="475" reactiontime="+93" swimtime="00:01:26.11" resultid="9042" heatid="10202" lane="7" entrytime="00:01:25.00" />
                <RESULT eventid="1465" points="401" swimtime="00:02:48.44" resultid="9043" heatid="10221" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="551" swimtime="00:00:30.93" resultid="9044" heatid="10250" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1654" points="520" swimtime="00:01:30.48" resultid="9045" heatid="10278" lane="2" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-06" firstname="Arkadiusz" gender="M" lastname="Bednarek" nation="POL" athleteid="2547">
              <RESULTS>
                <RESULT eventid="1077" points="220" swimtime="00:00:44.11" resultid="9046" heatid="10102" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1228" points="233" swimtime="00:01:26.79" resultid="9047" heatid="10149" lane="6" entrytime="00:01:22.00" />
                <RESULT eventid="1369" points="282" swimtime="00:00:44.97" resultid="9048" heatid="10185" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1574" points="267" swimtime="00:00:37.92" resultid="9049" heatid="10247" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+80" swimtime="00:02:40.08" resultid="9050" heatid="10268" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2540" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2529" number="2" />
                    <RELAYPOSITION athleteid="2536" number="3" />
                    <RELAYPOSITION athleteid="2522" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" status="DSQ" swimtime="00:02:20.99" resultid="9051" heatid="10124" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2522" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2540" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2529" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2536" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AJCZE" name="KU AZS AJD Częstochowa" nation="POL" shortname="AJD Częstochowa">
          <CONTACT city="Częstochowa" name="Klub Uczelniany AZS AJD Częstochowa" street="Armii Krajowej" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-28" firstname="Piotr" gender="M" lastname="Trzcionka" nation="POL" athleteid="2558">
              <RESULTS>
                <RESULT eventid="1109" points="531" swimtime="00:02:32.43" resultid="2559" heatid="10121" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="540" swimtime="00:01:00.63" resultid="2560" heatid="10157" lane="3" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1401" points="470" swimtime="00:01:09.91" resultid="2561" heatid="10205" lane="1" entrytime="00:01:08.00" entrycourse="LCM" />
                <RESULT eventid="1606" points="481" reactiontime="+72" swimtime="00:02:35.32" resultid="2562" heatid="10266" lane="3" entrytime="00:02:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKUT" name="WOPR Kutno" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1932-03-11" firstname="Kazimierz" gender="M" lastname="From" nation="POL" athleteid="2563">
              <RESULTS>
                <RESULT eventid="1195" points="160" swimtime="00:01:15.35" resultid="2565" heatid="10131" lane="4" />
                <RESULT eventid="1228" points="176" swimtime="00:02:17.85" resultid="2566" heatid="10147" lane="7" />
                <RESULT eventid="1401" points="160" reactiontime="+96" swimtime="00:02:51.08" resultid="2567" heatid="10198" lane="1" />
                <RESULT eventid="1465" points="213" swimtime="00:05:22.27" resultid="2568" heatid="10214" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="182" swimtime="00:00:58.44" resultid="2569" heatid="10246" lane="6" />
                <RESULT eventid="1606" points="157" reactiontime="+96" swimtime="00:06:20.34" resultid="2570" heatid="10261" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:03:01.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MACHE" name="Masters Chełm" nation="POL" region="LBL">
          <CONTACT city="Chełm" email="elzbietadz@gmail.com" name="Dziwisz Elżbieta" phone="660429651" state="LUB" street="Lubelska 139 D/13" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-01" firstname="Ireneusz" gender="M" lastname="Sokołowski" nation="POL" athleteid="2586">
              <RESULTS>
                <RESULT eventid="1195" points="170" swimtime="00:00:57.52" resultid="2587" heatid="10131" lane="3" />
                <RESULT eventid="1369" points="306" swimtime="00:00:49.27" resultid="2588" heatid="10183" lane="5" />
                <RESULT eventid="1654" points="240" swimtime="00:01:59.40" resultid="2589" heatid="10274" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Leszek" gender="M" lastname="Masłowski" nation="POL" athleteid="2590">
              <RESULTS>
                <RESULT eventid="1077" points="97" swimtime="00:01:09.13" resultid="2591" heatid="10100" lane="3" />
                <RESULT eventid="1109" points="148" swimtime="00:05:26.86" resultid="2592" heatid="10114" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="150" swimtime="00:02:04.27" resultid="2593" heatid="10147" lane="8" />
                <RESULT eventid="1324" points="188" swimtime="00:05:21.57" resultid="2594" heatid="10170" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="175" reactiontime="+91" swimtime="00:02:22.80" resultid="2595" heatid="10198" lane="7" />
                <RESULT eventid="1465" points="149" swimtime="00:04:40.04" resultid="2596" heatid="10214" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="90" swimtime="00:02:49.31" resultid="2597" heatid="10234" lane="3" />
                <RESULT eventid="1606" points="135" reactiontime="+103" swimtime="00:05:40.23" resultid="2598" heatid="10261" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:41.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Piotr" gender="M" lastname="Gryciuk" nation="POL" athleteid="2599">
              <RESULTS>
                <RESULT eventid="1077" points="749" swimtime="00:00:29.35" resultid="2600" heatid="10108" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1228" points="658" swimtime="00:01:01.41" resultid="2601" heatid="10155" lane="2" entrytime="00:01:03.00" />
                <RESULT eventid="1401" points="488" swimtime="00:01:17.12" resultid="2602" heatid="10203" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1542" points="520" swimtime="00:01:12.95" resultid="2603" heatid="10238" lane="7" entrytime="00:01:17.00" />
                <RESULT eventid="1574" points="633" swimtime="00:00:28.44" resultid="2604" heatid="10255" lane="1" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Elżbieta" gender="F" lastname="Dziwisz" nation="POL" athleteid="2605">
              <RESULTS>
                <RESULT eventid="1178" points="151" swimtime="00:01:09.47" resultid="2606" heatid="10126" lane="8" />
                <RESULT eventid="1308" points="215" swimtime="00:05:16.54" resultid="2607" heatid="10167" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" status="DSQ" swimtime="00:01:04.43" resultid="2608" heatid="10178" lane="4" />
                <RESULT eventid="1385" points="236" reactiontime="+70" swimtime="00:02:12.62" resultid="2609" heatid="10193" lane="1" />
                <RESULT eventid="1558" points="186" swimtime="00:00:54.29" resultid="2610" heatid="10241" lane="8" />
                <RESULT eventid="1638" points="226" swimtime="00:02:23.13" resultid="2611" heatid="10270" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Alicja" gender="F" lastname="Wątrobińska" nation="POL" athleteid="2612">
              <RESULTS>
                <RESULT eventid="1178" points="144" swimtime="00:01:13.22" resultid="2613" heatid="10126" lane="7" />
                <RESULT eventid="1352" points="168" swimtime="00:01:09.92" resultid="2614" heatid="10178" lane="5" />
                <RESULT eventid="1385" points="115" reactiontime="+91" swimtime="00:02:53.67" resultid="2615" heatid="10193" lane="7" />
                <RESULT eventid="1558" points="136" swimtime="00:01:02.43" resultid="2616" heatid="10241" lane="1" />
                <RESULT eventid="1638" points="147" swimtime="00:02:43.61" resultid="2617" heatid="10270" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="2622">
              <RESULTS>
                <RESULT eventid="1195" points="256" swimtime="00:01:00.16" resultid="2623" heatid="10132" lane="7" />
                <RESULT eventid="1228" points="252" swimtime="00:01:46.09" resultid="2624" heatid="10147" lane="3" entrytime="00:01:49.00" />
                <RESULT eventid="1324" points="486" swimtime="00:04:07.89" resultid="2625" heatid="10171" lane="7" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="593" swimtime="00:00:45.48" resultid="2626" heatid="10186" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1465" points="168" swimtime="00:04:40.33" resultid="2627" heatid="10214" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="546" swimtime="00:01:47.08" resultid="2628" heatid="10275" lane="5" entrytime="00:01:47.00" />
                <RESULT eventid="1606" points="266" reactiontime="+111" swimtime="00:04:47.89" resultid="10310" heatid="10261" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:16.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00305" name="UKS NAWA Skierniewice" nation="POL" region="LOD" shortname="NAWA Skierniewice">
          <CONTACT name="Marcin Sarna" phone="603331973" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-11" firstname="Sebastian" gender="M" lastname="Krawczyk" nation="POL" license="S00305200017" athleteid="2630">
              <RESULTS>
                <RESULT eventid="1109" points="600" swimtime="00:02:26.37" resultid="2631" heatid="10122" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="591" swimtime="00:02:40.66" resultid="2632" heatid="10177" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="742" swimtime="00:00:31.28" resultid="2633" heatid="10192" lane="4" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WEZAB" name="Weteran Zabrze" nation="POL">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW. JANA  4A/4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-01" firstname="MACIEJ" gender="M" lastname="KUNICKI" nation="POL" athleteid="2635">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:31.87" resultid="2636" heatid="10107" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1162" points="383" swimtime="00:23:26.14" resultid="2637" heatid="10297" lane="8" entrytime="00:22:30.00" />
                <RESULT eventid="1292" points="401" swimtime="00:02:56.77" resultid="2638" heatid="10165" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="473" swimtime="00:01:15.28" resultid="2639" heatid="10239" lane="7" entrytime="00:01:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="DANIEL" gender="M" lastname="FECICA" nation="POL" athleteid="2640">
              <RESULTS>
                <RESULT eventid="1077" points="469" swimtime="00:00:43.90" resultid="2641" heatid="10102" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1324" points="737" swimtime="00:03:35.73" resultid="2642" heatid="10172" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="499" swimtime="00:00:48.19" resultid="2643" heatid="10187" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1654" points="628" swimtime="00:01:42.19" resultid="2644" heatid="10277" lane="8" entrytime="00:01:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="WIESŁAW" gender="M" lastname="KORNICKI" nation="POL" athleteid="2645">
              <RESULTS>
                <RESULT eventid="1077" points="578" swimtime="00:00:36.45" resultid="2646" heatid="10104" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1228" points="433" swimtime="00:01:22.40" resultid="2647" heatid="10150" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1574" status="DSQ" swimtime="00:00:31.60" resultid="2648" heatid="10250" lane="7" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="KRYSTYNA" gender="F" lastname="FECICA" nation="POL" athleteid="2649">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1141" points="797" swimtime="00:16:08.91" resultid="2650" heatid="10294" lane="1" entrytime="00:16:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.75" />
                    <SPLIT distance="200" swimtime="00:06:00.14" />
                    <SPLIT distance="300" swimtime="00:08:03.32" />
                    <SPLIT distance="400" swimtime="00:10:04.04" />
                    <SPLIT distance="500" swimtime="00:12:06.45" />
                    <SPLIT distance="600" swimtime="00:14:07.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1308" points="781" swimtime="00:04:05.83" resultid="2651" heatid="10168" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="531" swimtime="00:00:54.97" resultid="2652" heatid="10180" lane="2" entrytime="00:00:50.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1449" points="642" swimtime="00:03:47.03" resultid="2653" heatid="10209" lane="4" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Pierwszy wynik w kategorii" eventid="1525" points="494" swimtime="00:01:58.03" resultid="2654" heatid="10232" lane="3" entrytime="00:01:50.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1638" points="630" swimtime="00:01:56.33" resultid="2655" heatid="10272" lane="8" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="BERNARD" gender="M" lastname="POLOCZEK" nation="POL" athleteid="2656">
              <RESULTS>
                <RESULT eventid="1195" points="575" swimtime="00:00:42.41" resultid="2657" heatid="10135" lane="5" entrytime="00:00:43.22" />
                <RESULT eventid="1401" points="509" reactiontime="+70" swimtime="00:01:40.11" resultid="2658" heatid="10200" lane="3" entrytime="00:01:39.21" />
                <RESULT eventid="1606" points="457" reactiontime="+75" swimtime="00:03:46.50" resultid="2659" heatid="10262" lane="4" entrytime="00:03:47.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="EWALD" gender="M" lastname="BASTEK" nation="POL" athleteid="2660">
              <RESULTS>
                <RESULT eventid="1077" points="589" swimtime="00:00:40.68" resultid="2661" heatid="10102" lane="2" entrytime="00:00:43.50" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1162" points="622" swimtime="00:26:01.92" resultid="2662" heatid="10299" lane="7" entrytime="00:26:00.00" />
                <RESULT eventid="1195" points="614" swimtime="00:00:44.96" resultid="2663" heatid="10134" lane="4" entrytime="00:00:46.50" />
                <RESULT eventid="1228" points="594" swimtime="00:01:19.73" resultid="2664" heatid="10149" lane="2" entrytime="00:01:22.50" />
                <RESULT eventid="1401" points="522" reactiontime="+50" swimtime="00:01:45.00" resultid="2665" heatid="10199" lane="4" entrytime="00:01:48.00" />
                <RESULT eventid="1465" points="584" swimtime="00:03:05.04" resultid="2666" heatid="10216" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="591" swimtime="00:00:35.91" resultid="2667" heatid="10248" lane="3" entrytime="00:00:36.50" />
                <RESULT eventid="1686" points="577" swimtime="00:06:41.17" resultid="2668" heatid="10287" lane="2" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.09" />
                    <SPLIT distance="200" swimtime="00:03:21.38" />
                    <SPLIT distance="300" swimtime="00:05:03.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="RENATA" gender="F" lastname="BASTEK" nation="POL" athleteid="2669">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1061" points="981" swimtime="00:00:42.89" resultid="2670" heatid="10097" lane="8" entrytime="00:00:47.50" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1178" points="1040" swimtime="00:00:42.96" resultid="2671" heatid="10127" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="1161" swimtime="00:01:22.09" resultid="2672" heatid="10143" lane="7" entrytime="00:01:25.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1385" points="1069" reactiontime="+72" swimtime="00:01:38.99" resultid="2673" heatid="10194" lane="6" entrytime="00:01:45.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1558" points="1064" swimtime="00:00:36.90" resultid="2674" heatid="10243" lane="2" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="BEATA" gender="F" lastname="SULEWSKA" nation="POL" athleteid="2675">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1093" points="672" swimtime="00:02:48.67" resultid="2676" heatid="10113" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="563" swimtime="00:01:11.40" resultid="2677" heatid="10145" lane="4" entrytime="00:01:09.50" />
                <RESULT eventid="1308" points="616" swimtime="00:03:11.89" resultid="2678" heatid="10169" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1481" points="657" swimtime="00:06:05.99" resultid="2679" heatid="10225" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="200" swimtime="00:03:01.93" />
                    <SPLIT distance="300" swimtime="00:04:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="538" swimtime="00:01:20.77" resultid="2680" heatid="10233" lane="3" entrytime="00:01:22.00" />
                <RESULT eventid="1638" points="564" swimtime="00:01:30.91" resultid="2681" heatid="10273" lane="6" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="BARBARA" gender="F" lastname="BRENDLER" nation="POL" athleteid="2682">
              <RESULTS>
                <RESULT eventid="1061" points="236" swimtime="00:00:59.16" resultid="2683" heatid="10096" lane="6" entrytime="00:00:56.00" />
                <RESULT eventid="1212" points="418" swimtime="00:01:35.46" resultid="2684" heatid="10142" lane="1" entrytime="00:01:32.00" />
                <RESULT eventid="1449" points="380" swimtime="00:03:43.45" resultid="2685" heatid="10210" lane="5" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="486" swimtime="00:00:40.88" resultid="2686" heatid="10242" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="TADEUSZ" gender="M" lastname="STUCHLIK" nation="POL" athleteid="2687">
              <RESULTS>
                <RESULT eventid="1077" points="716" swimtime="00:00:29.80" resultid="2688" heatid="10109" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="1109" points="758" swimtime="00:02:29.55" resultid="2689" heatid="10122" lane="7" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="689" swimtime="00:00:31.72" resultid="2690" heatid="10140" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1401" points="728" reactiontime="+88" swimtime="00:01:07.50" resultid="2691" heatid="10205" lane="3" entrytime="00:01:06.50" />
                <RESULT eventid="1606" points="733" reactiontime="+93" swimtime="00:02:30.23" resultid="2692" heatid="10266" lane="5" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="GRAŻYNA" gender="F" lastname="KISZCZAK" nation="POL" athleteid="2693">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1061" points="879" swimtime="00:00:38.19" resultid="2694" heatid="10098" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1178" points="894" swimtime="00:00:39.88" resultid="2695" heatid="10129" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1385" points="824" reactiontime="+80" swimtime="00:01:30.12" resultid="2696" heatid="10196" lane="6" entrytime="00:01:28.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1481" points="591" swimtime="00:07:37.36" resultid="2697" heatid="10225" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.10" />
                    <SPLIT distance="200" swimtime="00:03:44.27" />
                    <SPLIT distance="300" swimtime="00:05:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="886" reactiontime="+73" swimtime="00:03:16.88" resultid="2698" heatid="10259" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="STANISŁAW" gender="M" lastname="KISZCZAK" nation="POL" athleteid="2699">
              <RESULTS>
                <RESULT eventid="1077" points="492" swimtime="00:00:40.32" resultid="2700" heatid="10103" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1574" points="633" swimtime="00:00:32.92" resultid="2701" heatid="10249" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="ULASZ" gender="M" lastname="SZANLI" nation="POL" athleteid="2702">
              <RESULTS>
                <RESULT eventid="1228" status="DSQ" swimtime="00:02:13.63" resultid="2703" heatid="10147" lane="4" entrytime="00:01:38.00" />
                <RESULT eventid="1574" points="246" swimtime="00:00:36.77" resultid="2704" heatid="10248" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="JAN" gender="M" lastname="BARUCHA" nation="POL" athleteid="2705">
              <RESULTS>
                <RESULT eventid="1077" points="334" swimtime="00:00:39.94" resultid="2706" heatid="10105" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1195" points="458" swimtime="00:00:39.70" resultid="2707" heatid="10137" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1574" points="508" swimtime="00:00:31.78" resultid="2708" heatid="10252" lane="6" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="WŁODZIMIERZ" gender="M" lastname="BOSOWSKI" nation="POL" athleteid="2709">
              <RESULTS>
                <RESULT eventid="1077" points="331" swimtime="00:00:46.02" resultid="2710" heatid="10103" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1195" points="266" swimtime="00:00:54.84" resultid="2711" heatid="10134" lane="1" entrytime="00:00:52.50" />
                <RESULT eventid="1401" points="207" reactiontime="+121" swimtime="00:02:15.13" resultid="2712" heatid="10200" lane="8" entrytime="00:01:48.00" />
                <RESULT eventid="1574" points="422" swimtime="00:00:37.69" resultid="2713" heatid="10248" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="JANINA" gender="F" lastname="BOSOWSKA" nation="POL" athleteid="2714">
              <RESULTS>
                <RESULT eventid="1061" status="DSQ" swimtime="00:01:01.63" resultid="2715" heatid="10096" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="1178" points="461" swimtime="00:00:53.23" resultid="2716" heatid="10127" lane="1" entrytime="00:00:54.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1352" points="449" swimtime="00:00:57.25" resultid="2717" heatid="10180" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="1558" points="401" swimtime="00:00:47.17" resultid="2718" heatid="10242" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+83" swimtime="00:02:27.40" resultid="2724" heatid="10160" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2687" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2640" number="2" />
                    <RELAYPOSITION athleteid="2645" number="3" />
                    <RELAYPOSITION athleteid="2699" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+76" swimtime="00:02:42.08" resultid="2725" heatid="10160" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2656" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2660" number="2" />
                    <RELAYPOSITION athleteid="2635" number="3" />
                    <RELAYPOSITION athleteid="2709" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1433" swimtime="00:02:18.70" resultid="2727" heatid="10207" lane="3" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2705" number="1" />
                    <RELAYPOSITION athleteid="2709" number="2" />
                    <RELAYPOSITION athleteid="2645" number="3" />
                    <RELAYPOSITION athleteid="2699" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="4">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1244" reactiontime="+80" swimtime="00:02:43.96" resultid="2723" heatid="10159" lane="7" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2693" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2649" number="2" />
                    <RELAYPOSITION athleteid="2675" number="3" />
                    <RELAYPOSITION athleteid="2669" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1417" swimtime="00:02:42.95" resultid="2726" heatid="10206" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2682" number="1" />
                    <RELAYPOSITION athleteid="2714" number="2" />
                    <RELAYPOSITION athleteid="2693" number="3" />
                    <RELAYPOSITION athleteid="2669" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1125" swimtime="00:02:25.21" resultid="2719" heatid="10124" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2669" number="1" />
                    <RELAYPOSITION athleteid="2660" number="2" />
                    <RELAYPOSITION athleteid="2640" number="3" />
                    <RELAYPOSITION athleteid="2693" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:33.09" resultid="2721" heatid="10124" lane="7" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2705" number="1" />
                    <RELAYPOSITION athleteid="2714" number="2" />
                    <RELAYPOSITION athleteid="2682" number="3" />
                    <RELAYPOSITION athleteid="2645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:35.61" resultid="2722" heatid="10124" lane="1" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2649" number="1" />
                    <RELAYPOSITION athleteid="2709" number="2" />
                    <RELAYPOSITION athleteid="2656" number="3" />
                    <RELAYPOSITION athleteid="2675" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="9">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+82" swimtime="00:02:56.54" resultid="2720" heatid="10268" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2693" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="2640" number="2" />
                    <RELAYPOSITION athleteid="2660" number="3" />
                    <RELAYPOSITION athleteid="2669" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="10">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+74" swimtime="00:02:50.64" resultid="2728" heatid="10268" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2656" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2649" number="2" />
                    <RELAYPOSITION athleteid="2645" number="3" />
                    <RELAYPOSITION athleteid="2675" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" name="TS MASTERS WISŁA KRAKÓW" nation="POL" shortname="WISŁA KRAKÓW">
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="2748">
              <RESULTS>
                <RESULT eventid="1109" points="1014" swimtime="00:04:01.47" resultid="2750" heatid="10116" lane="2" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:03.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="823" swimtime="00:04:19.97" resultid="2751" heatid="10170" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:05.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="595" swimtime="00:00:53.53" resultid="2752" heatid="10184" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1574" points="627" swimtime="00:00:38.72" resultid="2754" heatid="10247" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1686" points="758" swimtime="00:07:31.95" resultid="2755" heatid="10287" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.49" />
                    <SPLIT distance="200" swimtime="00:03:38.11" />
                    <SPLIT distance="300" swimtime="00:05:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="639" swimtime="00:01:29.80" resultid="2756" heatid="10148" lane="6" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Janusz" gender="M" lastname="Konstanty" nation="POL" athleteid="2757">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2758" heatid="10118" lane="1" entrytime="00:03:15.00" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="2759" heatid="10137" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="2760" heatid="10202" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1606" status="DNS" swimtime="00:00:00.00" resultid="2761" heatid="10263" lane="4" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="2762">
              <RESULTS>
                <RESULT eventid="1093" points="524" swimtime="00:02:52.28" resultid="2763" heatid="10113" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="606" swimtime="00:00:35.20" resultid="2764" heatid="10130" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1385" points="640" reactiontime="+63" swimtime="00:01:14.33" resultid="2765" heatid="10197" lane="5" entrytime="00:01:16.00" />
                <RESULT eventid="1590" points="556" reactiontime="+63" swimtime="00:02:44.86" resultid="2766" heatid="10260" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Pawel" gender="M" lastname="Lesiakowski" nation="POL" athleteid="2767">
              <RESULTS>
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="2768" heatid="10187" lane="7" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="2769">
              <RESULTS>
                <RESULT eventid="1162" points="357" swimtime="00:23:06.00" resultid="2770" heatid="10298" lane="1" entrytime="00:24:00.00" />
                <RESULT eventid="1465" points="436" swimtime="00:02:27.19" resultid="2771" heatid="10220" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="594" swimtime="00:01:00.23" resultid="2772" heatid="10153" lane="4" entrytime="00:01:05.00" />
                <RESULT eventid="1574" points="615" swimtime="00:00:27.12" resultid="2773" heatid="10254" lane="5" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MARZE" name="Masters Rzeszów" nation="POL">
          <CONTACT city="Rzeszów" email="wieslawcieklinski@wp.pl" name="Ciekliński" phone="602682904" street="Jagiellońska 7/3" zip="35-025" />
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="2775">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:39.47" resultid="2776" heatid="10103" lane="4" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2777" heatid="10117" lane="4" entrytime="00:03:15.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="560" swimtime="00:01:11.20" resultid="2778" heatid="10151" lane="6" entrytime="00:01:11.50" entrycourse="LCM" />
                <RESULT eventid="1465" points="499" swimtime="00:02:46.06" resultid="2779" heatid="10217" lane="2" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" status="DSQ" swimtime="00:00:32.07" resultid="2780" heatid="10251" lane="2" entrytime="00:00:31.20" entrycourse="LCM" />
                <RESULT eventid="1686" points="492" swimtime="00:06:02.52" resultid="2781" heatid="10289" lane="8" entrytime="00:06:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="200" swimtime="00:02:58.69" />
                    <SPLIT distance="300" swimtime="00:04:32.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" name="Ks Warta Poznań" nation="POL" region="WIE" shortname="Warta Poznań">
          <CONTACT city="Poznań" email="j.thiem@glos.com" name="Thiem Jacek" phone="502499565" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1965-05-08" firstname="ANNA" gender="F" lastname="KOTECKA" nation="POL" athleteid="2783">
              <RESULTS>
                <RESULT eventid="1141" points="486" swimtime="00:13:04.13" resultid="2784" heatid="10294" lane="5" entrytime="00:13:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.07" />
                    <SPLIT distance="200" swimtime="00:03:02.77" />
                    <SPLIT distance="300" swimtime="00:04:43.98" />
                    <SPLIT distance="400" swimtime="00:06:24.58" />
                    <SPLIT distance="500" swimtime="00:08:05.23" />
                    <SPLIT distance="600" swimtime="00:09:45.30" />
                    <SPLIT distance="700" swimtime="00:11:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="392" swimtime="00:00:45.59" resultid="2785" heatid="10127" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1212" points="462" swimtime="00:01:22.15" resultid="2786" heatid="10143" lane="2" entrytime="00:01:22.00" />
                <RESULT eventid="1385" points="460" reactiontime="+50" swimtime="00:01:34.69" resultid="2787" heatid="10195" lane="7" entrytime="00:01:38.00" />
                <RESULT eventid="1449" points="443" swimtime="00:03:00.92" resultid="2788" heatid="10211" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="494" reactiontime="+67" swimtime="00:03:25.38" resultid="2789" heatid="10259" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="468" swimtime="00:06:17.11" resultid="2790" heatid="10284" lane="7" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.97" />
                    <SPLIT distance="200" swimtime="00:03:02.71" />
                    <SPLIT distance="300" swimtime="00:04:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="JACEK" gender="M" lastname="THIEM" nation="POL" athleteid="2791">
              <RESULTS>
                <RESULT eventid="1162" points="339" swimtime="00:26:10.88" resultid="2792" heatid="10299" lane="3" entrytime="00:25:00.00" />
                <RESULT eventid="1292" points="474" swimtime="00:03:12.69" resultid="2793" heatid="10165" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="414" swimtime="00:02:46.74" resultid="2794" heatid="10217" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="393" swimtime="00:01:26.17" resultid="2795" heatid="10237" lane="7" entrytime="00:01:28.00" />
                <RESULT eventid="1686" points="352" swimtime="00:06:19.86" resultid="2796" heatid="10288" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                    <SPLIT distance="200" swimtime="00:03:11.16" />
                    <SPLIT distance="300" swimtime="00:04:50.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="DARIUSZ" gender="M" lastname="JANYGA" nation="POL" athleteid="2797">
              <RESULTS>
                <RESULT eventid="1195" points="610" swimtime="00:00:34.02" resultid="2798" heatid="10138" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1228" points="558" swimtime="00:01:06.52" resultid="2799" heatid="10155" lane="8" entrytime="00:01:03.50" />
                <RESULT eventid="1401" points="629" reactiontime="+84" swimtime="00:01:15.91" resultid="2800" heatid="10204" lane="1" entrytime="00:01:14.50" />
                <RESULT eventid="1574" points="584" swimtime="00:00:29.34" resultid="2801" heatid="10254" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="1606" points="582" reactiontime="+95" swimtime="00:02:48.78" resultid="2802" heatid="10265" lane="7" entrytime="00:02:47.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-11-17" firstname="ZBIGNIEW" gender="M" lastname="LIBER" nation="POL" athleteid="2803">
              <RESULTS>
                <RESULT eventid="1369" points="190" swimtime="00:00:55.98" resultid="2804" heatid="10184" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1574" points="125" swimtime="00:00:50.66" resultid="2805" heatid="10247" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="PAWEŁ" gender="M" lastname="OLSZEWSKI" nation="POL" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1228" points="807" swimtime="00:01:01.09" resultid="2807" heatid="10156" lane="6" entrytime="00:01:01.50" />
                <RESULT eventid="1465" points="762" swimtime="00:02:16.06" resultid="2808" heatid="10222" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="668" swimtime="00:00:29.02" resultid="2809" heatid="10254" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1686" points="749" swimtime="00:04:55.49" resultid="2810" heatid="10292" lane="8" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="200" swimtime="00:02:25.41" />
                    <SPLIT distance="300" swimtime="00:03:40.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="PRZEMYSŁAW" gender="M" lastname="WARACZEWSKI" nation="POL" athleteid="2811">
              <RESULTS>
                <RESULT eventid="1195" points="464" swimtime="00:00:39.54" resultid="2812" heatid="10135" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1324" points="569" swimtime="00:03:14.52" resultid="2813" heatid="10174" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="612" swimtime="00:00:37.91" resultid="2814" heatid="10187" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1574" points="463" swimtime="00:00:32.78" resultid="2815" heatid="10250" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1654" points="550" swimtime="00:01:28.78" resultid="2816" heatid="10278" lane="7" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04514" name="UKS 307" nation="POL" region="MAZ">
          <CONTACT name="ILCZYSZYN" />
          <ATHLETES>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="Ziółkowski" nation="POL" athleteid="2820">
              <RESULTS>
                <RESULT eventid="1228" points="520" swimtime="00:01:03.95" resultid="2821" heatid="10154" lane="5" entrytime="00:01:03.90" />
                <RESULT eventid="1465" points="494" swimtime="00:02:26.90" resultid="2822" heatid="10219" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="389" swimtime="00:01:18.14" resultid="2823" heatid="10238" lane="2" entrytime="00:01:17.00" />
                <RESULT eventid="1574" points="497" swimtime="00:00:29.22" resultid="2824" heatid="10254" lane="1" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-13" firstname="Krzysztof" gender="M" lastname="Ilczyszyn" nation="POL" athleteid="2825">
              <RESULTS>
                <RESULT eventid="1228" points="478" swimtime="00:01:04.75" resultid="2826" heatid="10154" lane="4" entrytime="00:01:03.90" />
                <RESULT eventid="1465" points="394" swimtime="00:02:32.19" resultid="2827" heatid="10219" lane="7" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="370" swimtime="00:01:17.55" resultid="2828" heatid="10238" lane="6" entrytime="00:01:17.00" />
                <RESULT eventid="1574" status="DSQ" swimtime="00:00:29.65" resultid="2829" heatid="10253" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STPOZ" name="Start Poznań" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1967-07-02" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="2830">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2832" heatid="10121" lane="5" entrytime="00:02:31.00" />
                <RESULT eventid="1228" points="797" swimtime="00:00:59.07" resultid="2833" heatid="10157" lane="2" entrytime="00:00:59.30" />
                <RESULT eventid="1465" points="728" swimtime="00:02:16.23" resultid="2834" heatid="10214" lane="6" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1497" points="752" swimtime="00:05:34.05" resultid="2835" heatid="10231" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="200" swimtime="00:02:46.47" />
                    <SPLIT distance="300" swimtime="00:04:22.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="722" swimtime="00:00:27.34" resultid="2836" heatid="10256" lane="4" entrytime="00:00:26.80" />
                <RESULT eventid="1686" points="728" swimtime="00:04:52.07" resultid="2837" heatid="10292" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                    <SPLIT distance="200" swimtime="00:02:24.14" />
                    <SPLIT distance="300" swimtime="00:03:38.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="3823">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="3824" heatid="10106" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3825" heatid="10120" lane="8" entrytime="00:02:50.00" />
                <RESULT eventid="1195" points="616" swimtime="00:00:32.92" resultid="3826" heatid="10138" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1228" status="DSQ" swimtime="00:01:00.40" resultid="3827" heatid="10154" lane="8" entrytime="00:01:05.00" />
                <RESULT eventid="1401" points="649" reactiontime="+83" swimtime="00:01:10.13" resultid="3828" heatid="10204" lane="7" entrytime="00:01:12.00" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="3829" heatid="10221" lane="5" entrytime="00:02:22.00" />
                <RESULT eventid="1574" points="668" swimtime="00:00:27.93" resultid="3830" heatid="10252" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1606" status="DNS" swimtime="00:00:00.00" resultid="3831" heatid="10265" lane="3" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ENZGO" name="UKS Energetyk Zgorzelec" nation="POL" shortname="Energetyk Zgorzelec">
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="3076">
              <RESULTS>
                <RESULT eventid="1077" points="199" swimtime="00:00:54.47" resultid="3078" heatid="10101" lane="8" entrytime="00:00:57.00" />
                <RESULT eventid="1109" points="330" swimtime="00:04:10.02" resultid="3079" heatid="10115" lane="3" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="341" swimtime="00:00:50.48" resultid="3080" heatid="10133" lane="5" entrytime="00:00:53.00" />
                <RESULT eventid="1292" points="262" swimtime="00:04:46.70" resultid="3081" heatid="10163" lane="2" entrytime="00:04:29.00" />
                <RESULT eventid="1401" points="340" reactiontime="+86" swimtime="00:01:54.45" resultid="3082" heatid="10199" lane="3" entrytime="00:01:52.00" />
                <RESULT eventid="1497" points="310" swimtime="00:09:12.13" resultid="3083" heatid="10227" lane="6" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.06" />
                    <SPLIT distance="200" swimtime="00:04:32.51" />
                    <SPLIT distance="300" swimtime="00:07:13.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="193" swimtime="00:02:11.52" resultid="3084" heatid="10235" lane="7" entrytime="00:02:05.00" />
                <RESULT eventid="1606" points="370" reactiontime="+83" swimtime="00:04:03.06" resultid="3085" heatid="10262" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:00.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WPOZO" name="Zgiersko - Łęczyckie WOPR - Ozorków" nation="POL" region="LOD" shortname="WOPR Ozorków">
          <CONTACT city="OZORKÓW" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁODZK" street="Lotnicza 1 a" zip="95-035" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-22" firstname="ROMAN" gender="M" lastname="WICZEL" nation="POL" license="M0180520003" athleteid="3087">
              <RESULTS>
                <RESULT eventid="1324" points="652" swimtime="00:03:32.74" resultid="3088" heatid="10173" lane="3" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="791" swimtime="00:00:39.13" resultid="3089" heatid="10188" lane="6" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1654" points="717" swimtime="00:01:30.98" resultid="3090" heatid="10278" lane="6" entrytime="00:01:30.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-03-14" firstname="ALEKSANDER" gender="M" lastname="OSSOWSKI" nation="POL" license="M0180520001" athleteid="3091">
              <RESULTS>
                <RESULT eventid="1162" points="449" swimtime="00:26:34.76" resultid="3092" heatid="10300" lane="4" entrytime="00:27:00.00" entrycourse="LCM" />
                <RESULT eventid="1195" points="567" swimtime="00:00:40.40" resultid="3093" heatid="10136" lane="3" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1401" points="500" reactiontime="+82" swimtime="00:01:32.70" resultid="3094" heatid="10201" lane="7" entrytime="00:01:31.00" entrycourse="LCM" />
                <RESULT eventid="1497" points="402" swimtime="00:07:51.75" resultid="3095" heatid="10228" lane="7" entrytime="00:07:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.37" />
                    <SPLIT distance="200" swimtime="00:04:06.34" />
                    <SPLIT distance="300" swimtime="00:06:15.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="426" reactiontime="+89" swimtime="00:03:35.04" resultid="3096" heatid="10263" lane="7" entrytime="00:03:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-20" firstname="BOGDAN" gender="M" lastname="WĄSIK" nation="POL" license="M0180520002" athleteid="3097">
              <RESULTS>
                <RESULT eventid="1324" points="568" swimtime="00:03:18.85" resultid="3098" heatid="10174" lane="4" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="555" swimtime="00:00:40.41" resultid="3099" heatid="10188" lane="5" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1654" points="536" swimtime="00:01:31.41" resultid="3100" heatid="10278" lane="3" entrytime="00:01:28.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-13" firstname="MIROSŁAWA" gender="F" lastname="RAJTAR" nation="POL" license="M0180510004" athleteid="3101">
              <RESULTS>
                <RESULT eventid="1558" points="570" swimtime="00:00:37.41" resultid="3105" heatid="10243" lane="8" entrytime="00:00:37.60" entrycourse="LCM" />
                <RESULT eventid="1061" points="403" swimtime="00:00:45.43" resultid="3102" heatid="10097" lane="3" entrytime="00:00:43.60" entrycourse="LCM" />
                <RESULT eventid="1178" points="514" swimtime="00:00:46.25" resultid="3103" heatid="10127" lane="6" entrytime="00:00:46.60" entrycourse="LCM" />
                <RESULT eventid="1385" points="493" swimtime="00:01:43.73" resultid="3104" heatid="10194" lane="4" entrytime="00:01:40.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="URSZULA" gender="F" lastname="MRÓZ" nation="POL" license="M0180510002" athleteid="3106">
              <RESULTS>
                <RESULT eventid="1061" points="625" swimtime="00:00:38.56" resultid="3107" heatid="10098" lane="5" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1178" status="DSQ" swimtime="00:00:40.46" resultid="3108" heatid="10129" lane="2" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1385" points="593" reactiontime="+80" swimtime="00:01:31.90" resultid="3109" heatid="10195" lane="5" entrytime="00:01:31.00" entrycourse="LCM" />
                <RESULT eventid="1525" points="489" swimtime="00:01:33.29" resultid="3110" heatid="10233" lane="2" entrytime="00:01:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="EWA" gender="F" lastname="STĘPIEŃ" nation="POL" license="M0180510003" athleteid="3111">
              <RESULTS>
                <RESULT eventid="1093" points="649" swimtime="00:03:08.41" resultid="3112" heatid="10112" lane="2" entrytime="00:03:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="644" swimtime="00:01:15.30" resultid="3113" heatid="10144" lane="6" entrytime="00:01:16.00" entrycourse="LCM" />
                <RESULT eventid="1308" points="617" swimtime="00:03:29.60" resultid="3114" heatid="10169" lane="7" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1352" points="840" swimtime="00:00:40.17" resultid="3115" heatid="10182" lane="8" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1558" points="697" swimtime="00:00:32.86" resultid="3116" heatid="10244" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1638" points="771" swimtime="00:01:30.88" resultid="3117" heatid="10272" lane="5" entrytime="00:01:32.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="TOMASZ" gender="M" lastname="NIEDZWIEDZ" nation="POL" license="M01805200" athleteid="3118">
              <RESULTS>
                <RESULT eventid="1109" points="320" swimtime="00:03:37.08" resultid="3119" heatid="10115" lane="4" entrytime="00:03:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="246" swimtime="00:03:59.58" resultid="3120" heatid="10164" lane="1" entrytime="00:04:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="309" swimtime="00:07:47.81" resultid="3121" heatid="10227" lane="5" entrytime="00:08:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.47" />
                    <SPLIT distance="200" swimtime="00:03:55.66" />
                    <SPLIT distance="300" swimtime="00:06:04.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="207" swimtime="00:01:46.77" resultid="3122" heatid="10236" lane="8" entrytime="00:01:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="WŁODZIMIERZ" gender="M" lastname="PRZYTULSKI" nation="POL" license="M0180520005" athleteid="3123">
              <RESULTS>
                <RESULT eventid="1077" points="659" swimtime="00:00:32.26" resultid="3124" heatid="10107" lane="7" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3125" heatid="10118" lane="4" entrytime="00:03:02.00" entrycourse="LCM" />
                <RESULT eventid="1195" points="654" swimtime="00:00:36.75" resultid="3126" heatid="10138" lane="7" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="3127" heatid="10165" lane="7" entrytime="00:03:10.00" entrycourse="LCM" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="3128" heatid="10202" lane="3" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="581" swimtime="00:02:37.88" resultid="3129" heatid="10219" lane="5" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="3130" heatid="10237" lane="4" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="1606" points="525" reactiontime="+88" swimtime="00:03:06.66" resultid="3131" heatid="10264" lane="7" entrytime="00:03:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="MAŁGORZATA" gender="F" lastname="ŚCIBIOREK" nation="POL" license="M01805100" athleteid="3132">
              <RESULTS>
                <RESULT eventid="1061" points="746" swimtime="00:00:32.70" resultid="3133" heatid="10099" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1093" points="652" swimtime="00:02:50.39" resultid="3134" heatid="10113" lane="1" entrytime="00:02:51.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="585" swimtime="00:00:37.56" resultid="3135" heatid="10130" lane="6" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1385" points="561" reactiontime="+90" swimtime="00:01:20.86" resultid="3136" heatid="10197" lane="8" entrytime="00:01:21.00" entrycourse="LCM" />
                <RESULT eventid="1670" points="536" swimtime="00:05:34.74" resultid="3137" heatid="10285" lane="8" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="200" swimtime="00:02:41.71" />
                    <SPLIT distance="300" swimtime="00:04:08.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="TOMASZ" gender="M" lastname="CAJDLER" nation="POL" license="M0180520006" athleteid="3138">
              <RESULTS>
                <RESULT eventid="1228" points="450" swimtime="00:01:14.20" resultid="3139" heatid="10151" lane="1" entrytime="00:01:13.00" entrycourse="LCM" />
                <RESULT eventid="1369" points="487" swimtime="00:00:40.92" resultid="3140" heatid="10188" lane="8" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1574" points="492" swimtime="00:00:32.12" resultid="3141" heatid="10250" lane="4" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1654" points="349" swimtime="00:01:43.33" resultid="3142" heatid="10277" lane="5" entrytime="00:01:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Z - Ł WOPR" number="1">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+82" swimtime="00:02:30.19" resultid="3147" heatid="10160" lane="5" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3091" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3087" number="2" />
                    <RELAYPOSITION athleteid="3123" number="3" />
                    <RELAYPOSITION athleteid="3138" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Z - Ł WOPR" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1244" reactiontime="+74" swimtime="00:02:35.88" resultid="3145" heatid="10159" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3106" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3111" number="2" />
                    <RELAYPOSITION athleteid="3132" number="3" />
                    <RELAYPOSITION athleteid="3101" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1417" swimtime="00:02:20.78" resultid="3146" heatid="10206" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3132" number="1" />
                    <RELAYPOSITION athleteid="3101" number="2" />
                    <RELAYPOSITION athleteid="3106" number="3" />
                    <RELAYPOSITION athleteid="3111" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Z - Ł WOPR" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:11.07" resultid="3143" heatid="10125" lane="8" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3111" number="1" />
                    <RELAYPOSITION athleteid="3091" number="2" />
                    <RELAYPOSITION athleteid="3132" number="3" />
                    <RELAYPOSITION athleteid="3123" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+77" swimtime="00:02:29.93" resultid="3144" heatid="10269" lane="1" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3123" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3111" number="2" />
                    <RELAYPOSITION athleteid="3132" number="3" />
                    <RELAYPOSITION athleteid="3091" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASTKRAŚ" name="Masters Kraśnik" nation="POL" region="LBL">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="3158">
              <RESULTS>
                <RESULT eventid="1324" points="461" swimtime="00:03:14.60" resultid="3159" heatid="10174" lane="8" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="377" swimtime="00:00:40.82" resultid="3160" heatid="10188" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1654" points="411" swimtime="00:01:30.35" resultid="3161" heatid="10278" lane="1" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="3162">
              <RESULTS>
                <RESULT eventid="1077" points="366" swimtime="00:00:38.75" resultid="3163" heatid="10103" lane="3" entrytime="00:00:38.57" />
                <RESULT eventid="1109" points="362" swimtime="00:03:28.32" resultid="3164" heatid="10118" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="485" swimtime="00:00:38.97" resultid="3165" heatid="10137" lane="7" entrytime="00:00:39.13" />
                <RESULT eventid="1228" points="457" swimtime="00:01:13.82" resultid="3166" heatid="10152" lane="8" entrytime="00:01:10.00" />
                <RESULT eventid="1401" points="474" reactiontime="+81" swimtime="00:01:26.14" resultid="3167" heatid="10201" lane="5" entrytime="00:01:27.86" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="3168" heatid="10218" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="362" swimtime="00:00:35.59" resultid="3169" heatid="10251" lane="4" entrytime="00:00:30.70" />
                <RESULT eventid="1606" points="180" reactiontime="+106" swimtime="00:04:23.46" resultid="3170" heatid="10263" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-17" firstname="Jacek" gender="M" lastname="Janik" nation="POL" athleteid="3171">
              <RESULTS>
                <RESULT eventid="1077" points="195" swimtime="00:00:47.23" resultid="3172" heatid="10103" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1228" points="325" swimtime="00:01:19.62" resultid="3173" heatid="10149" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1324" points="300" swimtime="00:03:49.85" resultid="3174" heatid="10171" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="288" swimtime="00:00:46.47" resultid="3175" heatid="10186" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1465" points="276" swimtime="00:03:08.04" resultid="3176" heatid="10216" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="274" swimtime="00:00:37.76" resultid="3177" heatid="10249" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1654" points="274" swimtime="00:01:45.80" resultid="3178" heatid="10276" lane="8" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:44.46" resultid="3180" heatid="10101" lane="5" entrytime="00:00:46.02" />
                <RESULT eventid="1109" points="273" swimtime="00:03:58.49" resultid="3181" heatid="10115" lane="5" entrytime="00:03:52.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="338" swimtime="00:00:45.79" resultid="3182" heatid="10135" lane="8" entrytime="00:00:46.20" />
                <RESULT eventid="1401" points="282" reactiontime="+94" swimtime="00:01:43.00" resultid="3183" heatid="10200" lane="1" entrytime="00:01:47.20" />
                <RESULT eventid="1542" points="179" swimtime="00:01:54.21" resultid="3184" heatid="10235" lane="5" entrytime="00:01:52.00" />
                <RESULT eventid="1606" points="259" reactiontime="+107" swimtime="00:03:56.25" resultid="3185" heatid="10262" lane="5" entrytime="00:03:52.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="3186">
              <RESULTS>
                <RESULT eventid="1109" points="332" swimtime="00:03:52.60" resultid="3187" heatid="10115" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="179" swimtime="00:04:47.27" resultid="3188" heatid="10163" lane="7" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="446" swimtime="00:03:50.97" resultid="3189" heatid="10171" lane="6" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="247" swimtime="00:03:44.84" resultid="3190" heatid="10215" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="282" swimtime="00:08:50.64" resultid="3191" heatid="10227" lane="2" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:11.18" />
                    <SPLIT distance="200" swimtime="00:04:41.35" />
                    <SPLIT distance="300" swimtime="00:06:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="205" reactiontime="+121" swimtime="00:04:34.41" resultid="3192" heatid="10262" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="189" swimtime="00:08:33.84" resultid="3193" heatid="10286" lane="2" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:06.24" />
                    <SPLIT distance="200" swimtime="00:04:20.92" />
                    <SPLIT distance="300" swimtime="00:06:34.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="3194">
              <RESULTS>
                <RESULT eventid="1077" points="211" swimtime="00:00:47.14" resultid="3195" heatid="10101" lane="3" entrytime="00:00:46.30" />
                <RESULT eventid="1195" points="244" swimtime="00:00:51.05" resultid="3196" heatid="10134" lane="7" entrytime="00:00:50.20" />
                <RESULT eventid="1292" points="102" swimtime="00:05:24.98" resultid="3197" heatid="10163" lane="1" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:24.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="251" swimtime="00:00:52.63" resultid="3198" heatid="10185" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1654" points="294" swimtime="00:01:51.70" resultid="3199" heatid="10275" lane="2" entrytime="00:01:58.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GDMAS" name="Gdynia Masters" nation="POL">
          <CONTACT name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1061" points="413" swimtime="00:00:44.28" resultid="3202" heatid="10097" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1141" points="389" swimtime="00:14:23.01" resultid="3203" heatid="10294" lane="6" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.79" />
                    <SPLIT distance="200" swimtime="00:03:23.94" />
                    <SPLIT distance="300" swimtime="00:05:14.84" />
                    <SPLIT distance="400" swimtime="00:07:06.51" />
                    <SPLIT distance="500" swimtime="00:08:58.02" />
                    <SPLIT distance="600" swimtime="00:10:49.13" />
                    <SPLIT distance="700" swimtime="00:12:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="466" swimtime="00:00:44.61" resultid="3204" heatid="10128" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1212" points="463" swimtime="00:01:24.06" resultid="3205" heatid="10142" lane="3" entrytime="00:01:27.00" />
                <RESULT eventid="1449" points="410" swimtime="00:03:12.86" resultid="3206" heatid="10211" lane="6" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="511" swimtime="00:00:36.44" resultid="3207" heatid="10243" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1670" points="422" swimtime="00:06:52.02" resultid="3208" heatid="10283" lane="4" entrytime="00:06:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.35" />
                    <SPLIT distance="200" swimtime="00:03:22.21" />
                    <SPLIT distance="300" swimtime="00:05:10.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1195" points="526" swimtime="00:00:48.95" resultid="3210" heatid="10133" lane="2" entrytime="00:00:57.00" />
                <RESULT eventid="1324" points="597" swimtime="00:03:59.18" resultid="3211" heatid="10171" lane="3" entrytime="00:03:53.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="597" swimtime="00:00:47.61" resultid="3212" heatid="10185" lane="5" entrytime="00:00:46.49" />
                <RESULT eventid="1654" status="DSQ" swimtime="00:01:54.35" resultid="3213" heatid="10276" lane="1" entrytime="00:01:44.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="3214">
              <RESULTS>
                <RESULT eventid="1077" points="408" swimtime="00:00:45.99" resultid="3215" heatid="10101" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1109" points="481" swimtime="00:03:57.09" resultid="3216" heatid="10116" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="517" swimtime="00:00:47.60" resultid="3217" heatid="10134" lane="5" entrytime="00:00:47.00" />
                <RESULT eventid="1324" points="567" swimtime="00:03:55.39" resultid="3218" heatid="10171" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="698" swimtime="00:00:43.09" resultid="3219" heatid="10187" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1465" points="389" swimtime="00:03:31.77" resultid="3220" heatid="10216" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="499" swimtime="00:00:38.00" resultid="3221" heatid="10248" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1654" points="611" swimtime="00:01:43.17" resultid="3222" heatid="10276" lane="7" entrytime="00:01:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="3223">
              <RESULTS>
                <RESULT eventid="1109" points="398" swimtime="00:03:38.92" resultid="3224" heatid="10116" lane="6" entrytime="00:03:40.00" />
                <RESULT eventid="1324" points="492" swimtime="00:03:43.54" resultid="3225" heatid="10172" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="344" swimtime="00:00:48.88" resultid="3226" heatid="10186" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1497" points="399" swimtime="00:07:52.68" resultid="3227" heatid="10228" lane="2" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.62" />
                    <SPLIT distance="200" swimtime="00:04:05.99" />
                    <SPLIT distance="300" swimtime="00:06:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="422" swimtime="00:01:45.26" resultid="3228" heatid="10276" lane="5" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGOR" name="MASTERS Gorzów Wlkp." nation="POL" region="LBS" shortname="MASTERS Gorzów">
          <CONTACT city="Kłodawa" email="mastersgorzow@onet.eu" name="Marek Wojciechowicz" phone="602891603" state="LUB" street="Skalna 2" zip="66-415" />
          <ATHLETES>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="Wojciechowicz" nation="POL" license="500604200002" athleteid="3230">
              <RESULTS>
                <RESULT eventid="1109" points="597" swimtime="00:02:41.95" resultid="3231" heatid="10119" lane="4" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="499" swimtime="00:21:26.89" resultid="3232" heatid="10297" lane="5" entrytime="00:21:00.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="608" swimtime="00:01:03.04" resultid="3233" heatid="10156" lane="2" entrytime="00:01:01.50" entrycourse="LCM" />
                <RESULT eventid="1465" points="579" swimtime="00:02:22.03" resultid="3234" heatid="10222" lane="5" entrytime="00:02:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="671" swimtime="00:00:27.89" resultid="3235" heatid="10255" lane="4" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="1686" points="507" swimtime="00:05:15.03" resultid="3236" heatid="10291" lane="6" entrytime="00:05:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:02:33.54" />
                    <SPLIT distance="300" swimtime="00:03:55.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" license="500604200001" athleteid="3237">
              <RESULTS>
                <RESULT eventid="1162" points="335" swimtime="00:28:15.75" resultid="3238" heatid="10300" lane="7" entrytime="00:29:00.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="332" swimtime="00:01:24.71" resultid="3239" heatid="10148" lane="5" entrytime="00:01:25.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="290" swimtime="00:03:19.00" resultid="3240" heatid="10216" lane="6" entrytime="00:03:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="378" swimtime="00:00:36.10" resultid="3241" heatid="10248" lane="8" entrytime="00:00:37.50" entrycourse="LCM" />
                <RESULT eventid="1686" points="333" swimtime="00:06:52.93" resultid="3242" heatid="10287" lane="1" entrytime="00:06:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.05" />
                    <SPLIT distance="200" swimtime="00:03:17.43" />
                    <SPLIT distance="300" swimtime="00:05:06.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NARUD" name="Naprzód RYDUŁTOWY" nation="POL">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK  Marian" phone="530556313" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="RUDOLF" gender="M" lastname="BUGLA" nation="POL" athleteid="3244">
              <RESULTS>
                <RESULT eventid="1077" points="225" swimtime="00:00:56.05" resultid="3245" heatid="10101" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1109" points="291" swimtime="00:04:40.34" resultid="3246" heatid="10115" lane="7" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="272" swimtime="00:00:58.92" resultid="3247" heatid="10133" lane="8" entrytime="00:00:58.00" />
                <RESULT eventid="1292" points="232" swimtime="00:05:14.86" resultid="3248" heatid="10163" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="279" reactiontime="+88" swimtime="00:02:09.39" resultid="3249" heatid="10199" lane="1" entrytime="00:02:00.00" />
                <RESULT eventid="1497" points="247" swimtime="00:10:30.85" resultid="3250" heatid="10227" lane="7" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:28.95" />
                    <SPLIT distance="200" swimtime="00:05:09.97" />
                    <SPLIT distance="300" swimtime="00:07:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="203" swimtime="00:02:16.96" resultid="3251" heatid="10235" lane="3" entrytime="00:02:00.00" />
                <RESULT eventid="1606" points="317" reactiontime="+97" swimtime="00:04:31.64" resultid="3252" heatid="10262" lane="7" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZKS DRZ" name="ZKS Drzonków" nation="POL" region="ZG">
          <CONTACT city="ŁĘŻYCA" email="piotrbarta@o2.pl" name="BARTA PIOTR" phone="602347348" state="LUB" street="ODRZAŃSKA 21" zip="66-016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="PIOTR" gender="M" lastname="BARTA" nation="POL" athleteid="3254">
              <RESULTS>
                <RESULT eventid="1109" points="681" swimtime="00:02:34.97" resultid="3255" heatid="10120" lane="6" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="746" swimtime="00:02:45.76" resultid="3256" heatid="10177" lane="7" entrytime="00:02:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="641" swimtime="00:00:34.21" resultid="3257" heatid="10191" lane="7" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1497" points="646" swimtime="00:05:39.29" resultid="3258" heatid="10230" lane="6" entrytime="00:06:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="200" swimtime="00:02:48.76" />
                    <SPLIT distance="300" swimtime="00:04:20.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="675" swimtime="00:01:16.57" resultid="3259" heatid="10275" lane="4" entrytime="00:01:45.00" entrycourse="LCM" />
                <RESULT eventid="1686" points="602" swimtime="00:04:57.51" resultid="3260" heatid="10291" lane="7" entrytime="00:05:05.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="200" swimtime="00:02:26.57" />
                    <SPLIT distance="300" swimtime="00:03:42.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-16" firstname="MARCIN" gender="M" lastname="HORBACZ" nation="POL" athleteid="3261">
              <RESULTS>
                <RESULT eventid="1109" points="683" swimtime="00:02:22.38" resultid="3262" heatid="10122" lane="2" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="707" swimtime="00:00:57.71" resultid="3263" heatid="10157" lane="4" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1465" points="805" swimtime="00:02:04.85" resultid="3264" heatid="10223" lane="4" entrytime="00:02:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="607" swimtime="00:00:27.33" resultid="3265" heatid="10256" lane="3" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1686" points="754" swimtime="00:04:29.56" resultid="3266" heatid="10292" lane="4" entrytime="00:04:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="200" swimtime="00:02:14.61" />
                    <SPLIT distance="300" swimtime="00:03:22.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" name="UKS Victoria Józefów" nation="POL" region="MAZ" shortname="Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="KOWALCZYK ALICJA" />
          <ATHLETES>
            <ATHLETE birthdate="1980-11-08" firstname="Alicja" gender="F" lastname="Kowalczyk-Kędzierska" nation="POL" athleteid="3268">
              <RESULTS>
                <RESULT eventid="1061" points="629" swimtime="00:00:33.65" resultid="3269" heatid="10099" lane="8" entrytime="00:00:35.80" />
                <RESULT eventid="1178" points="503" swimtime="00:00:38.32" resultid="3270" heatid="10129" lane="3" entrytime="00:00:38.20" />
                <RESULT eventid="1352" points="442" swimtime="00:00:43.67" resultid="3271" heatid="10181" lane="8" entrytime="00:00:44.34" />
                <RESULT eventid="1385" points="477" reactiontime="+90" swimtime="00:01:23.88" resultid="3272" heatid="10196" lane="5" entrytime="00:01:22.20" />
                <RESULT eventid="1525" points="389" swimtime="00:01:27.57" resultid="3273" heatid="10233" lane="7" entrytime="00:01:28.90" />
                <RESULT eventid="1590" points="398" reactiontime="+96" swimtime="00:03:08.98" resultid="3274" heatid="10260" lane="1" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORMAS" name="Orka Masters" nation="POL">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK MARIAN" phone="530556313" />
          <ATHLETES>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="OTLIK" nation="POL" athleteid="3554">
              <RESULTS>
                <RESULT eventid="1077" points="422" swimtime="00:00:36.50" resultid="3555" heatid="10104" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1109" points="411" swimtime="00:03:07.94" resultid="3556" heatid="10117" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="494" swimtime="00:01:09.28" resultid="3557" heatid="10151" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1324" points="332" swimtime="00:03:42.18" resultid="3558" heatid="10173" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="289" swimtime="00:00:46.46" resultid="3559" heatid="10188" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1465" points="388" swimtime="00:02:48.01" resultid="3560" heatid="10218" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="272" swimtime="00:01:34.60" resultid="3561" heatid="10237" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1574" points="474" status="EXH" swimtime="00:00:31.45" resultid="3562" heatid="10252" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1686" points="345" swimtime="00:06:14.32" resultid="3563" heatid="10288" lane="3" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="200" swimtime="00:03:01.75" />
                    <SPLIT distance="300" swimtime="00:04:40.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="CIECIOR" nation="POL" athleteid="3564">
              <RESULTS>
                <RESULT eventid="1077" points="587" swimtime="00:00:36.26" resultid="3565" heatid="10104" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1109" points="517" swimtime="00:03:20.67" resultid="3566" heatid="10117" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="427" swimtime="00:00:44.39" resultid="3567" heatid="10136" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1228" points="519" swimtime="00:01:17.58" resultid="3568" heatid="10150" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="1401" points="461" reactiontime="+90" swimtime="00:01:35.24" resultid="3569" heatid="10201" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1497" points="487" swimtime="00:07:22.47" resultid="3570" heatid="10228" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                    <SPLIT distance="200" swimtime="00:03:36.34" />
                    <SPLIT distance="300" swimtime="00:05:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="394" swimtime="00:01:35.52" resultid="3571" heatid="10236" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="1686" points="445" swimtime="00:06:26.49" resultid="3572" heatid="10288" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="200" swimtime="00:03:07.28" />
                    <SPLIT distance="300" swimtime="00:04:48.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-08-10" firstname="Jan" gender="M" lastname="KLAPSIA" nation="POL" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1195" points="154" swimtime="00:01:11.21" resultid="3574" heatid="10131" lane="5" />
                <RESULT eventid="1228" points="59" swimtime="00:02:52.02" resultid="3575" heatid="10147" lane="1" />
                <RESULT eventid="1369" points="140" swimtime="00:01:13.56" resultid="3576" heatid="10183" lane="4" />
                <RESULT eventid="1401" points="124" reactiontime="+120" swimtime="00:02:49.16" resultid="3577" heatid="10198" lane="2" />
                <RESULT eventid="1574" points="67" swimtime="00:01:13.96" resultid="3578" heatid="10246" lane="3" />
                <RESULT eventid="1654" points="115" swimtime="00:02:59.68" resultid="3579" heatid="10274" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="IRCZYK" nation="POL" athleteid="3580">
              <RESULTS>
                <RESULT eventid="1109" points="256" swimtime="00:04:13.71" resultid="3581" heatid="10115" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="255" swimtime="00:32:06.43" resultid="3582" heatid="10300" lane="6" entrytime="00:29:00.00" />
                <RESULT eventid="1292" points="152" swimtime="00:05:03.28" resultid="3583" heatid="10163" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="441" swimtime="00:03:51.93" resultid="3584" heatid="10172" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="238" swimtime="00:03:47.84" resultid="3585" heatid="10216" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="272" swimtime="00:08:57.18" resultid="3586" heatid="10227" lane="3" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.64" />
                    <SPLIT distance="200" swimtime="00:04:55.14" />
                    <SPLIT distance="300" swimtime="00:06:55.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="152" swimtime="00:02:11.03" resultid="3587" heatid="10235" lane="6" entrytime="00:02:00.00" />
                <RESULT eventid="1686" points="218" swimtime="00:08:09.91" resultid="3588" heatid="10286" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.63" />
                    <SPLIT distance="200" swimtime="00:03:59.03" />
                    <SPLIT distance="300" swimtime="00:06:06.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WAMAS" name="Warsaw Masters Team" nation="POL" shortname="Warsaw Masters">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 4444" />
          <ATHLETES>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="3590">
              <RESULTS>
                <RESULT eventid="1109" points="936" swimtime="00:02:31.86" resultid="6666" heatid="10120" lane="4" entrytime="00:02:37.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="891" swimtime="00:00:59.10" resultid="6667" heatid="10158" lane="1" entrytime="00:00:58.59" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1465" points="841" swimtime="00:02:11.67" resultid="6668" heatid="10223" lane="1" entrytime="00:02:13.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="747" swimtime="00:00:27.96" resultid="6669" heatid="10256" lane="2" entrytime="00:00:27.31" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1686" points="750" swimtime="00:04:55.34" resultid="6670" heatid="10291" lane="4" entrytime="00:04:57.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="200" swimtime="00:02:29.82" />
                    <SPLIT distance="300" swimtime="00:03:44.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="Michalczyk" nation="POL" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1212" points="445" swimtime="00:01:15.23" resultid="6671" heatid="10144" lane="4" entrytime="00:01:13.80" entrycourse="LCM" />
                <RESULT eventid="1308" points="428" swimtime="00:03:29.36" resultid="6672" heatid="10168" lane="4" entrytime="00:03:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="413" swimtime="00:00:45.77" resultid="6673" heatid="10181" lane="2" entrytime="00:00:43.90" />
                <RESULT eventid="1449" points="409" swimtime="00:02:45.54" resultid="6674" heatid="10212" lane="3" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="438" swimtime="00:01:23.15" resultid="6675" heatid="10233" lane="5" entrytime="00:01:20.60" entrycourse="LCM" />
                <RESULT eventid="1638" points="393" swimtime="00:01:36.53" resultid="6676" heatid="10272" lane="4" entrytime="00:01:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1162" points="347" swimtime="00:23:19.39" resultid="6677" heatid="10298" lane="4" entrytime="00:22:30.00" />
                <RESULT eventid="1195" points="275" swimtime="00:00:40.11" resultid="6678" heatid="10137" lane="5" entrytime="00:00:37.89" entrycourse="LCM" />
                <RESULT eventid="1228" points="390" swimtime="00:01:09.31" resultid="6679" heatid="10153" lane="8" entrytime="00:01:07.57" entrycourse="LCM" />
                <RESULT eventid="1401" points="247" reactiontime="+90" swimtime="00:01:30.30" resultid="6680" heatid="10202" lane="2" entrytime="00:01:24.32" entrycourse="LCM" />
                <RESULT eventid="1465" points="335" swimtime="00:02:40.73" resultid="6681" heatid="10220" lane="8" entrytime="00:02:34.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="403" swimtime="00:00:31.21" resultid="6682" heatid="10252" lane="8" entrytime="00:00:30.51" entrycourse="LCM" />
                <RESULT eventid="1686" points="346" swimtime="00:05:42.63" resultid="6683" heatid="10290" lane="7" entrytime="00:05:36.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="200" swimtime="00:02:47.57" />
                    <SPLIT distance="300" swimtime="00:04:16.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan" gender="M" lastname="Boboli" nation="POL" athleteid="3611">
              <RESULTS>
                <RESULT eventid="1077" points="515" swimtime="00:00:39.72" resultid="6684" heatid="10104" lane="8" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1195" points="198" swimtime="00:01:00.53" resultid="6685" heatid="10133" lane="6" entrytime="00:00:56.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="362" swimtime="00:01:32.65" resultid="6686" heatid="10148" lane="3" entrytime="00:01:26.00" entrycourse="LCM" />
                <RESULT eventid="1369" points="46" swimtime="00:01:40.87" resultid="6687" heatid="10184" lane="1" entrytime="00:00:58.00" entrycourse="LCM" />
                <RESULT eventid="1574" points="455" swimtime="00:00:36.73" resultid="6688" heatid="10248" lane="5" entrytime="00:00:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="3617">
              <RESULTS>
                <RESULT eventid="1109" points="231" swimtime="00:03:47.62" resultid="6689" heatid="10114" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="271" swimtime="00:01:24.56" resultid="6690" heatid="10148" lane="2" entrytime="00:01:29.01" entrycourse="LCM" />
                <RESULT eventid="1324" points="363" swimtime="00:03:35.82" resultid="6691" heatid="10173" lane="1" entrytime="00:03:37.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="310" swimtime="00:00:45.37" resultid="6692" heatid="10186" lane="3" entrytime="00:00:44.96" entrycourse="LCM" />
                <RESULT eventid="1574" points="256" swimtime="00:00:38.59" resultid="6693" heatid="10247" lane="3" entrytime="00:00:38.52" entrycourse="LCM" />
                <RESULT eventid="1654" points="344" swimtime="00:01:38.06" resultid="6694" heatid="10276" lane="4" entrytime="00:01:39.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="3624">
              <RESULTS>
                <RESULT eventid="1077" points="686" swimtime="00:00:31.05" resultid="6695" heatid="10108" lane="4" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1109" points="678" swimtime="00:02:39.17" resultid="6696" heatid="10121" lane="3" entrytime="00:02:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="693" swimtime="00:00:32.60" resultid="6697" heatid="10139" lane="5" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="681" swimtime="00:01:02.25" resultid="6698" heatid="10157" lane="7" entrytime="00:00:59.59" entrycourse="LCM" />
                <RESULT eventid="1401" points="788" reactiontime="+81" swimtime="00:01:10.43" resultid="6699" heatid="10205" lane="6" entrytime="00:01:07.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="440" swimtime="00:02:41.07" resultid="6700" heatid="10222" lane="7" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="612" swimtime="00:00:28.89" resultid="6701" heatid="10254" lane="4" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1606" points="684" reactiontime="+94" swimtime="00:02:39.88" resultid="6702" heatid="10266" lane="8" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-06" firstname="Paweł" gender="M" lastname="Gajewski" nation="POL" athleteid="3633">
              <RESULTS>
                <RESULT eventid="1162" points="163" swimtime="00:29:56.84" resultid="6703" heatid="10301" lane="4" entrytime="00:30:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Stanisławska" nation="POL" athleteid="3635">
              <RESULTS>
                <RESULT eventid="1061" points="310" swimtime="00:00:43.03" resultid="6704" heatid="10097" lane="6" entrytime="00:00:45.00" entrycourse="LCM" />
                <RESULT eventid="1141" points="288" swimtime="00:14:00.64" resultid="6705" heatid="10294" lane="3" entrytime="00:14:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                    <SPLIT distance="200" swimtime="00:03:19.86" />
                    <SPLIT distance="300" swimtime="00:05:07.70" />
                    <SPLIT distance="400" swimtime="00:06:55.92" />
                    <SPLIT distance="500" swimtime="00:08:44.95" />
                    <SPLIT distance="600" swimtime="00:10:33.92" />
                    <SPLIT distance="700" swimtime="00:12:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="293" swimtime="00:01:26.47" resultid="6706" heatid="10142" lane="2" entrytime="00:01:30.00" entrycourse="LCM" />
                <RESULT eventid="1276" status="DSQ" swimtime="00:03:53.99" resultid="6707" heatid="10162" lane="4" entrytime="00:04:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="258" swimtime="00:03:12.87" resultid="6708" heatid="10211" lane="2" entrytime="00:03:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="275" swimtime="00:07:46.05" resultid="6709" heatid="10224" lane="5" entrytime="00:08:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.78" />
                    <SPLIT distance="200" swimtime="00:03:53.00" />
                    <SPLIT distance="300" swimtime="00:06:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="176" swimtime="00:01:52.56" resultid="6710" heatid="10232" lane="6" entrytime="00:01:50.00" entrycourse="LCM" />
                <RESULT eventid="1670" points="266" swimtime="00:06:53.22" resultid="6711" heatid="10283" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.74" />
                    <SPLIT distance="200" swimtime="00:03:23.10" />
                    <SPLIT distance="300" swimtime="00:05:11.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="3644">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1109" points="912" swimtime="00:02:46.11" resultid="6712" heatid="10120" lane="1" entrytime="00:02:46.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1228" points="913" swimtime="00:01:04.29" resultid="6713" heatid="10153" lane="3" entrytime="00:01:05.80" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1401" points="855" reactiontime="+83" swimtime="00:01:17.53" resultid="6714" heatid="10203" lane="7" entrytime="00:01:16.80" entrycourse="LCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1465" points="955" swimtime="00:02:23.35" resultid="6715" heatid="10221" lane="6" entrytime="00:02:23.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="898" reactiontime="+77" swimtime="00:02:47.79" resultid="6716" heatid="10265" lane="2" entrytime="00:02:46.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-18" firstname="Robert" gender="M" lastname="Nowicki" nation="POL" athleteid="3650">
              <RESULTS>
                <RESULT eventid="1162" points="239" swimtime="00:29:23.49" resultid="6717" heatid="10300" lane="1" entrytime="00:29:30.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="223" swimtime="00:01:33.76" resultid="6718" heatid="10148" lane="7" entrytime="00:01:35.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="206" swimtime="00:03:30.27" resultid="6719" heatid="10215" lane="4" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" status="DNS" swimtime="00:00:00.00" resultid="6720" heatid="10286" lane="5" entrytime="00:07:20.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="3655">
              <RESULTS>
                <RESULT eventid="1212" points="331" swimtime="00:01:23.44" resultid="6721" heatid="10142" lane="6" entrytime="00:01:27.75" entrycourse="LCM" />
                <RESULT eventid="1385" points="331" reactiontime="+102" swimtime="00:01:33.51" resultid="6722" heatid="10195" lane="6" entrytime="00:01:35.89" entrycourse="LCM" />
                <RESULT eventid="1449" points="314" swimtime="00:03:05.00" resultid="6723" heatid="10211" lane="1" entrytime="00:03:10.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="315" reactiontime="+99" swimtime="00:03:23.46" resultid="6724" heatid="10259" lane="2" entrytime="00:03:29.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="3660">
              <RESULTS>
                <RESULT eventid="1077" points="195" swimtime="00:01:02.06" resultid="6725" heatid="10100" lane="5" entrytime="00:02:30.00" entrycourse="LCM" />
                <RESULT eventid="1109" points="312" swimtime="00:04:39.96" resultid="6726" heatid="10115" lane="1" entrytime="00:04:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="259" swimtime="00:01:01.96" resultid="6727" heatid="10133" lane="7" entrytime="00:00:58.00" entrycourse="LCM" />
                <RESULT eventid="1324" points="419" swimtime="00:04:29.15" resultid="6728" heatid="10170" lane="4" entrytime="00:04:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:08.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="424" swimtime="00:00:53.35" resultid="6729" heatid="10184" lane="7" entrytime="00:00:55.00" entrycourse="LCM" />
                <RESULT eventid="1401" points="173" reactiontime="+92" swimtime="00:02:37.84" resultid="6730" heatid="10198" lane="3" entrytime="00:02:30.00" entrycourse="LCM" />
                <RESULT eventid="1542" points="188" swimtime="00:02:40.47" resultid="6731" heatid="10235" lane="1" entrytime="00:02:35.00" entrycourse="LCM" />
                <RESULT eventid="1654" points="298" swimtime="00:02:12.56" resultid="6732" heatid="10274" lane="4" entrytime="00:02:15.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="3672">
              <RESULTS>
                <RESULT eventid="1061" points="387" swimtime="00:00:39.57" resultid="6733" heatid="10097" lane="7" entrytime="00:00:45.04" entrycourse="LCM" />
                <RESULT eventid="1212" points="343" swimtime="00:01:22.90" resultid="6734" heatid="10142" lane="5" entrytime="00:01:26.30" entrycourse="LCM" />
                <RESULT eventid="1449" points="301" swimtime="00:03:06.81" resultid="6735" heatid="10211" lane="5" entrytime="00:03:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="368" swimtime="00:00:37.07" resultid="6736" heatid="10242" lane="4" entrytime="00:00:37.88" entrycourse="LCM" />
                <RESULT eventid="1670" points="316" swimtime="00:06:33.27" resultid="6737" heatid="10283" lane="5" entrytime="00:06:44.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.08" />
                    <SPLIT distance="200" swimtime="00:03:17.44" />
                    <SPLIT distance="300" swimtime="00:04:58.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-06-16" firstname="Elżbieta" gender="F" lastname="Janik" nation="POL" athleteid="3678">
              <RESULTS>
                <RESULT eventid="1178" points="323" swimtime="00:01:09.82" resultid="6738" heatid="10126" lane="5" entrytime="00:01:07.30" entrycourse="LCM" />
                <RESULT eventid="1385" points="368" reactiontime="+71" swimtime="00:02:29.60" resultid="6739" heatid="10193" lane="4" entrytime="00:02:23.61" entrycourse="LCM" />
                <RESULT eventid="1590" points="381" reactiontime="+82" swimtime="00:05:21.75" resultid="6740" heatid="10258" lane="7" entrytime="00:04:59.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:39.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-14" firstname="Sebastian" gender="M" lastname="Wojciechowski" nation="POL" athleteid="3682">
              <RESULTS>
                <RESULT eventid="1162" points="273" swimtime="00:26:13.28" resultid="6741" heatid="10300" lane="5" entrytime="00:28:23.00" entrycourse="LCM" />
                <RESULT eventid="1465" points="268" swimtime="00:03:03.51" resultid="6742" heatid="10216" lane="5" entrytime="00:03:01.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="252" swimtime="00:06:37.34" resultid="6743" heatid="10287" lane="6" entrytime="00:06:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.48" />
                    <SPLIT distance="200" swimtime="00:03:15.51" />
                    <SPLIT distance="300" swimtime="00:05:00.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="3686">
              <RESULTS>
                <RESULT eventid="1093" points="645" swimtime="00:03:04.10" resultid="6744" heatid="10112" lane="3" entrytime="00:03:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="687" swimtime="00:03:13.98" resultid="6745" heatid="10169" lane="2" entrytime="00:03:12.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1352" points="747" swimtime="00:00:39.76" resultid="6746" heatid="10182" lane="7" entrytime="00:00:40.70" entrycourse="LCM" />
                <RESULT eventid="1449" points="491" swimtime="00:02:54.88" resultid="6747" heatid="10212" lane="6" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="674" swimtime="00:01:30.39" resultid="6748" heatid="10273" lane="7" entrytime="00:01:28.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="3692">
              <RESULTS>
                <RESULT eventid="1324" points="527" swimtime="00:02:55.74" resultid="6749" heatid="10177" lane="5" entrytime="00:02:40.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="744" swimtime="00:00:31.21" resultid="6750" heatid="10192" lane="5" entrytime="00:00:31.23" entrycourse="LCM" />
                <RESULT eventid="1654" points="607" swimtime="00:01:14.62" resultid="6751" heatid="10281" lane="4" entrytime="00:01:10.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-07-11" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="3696">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="6752" heatid="10105" lane="1" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="6753" heatid="10136" lane="1" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="6754" heatid="10151" lane="8" entrytime="00:01:13.14" entrycourse="SCM" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="6755" heatid="10190" lane="4" entrytime="00:00:35.94" entrycourse="LCM" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="6756" heatid="10252" lane="1" entrytime="00:00:30.31" entrycourse="LCM" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="6757" heatid="10279" lane="1" entrytime="00:01:25.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="3703">
              <RESULTS>
                <RESULT eventid="1228" status="DSQ" swimtime="00:01:00.26" resultid="6758" heatid="10157" lane="6" entrytime="00:00:59.24" entrycourse="LCM" />
                <RESULT eventid="1401" points="439" reactiontime="+89" swimtime="00:01:13.96" resultid="6759" heatid="10204" lane="3" entrytime="00:01:09.99" entrycourse="LCM" />
                <RESULT eventid="1574" points="632" swimtime="00:00:26.49" resultid="6760" heatid="10257" lane="8" entrytime="00:00:26.75" entrycourse="LCM" />
                <RESULT eventid="1686" points="436" swimtime="00:05:18.33" resultid="6761" heatid="10291" lane="3" entrytime="00:04:59.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="200" swimtime="00:02:37.37" />
                    <SPLIT distance="300" swimtime="00:04:00.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="3708">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="6762" heatid="10120" lane="5" entrytime="00:02:39.89" entrycourse="LCM" />
                <RESULT eventid="1162" status="DNS" swimtime="00:00:00.00" resultid="6763" heatid="10297" lane="7" entrytime="00:22:08.15" entrycourse="LCM" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="6764" heatid="10138" lane="1" entrytime="00:00:36.12" entrycourse="LCM" />
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="6765" heatid="10165" lane="4" entrytime="00:02:47.19" entrycourse="LCM" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="6766" heatid="10189" lane="4" entrytime="00:00:37.10" entrycourse="LCM" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="6767" heatid="10230" lane="5" entrytime="00:05:50.19" entrycourse="LCM" />
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="6768" heatid="10239" lane="1" entrytime="00:01:14.19" entrycourse="LCM" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="6769" heatid="10280" lane="8" entrytime="00:01:21.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+83" swimtime="00:02:18.12" resultid="6772" heatid="10161" lane="6" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3624" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3692" number="2" />
                    <RELAYPOSITION athleteid="3611" number="3" />
                    <RELAYPOSITION athleteid="3703" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1433" swimtime="00:01:55.86" resultid="6774" heatid="10208" lane="5" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3624" number="1" />
                    <RELAYPOSITION athleteid="3603" number="2" />
                    <RELAYPOSITION athleteid="3692" number="3" />
                    <RELAYPOSITION athleteid="3703" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1244" reactiontime="+90" swimtime="00:02:50.71" resultid="6771" heatid="10159" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3655" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="3672" number="2" />
                    <RELAYPOSITION athleteid="3596" number="3" />
                    <RELAYPOSITION athleteid="3635" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1417" swimtime="00:02:31.27" resultid="6773" heatid="10206" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3635" number="1" />
                    <RELAYPOSITION athleteid="3672" number="2" />
                    <RELAYPOSITION athleteid="3655" number="3" />
                    <RELAYPOSITION athleteid="3596" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:20.44" resultid="6770" heatid="10124" lane="3" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3635" number="1" />
                    <RELAYPOSITION athleteid="3672" number="2" />
                    <RELAYPOSITION athleteid="3611" number="3" />
                    <RELAYPOSITION athleteid="3624" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+91" swimtime="00:02:29.59" resultid="6775" heatid="10269" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3624" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="3672" number="2" />
                    <RELAYPOSITION athleteid="3703" number="3" />
                    <RELAYPOSITION athleteid="3635" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" name="MOTYL SENIOR MOSiR Stalowa Wola" nation="POL" region="PDK" shortname="SENIOR Stalowa Wola">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="15-8422562 wew.45" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="3737">
              <RESULTS>
                <RESULT eventid="1109" points="545" swimtime="00:02:33.49" resultid="3738" heatid="10120" lane="2" entrytime="00:02:43.03">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="691" swimtime="00:00:31.07" resultid="3739" heatid="10140" lane="7" entrytime="00:00:31.18" />
                <RESULT eventid="1228" points="619" swimtime="00:01:00.33" resultid="3740" heatid="10156" lane="4" entrytime="00:01:00.66" />
                <RESULT eventid="1401" points="640" reactiontime="+86" swimtime="00:01:08.24" resultid="3741" heatid="10204" lane="5" entrytime="00:01:09.53" />
                <RESULT eventid="1574" points="654" swimtime="00:00:26.67" resultid="3742" heatid="10256" lane="7" entrytime="00:00:27.36" />
                <RESULT eventid="1606" points="583" reactiontime="+84" swimtime="00:02:32.22" resultid="3743" heatid="10265" lane="5" entrytime="00:02:36.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="3744">
              <RESULTS>
                <RESULT eventid="1077" points="834" swimtime="00:00:28.32" resultid="3745" heatid="10110" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="1109" points="846" swimtime="00:02:24.15" resultid="3746" heatid="10122" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="752" swimtime="00:02:23.39" resultid="3747" heatid="10166" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="601" swimtime="00:00:34.94" resultid="3748" heatid="10192" lane="1" entrytime="00:00:33.80" />
                <RESULT eventid="1497" points="780" swimtime="00:05:18.67" resultid="3749" heatid="10231" lane="3" entrytime="00:05:10.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="200" swimtime="00:02:32.61" />
                    <SPLIT distance="300" swimtime="00:04:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="880" swimtime="00:01:01.22" resultid="3750" heatid="10240" lane="5" entrytime="00:01:00.85" />
                <RESULT eventid="1654" points="721" swimtime="00:01:14.92" resultid="3751" heatid="10281" lane="2" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="3752">
              <RESULTS>
                <RESULT eventid="1109" points="471" swimtime="00:03:27.00" resultid="3753" heatid="10117" lane="8" entrytime="00:03:36.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="533" swimtime="00:00:41.24" resultid="3754" heatid="10135" lane="6" entrytime="00:00:44.07" />
                <RESULT eventid="1324" points="472" swimtime="00:03:46.62" resultid="3755" heatid="10172" lane="4" entrytime="00:03:39.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="485" reactiontime="+92" swimtime="00:01:33.67" resultid="3756" heatid="10201" lane="8" entrytime="00:01:33.65" />
                <RESULT eventid="1497" points="471" swimtime="00:07:27.29" resultid="3757" heatid="10228" lane="6" entrytime="00:07:26.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.92" />
                    <SPLIT distance="200" swimtime="00:03:48.82" />
                    <SPLIT distance="300" swimtime="00:05:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="485" reactiontime="+96" swimtime="00:03:26.08" resultid="3758" heatid="10263" lane="1" entrytime="00:03:39.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="422" swimtime="00:06:33.28" resultid="3759" heatid="10287" lane="4" entrytime="00:06:20.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="200" swimtime="00:03:14.47" />
                    <SPLIT distance="300" swimtime="00:04:58.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="Kalbarczyk" nation="POL" athleteid="3760">
              <RESULTS>
                <RESULT eventid="1077" points="494" swimtime="00:00:33.72" resultid="3761" heatid="10105" lane="4" entrytime="00:00:34.15" />
                <RESULT eventid="1109" points="497" swimtime="00:02:52.12" resultid="3762" heatid="10119" lane="3" entrytime="00:02:54.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="465" swimtime="00:01:08.95" resultid="3763" heatid="10151" lane="3" entrytime="00:01:10.71" />
                <RESULT eventid="1324" points="410" swimtime="00:03:22.25" resultid="3764" heatid="10173" lane="4" entrytime="00:03:25.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="434" swimtime="00:02:36.33" resultid="3765" heatid="10218" lane="3" entrytime="00:02:42.15">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="442" swimtime="00:06:24.90" resultid="3766" heatid="10229" lane="2" entrytime="00:06:35.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.02" />
                    <SPLIT distance="200" swimtime="00:03:10.52" />
                    <SPLIT distance="300" swimtime="00:05:00.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="469" reactiontime="+87" swimtime="00:02:54.37" resultid="3767" heatid="10264" lane="3" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="400" swimtime="00:05:40.71" resultid="3768" heatid="10290" lane="1" entrytime="00:05:37.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                    <SPLIT distance="200" swimtime="00:02:44.75" />
                    <SPLIT distance="300" swimtime="00:04:14.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="3769">
              <RESULTS>
                <RESULT eventid="1109" points="629" swimtime="00:02:53.32" resultid="3770" heatid="10119" lane="2" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="582" swimtime="00:01:08.13" resultid="3771" heatid="10152" lane="6" entrytime="00:01:09.54" />
                <RESULT eventid="1292" points="416" swimtime="00:03:21.12" resultid="3772" heatid="10164" lane="3" entrytime="00:03:25.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="494" swimtime="00:02:37.25" resultid="3773" heatid="10219" lane="8" entrytime="00:02:38.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="583" swimtime="00:06:18.53" resultid="3774" heatid="10229" lane="4" entrytime="00:06:24.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="200" swimtime="00:03:05.05" />
                    <SPLIT distance="300" swimtime="00:04:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="570" reactiontime="+90" swimtime="00:02:59.59" resultid="3775" heatid="10264" lane="1" entrytime="00:03:03.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="450" swimtime="00:05:50.16" resultid="3776" heatid="10289" lane="6" entrytime="00:05:48.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="200" swimtime="00:02:50.43" />
                    <SPLIT distance="300" swimtime="00:04:22.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-29" firstname="Jarosław" gender="M" lastname="Niedbałowski" nation="POL" athleteid="3777">
              <RESULTS>
                <RESULT eventid="1077" points="437" swimtime="00:00:36.98" resultid="3778" heatid="10103" lane="5" entrytime="00:00:38.25" />
                <RESULT eventid="1324" points="548" swimtime="00:03:21.22" resultid="3779" heatid="10174" lane="6" entrytime="00:03:16.41">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="593" swimtime="00:00:39.51" resultid="3780" heatid="10189" lane="3" entrytime="00:00:37.42" />
                <RESULT eventid="1574" points="571" swimtime="00:00:31.47" resultid="3781" heatid="10251" lane="8" entrytime="00:00:31.59" />
                <RESULT eventid="1654" points="580" swimtime="00:01:29.05" resultid="3782" heatid="10278" lane="5" entrytime="00:01:27.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="3783">
              <RESULTS>
                <RESULT eventid="1061" points="477" swimtime="00:00:39.03" resultid="3784" heatid="10098" lane="2" entrytime="00:00:39.11" />
                <RESULT eventid="1093" points="495" swimtime="00:03:21.12" resultid="3785" heatid="10112" lane="1" entrytime="00:03:13.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DSQ" swimtime="00:01:19.74" resultid="3786" heatid="10144" lane="8" entrytime="00:01:18.11" />
                <RESULT eventid="1308" points="515" swimtime="00:03:33.52" resultid="3787" heatid="10168" lane="7" entrytime="00:03:32.33">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="488" swimtime="00:00:45.81" resultid="3788" heatid="10180" lane="5" entrytime="00:00:46.11" />
                <RESULT eventid="1481" points="559" swimtime="00:06:57.00" resultid="3789" heatid="10225" lane="6" entrytime="00:06:57.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.12" />
                    <SPLIT distance="200" swimtime="00:03:32.25" />
                    <SPLIT distance="300" swimtime="00:05:24.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="424" swimtime="00:01:33.62" resultid="3790" heatid="10233" lane="1" entrytime="00:01:32.21" />
                <RESULT eventid="1638" points="458" swimtime="00:01:42.81" resultid="3791" heatid="10272" lane="7" entrytime="00:01:40.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="3792">
              <RESULTS>
                <RESULT eventid="1077" points="701" swimtime="00:00:30.82" resultid="3793" heatid="10107" lane="8" entrytime="00:00:32.40" />
                <RESULT eventid="1228" points="609" swimtime="00:01:04.60" resultid="3794" heatid="10151" lane="2" entrytime="00:01:12.67" />
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="3795" heatid="10164" lane="5" entrytime="00:03:20.12" />
                <RESULT eventid="1401" points="519" reactiontime="+74" swimtime="00:01:20.97" resultid="3796" heatid="10202" lane="4" entrytime="00:01:19.83" />
                <RESULT eventid="1465" points="439" swimtime="00:02:41.20" resultid="3797" heatid="10219" lane="6" entrytime="00:02:35.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="680" swimtime="00:00:27.89" resultid="3798" heatid="10249" lane="7" entrytime="00:00:34.07" />
                <RESULT eventid="1606" points="439" reactiontime="+82" swimtime="00:03:05.33" resultid="3799" heatid="10264" lane="6" entrytime="00:02:59.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="3800">
              <RESULTS>
                <RESULT eventid="1109" points="549" swimtime="00:02:33.13" resultid="3801" heatid="10121" lane="7" entrytime="00:02:35.39">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="572" swimtime="00:02:50.78" resultid="3802" heatid="10176" lane="4" entrytime="00:02:50.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="586" swimtime="00:00:34.42" resultid="3803" heatid="10191" lane="3" entrytime="00:00:34.30" />
                <RESULT eventid="1497" points="583" swimtime="00:05:41.57" resultid="3804" heatid="10230" lane="7" entrytime="00:06:00.19">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="200" swimtime="00:02:51.87" />
                    <SPLIT distance="300" swimtime="00:04:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="594" swimtime="00:01:15.26" resultid="3805" heatid="10281" lane="8" entrytime="00:01:17.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-04" firstname="Paweł" gender="M" lastname="Opaliński" nation="POL" athleteid="3806">
              <RESULTS>
                <RESULT eventid="1077" points="547" swimtime="00:00:30.73" resultid="3807" heatid="10107" lane="5" entrytime="00:00:31.12" />
                <RESULT eventid="1228" points="574" swimtime="00:01:01.85" resultid="3808" heatid="10156" lane="7" entrytime="00:01:01.59" />
                <RESULT eventid="1324" points="571" swimtime="00:02:50.92" resultid="3809" heatid="10176" lane="5" entrytime="00:02:57.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="612" swimtime="00:00:33.93" resultid="3810" heatid="10191" lane="8" entrytime="00:00:35.01" />
                <RESULT eventid="1465" points="602" swimtime="00:02:17.52" resultid="3811" heatid="10222" lane="2" entrytime="00:02:19.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="530" swimtime="00:01:18.17" resultid="3812" heatid="10280" lane="6" entrytime="00:01:18.36" />
                <RESULT eventid="1686" status="DNS" swimtime="00:00:00.00" resultid="3813" heatid="10290" lane="4" entrytime="00:05:19.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="3814">
              <RESULTS>
                <RESULT eventid="1195" points="489" swimtime="00:00:34.87" resultid="3815" heatid="10138" lane="3" entrytime="00:00:35.36" />
                <RESULT eventid="1324" status="DSQ" swimtime="00:03:10.76" resultid="3816" heatid="10175" lane="2" entrytime="00:03:12.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="469" swimtime="00:00:37.08" resultid="3817" heatid="10189" lane="6" entrytime="00:00:37.60" />
                <RESULT eventid="1497" points="374" swimtime="00:06:36.00" resultid="3818" heatid="10229" lane="7" entrytime="00:06:36.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="200" swimtime="00:03:20.13" />
                    <SPLIT distance="300" swimtime="00:05:06.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+80" swimtime="00:02:02.12" resultid="3819" heatid="10161" lane="5" entrytime="00:02:02.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3737" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3800" number="2" />
                    <RELAYPOSITION athleteid="3744" number="3" />
                    <RELAYPOSITION athleteid="3792" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+84" swimtime="00:02:22.92" resultid="3820" heatid="10160" lane="4" entrytime="00:02:22.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3760" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3777" number="2" />
                    <RELAYPOSITION athleteid="3806" number="3" />
                    <RELAYPOSITION athleteid="3752" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1433" swimtime="00:01:52.70" resultid="3821" heatid="10208" lane="3" entrytime="00:01:52.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3737" number="1" />
                    <RELAYPOSITION athleteid="3800" number="2" />
                    <RELAYPOSITION athleteid="3792" number="3" />
                    <RELAYPOSITION athleteid="3744" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1433" swimtime="00:02:04.76" resultid="3822" heatid="10208" lane="8" entrytime="00:02:02.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3760" number="1" />
                    <RELAYPOSITION athleteid="3777" number="2" />
                    <RELAYPOSITION athleteid="3752" number="3" />
                    <RELAYPOSITION athleteid="3806" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" name="K.S. niezrzeszeni.pl" nation="POL" region="WA" shortname="niezrzeszeni.pl">
          <CONTACT city="Warszawa" email="niezrzeszenipl@gmail.com" internet="niezrzeszeni.pl" name="Wawer Matylda Katarzyna" phone="505960036" />
          <ATHLETES>
            <ATHLETE birthdate="1960-07-16" firstname="Matylda Katarzyna" gender="F" lastname="Wawer" nation="POL" athleteid="3839">
              <RESULTS>
                <RESULT eventid="1061" points="435" swimtime="00:00:43.52" resultid="3840" heatid="10095" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="412" swimtime="00:01:27.39" resultid="3841" heatid="10142" lane="4" entrytime="00:01:26.00" />
                <RESULT eventid="1449" points="317" swimtime="00:03:30.06" resultid="3842" heatid="10210" lane="4" entrytime="00:03:24.93">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="505" swimtime="00:00:36.59" resultid="3843" heatid="10243" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1670" points="307" swimtime="00:07:38.06" resultid="3844" heatid="10282" lane="4" entrytime="00:07:46.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="200" swimtime="00:03:39.97" />
                    <SPLIT distance="300" swimtime="00:05:40.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-16" firstname="Paweł" gender="M" lastname="Borkowski" nation="POL" athleteid="3845">
              <RESULTS>
                <RESULT eventid="1228" points="445" swimtime="00:01:04.64" resultid="3846" heatid="10155" lane="4" entrytime="00:01:02.01" />
                <RESULT eventid="1465" points="372" swimtime="00:02:29.66" resultid="3847" heatid="10221" lane="3" entrytime="00:02:22.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="490" swimtime="00:00:28.30" resultid="3848" heatid="10256" lane="8" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="3849">
              <RESULTS>
                <RESULT eventid="1162" points="373" swimtime="00:27:15.89" resultid="3850" heatid="10299" lane="6" entrytime="00:25:30.00" />
                <RESULT eventid="1228" points="319" swimtime="00:01:25.86" resultid="3851" heatid="10149" lane="7" entrytime="00:01:23.00" />
                <RESULT eventid="1324" points="355" swimtime="00:03:52.65" resultid="3852" heatid="10172" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="377" swimtime="00:00:45.94" resultid="3853" heatid="10186" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1497" points="291" swimtime="00:08:29.94" resultid="3854" heatid="10227" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.52" />
                    <SPLIT distance="200" swimtime="00:04:38.63" />
                    <SPLIT distance="300" swimtime="00:06:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="156" swimtime="00:01:59.57" resultid="3855" heatid="10234" lane="4" />
                <RESULT eventid="1686" points="373" swimtime="00:06:37.64" resultid="3856" heatid="10287" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="200" swimtime="00:03:14.15" />
                    <SPLIT distance="300" swimtime="00:04:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-04-08" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="3857">
              <RESULTS>
                <RESULT eventid="1077" points="345" swimtime="00:00:40.03" resultid="3858" heatid="10104" lane="2" entrytime="00:00:37.21" />
                <RESULT eventid="1195" points="286" swimtime="00:00:48.38" resultid="3859" heatid="10135" lane="3" entrytime="00:00:43.71" />
                <RESULT eventid="1324" points="385" swimtime="00:03:46.38" resultid="3860" heatid="10173" lane="5" entrytime="00:03:29.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="519" swimtime="00:00:41.32" resultid="3861" heatid="10189" lane="8" entrytime="00:00:39.33" />
                <RESULT eventid="1465" points="254" swimtime="00:03:27.94" resultid="3862" heatid="10216" lane="2" entrytime="00:03:12.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="443" swimtime="00:00:34.24" resultid="3863" heatid="10250" lane="6" entrytime="00:00:32.30" />
                <RESULT eventid="1654" points="409" swimtime="00:01:40.05" resultid="3864" heatid="10277" lane="4" entrytime="00:01:31.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="3865">
              <RESULTS>
                <RESULT eventid="1141" points="154" swimtime="00:17:35.19" resultid="3866" heatid="10295" lane="4" entrytime="00:17:02.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.30" />
                    <SPLIT distance="200" swimtime="00:04:05.61" />
                    <SPLIT distance="300" swimtime="00:06:18.68" />
                    <SPLIT distance="400" swimtime="00:08:36.61" />
                    <SPLIT distance="500" swimtime="00:10:55.21" />
                    <SPLIT distance="600" swimtime="00:13:13.79" />
                    <SPLIT distance="700" swimtime="00:15:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="182" swimtime="00:01:44.03" resultid="3867" heatid="10141" lane="4" entrytime="00:01:38.00" />
                <RESULT eventid="1308" points="310" swimtime="00:04:01.08" resultid="3868" heatid="10168" lane="1" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="168" swimtime="00:03:55.19" resultid="3869" heatid="10210" lane="6" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="212" swimtime="00:00:45.57" resultid="3870" heatid="10241" lane="5" entrytime="00:00:47.00" />
                <RESULT eventid="1670" points="156" swimtime="00:08:24.99" resultid="3871" heatid="10282" lane="3" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.21" />
                    <SPLIT distance="200" swimtime="00:04:01.43" />
                    <SPLIT distance="300" swimtime="00:06:16.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:34.28" resultid="3872" heatid="10123" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3849" number="1" />
                    <RELAYPOSITION athleteid="3839" number="2" />
                    <RELAYPOSITION athleteid="3865" number="3" />
                    <RELAYPOSITION athleteid="3857" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+100" swimtime="00:02:57.65" resultid="3873" heatid="10267" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3857" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="3865" number="2" />
                    <RELAYPOSITION athleteid="3839" number="3" />
                    <RELAYPOSITION athleteid="3849" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MABIA" name="Masters Białystok" nation="POL">
          <CONTACT email="j.wasilewicz@biaform.com.pl" name="Joanna Wasilewicz" phone="601065257" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-01" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="4212">
              <RESULTS>
                <RESULT eventid="1077" points="641" swimtime="00:00:30.92" resultid="5993" heatid="10109" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1195" points="562" swimtime="00:00:33.94" resultid="5994" heatid="10139" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1324" points="510" swimtime="00:03:08.09" resultid="5995" heatid="10176" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="610" swimtime="00:00:34.78" resultid="5996" heatid="10191" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1574" points="633" swimtime="00:00:28.43" resultid="5997" heatid="10256" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1654" points="491" swimtime="00:01:25.13" resultid="5998" heatid="10280" lane="1" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="4219">
              <RESULTS>
                <RESULT eventid="1077" points="539" swimtime="00:00:34.49" resultid="5999" heatid="10106" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1195" points="479" swimtime="00:00:40.77" resultid="6000" heatid="10136" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1324" points="533" swimtime="00:03:23.14" resultid="6001" heatid="10175" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1369" points="762" swimtime="00:00:36.35" resultid="6002" heatid="10190" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1465" points="504" swimtime="00:02:45.54" resultid="6003" heatid="10217" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="629" swimtime="00:01:26.68" resultid="6004" heatid="10279" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1686" points="466" swimtime="00:06:09.13" resultid="6005" heatid="10289" lane="7" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.11" />
                    <SPLIT distance="200" swimtime="00:02:57.81" />
                    <SPLIT distance="300" swimtime="00:04:33.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Jarosław" gender="M" lastname="Pawlik" nation="POL" athleteid="4226">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="6006" heatid="10103" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="6007" heatid="10149" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="6008" heatid="10186" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="6009" heatid="10235" lane="4" entrytime="00:01:50.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="6010" heatid="10249" lane="3" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="4232">
              <RESULTS>
                <RESULT eventid="1077" points="347" swimtime="00:00:38.95" resultid="6011" heatid="10104" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1162" points="284" swimtime="00:26:41.10" resultid="6012" heatid="10300" lane="2" entrytime="00:29:00.00" />
                <RESULT eventid="1195" points="444" swimtime="00:00:37.83" resultid="6013" heatid="10137" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1292" points="218" swimtime="00:03:55.58" resultid="6014" heatid="10164" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="417" reactiontime="+77" swimtime="00:01:27.03" resultid="6015" heatid="10202" lane="8" entrytime="00:01:26.00" />
                <RESULT eventid="1542" status="DSQ" swimtime="00:01:42.81" resultid="6016" heatid="10236" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="1606" points="344" reactiontime="+85" swimtime="00:03:21.02" resultid="6017" heatid="10263" lane="5" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="4240">
              <RESULTS>
                <RESULT eventid="1061" points="511" swimtime="00:00:38.15" resultid="6018" heatid="10098" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1178" points="577" swimtime="00:00:40.08" resultid="6019" heatid="10129" lane="7" entrytime="00:00:39.90" />
                <RESULT eventid="1212" points="595" swimtime="00:01:15.51" resultid="6020" heatid="10144" lane="5" entrytime="00:01:14.90" />
                <RESULT eventid="1385" points="574" reactiontime="+79" swimtime="00:01:27.99" resultid="6021" heatid="10196" lane="7" entrytime="00:01:29.90" />
                <RESULT eventid="1449" points="471" swimtime="00:02:57.27" resultid="6022" heatid="10212" lane="2" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="601" swimtime="00:00:33.36" resultid="6023" heatid="10244" lane="6" entrytime="00:00:33.90" />
                <RESULT eventid="1590" points="548" reactiontime="+74" swimtime="00:03:18.30" resultid="6024" heatid="10259" lane="3" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="4248">
              <RESULTS>
                <RESULT eventid="1212" points="420" swimtime="00:01:26.82" resultid="6025" heatid="10143" lane="8" entrytime="00:01:25.80" />
                <RESULT eventid="1449" points="387" swimtime="00:03:16.60" resultid="6026" heatid="10211" lane="8" entrytime="00:03:14.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="440" swimtime="00:00:38.30" resultid="6027" heatid="10243" lane="1" entrytime="00:00:37.50" />
                <RESULT eventid="1670" points="382" swimtime="00:07:05.64" resultid="6028" heatid="10283" lane="6" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.48" />
                    <SPLIT distance="200" swimtime="00:03:28.33" />
                    <SPLIT distance="300" swimtime="00:05:18.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="4253">
              <RESULTS>
                <RESULT eventid="1212" points="633" swimtime="00:01:07.61" resultid="6029" heatid="10145" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1449" points="632" swimtime="00:02:25.96" resultid="6030" heatid="10213" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1670" points="661" swimtime="00:05:07.67" resultid="6031" heatid="10285" lane="6" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="200" swimtime="00:02:31.50" />
                    <SPLIT distance="300" swimtime="00:03:50.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TWOPR" name="Tarnowskie WOPR Masters" nation="POL" region="MAL">
          <CONTACT city="zgłobice" email="kacermarcin@o2.pl" name="kacer" phone="607681313" state="MAL" street="rzemieślnicza 24" zip="33-113" />
          <ATHLETES>
            <ATHLETE birthdate="1979-10-26" firstname="Katarzyna" gender="F" lastname="Kacer" nation="POL" athleteid="4266">
              <RESULTS>
                <RESULT eventid="1178" points="326" swimtime="00:00:44.28" resultid="4267" heatid="10128" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1558" points="413" swimtime="00:00:35.68" resultid="4268" heatid="10243" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-15" firstname="Marcin" gender="M" lastname="Kacer" nation="POL" athleteid="4269">
              <RESULTS>
                <RESULT eventid="1077" points="627" swimtime="00:00:29.50" resultid="4270" heatid="10109" lane="4" entrytime="00:00:28.90" />
                <RESULT eventid="1542" points="551" swimtime="00:01:07.95" resultid="4271" heatid="10240" lane="8" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-16" firstname="Maciej" gender="M" lastname="Kacer" nation="POL" athleteid="4272" />
            <ATHLETE birthdate="1975-08-30" firstname="Norbert" gender="M" lastname="Charhouli" nation="POL" athleteid="4273">
              <RESULTS>
                <RESULT eventid="1109" points="186" swimtime="00:03:39.54" resultid="4274" heatid="10117" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="196" swimtime="00:00:47.27" resultid="4275" heatid="10135" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1401" points="201" reactiontime="+82" swimtime="00:01:40.31" resultid="4276" heatid="10200" lane="5" entrytime="00:01:36.00" />
                <RESULT eventid="1606" points="202" reactiontime="+79" swimtime="00:03:36.74" resultid="4277" heatid="10263" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-25" firstname="Adam" gender="M" lastname="Wytrwał" nation="POL" athleteid="4278">
              <RESULTS>
                <RESULT eventid="1162" points="317" swimtime="00:24:56.20" resultid="4279" heatid="10299" lane="2" entrytime="00:26:00.00" />
                <RESULT eventid="1324" points="330" swimtime="00:03:37.38" resultid="4280" heatid="10174" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4281" heatid="10218" lane="5" entrytime="00:02:40.00" />
                <RESULT eventid="1686" points="305" swimtime="00:06:13.21" resultid="4282" heatid="10289" lane="5" entrytime="00:05:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.20" />
                    <SPLIT distance="200" swimtime="00:03:04.25" />
                    <SPLIT distance="300" swimtime="00:04:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="271" swimtime="00:07:32.88" resultid="9054" heatid="10229" lane="3" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.78" />
                    <SPLIT distance="200" swimtime="00:03:48.81" />
                    <SPLIT distance="300" swimtime="00:05:56.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-13" firstname="Barbara" gender="F" lastname="Wytrwał" nation="POL" athleteid="4283">
              <RESULTS>
                <RESULT eventid="1212" points="52" swimtime="00:02:37.18" resultid="4284" heatid="10141" lane="3" entrytime="00:01:50.00" />
                <RESULT eventid="1449" points="46" swimtime="00:06:00.31" resultid="4285" heatid="10210" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="74" swimtime="00:01:04.76" resultid="4286" heatid="10241" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1670" points="60" swimtime="00:11:31.64" resultid="4287" heatid="10282" lane="1" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:52.93" />
                    <SPLIT distance="200" swimtime="00:05:51.36" />
                    <SPLIT distance="300" swimtime="00:08:51.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-24" firstname="Radosław" gender="M" lastname="Jurek" nation="POL" athleteid="4288">
              <RESULTS>
                <RESULT eventid="1077" points="555" swimtime="00:00:30.73" resultid="4289" heatid="10109" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1228" points="404" swimtime="00:01:08.49" resultid="4290" heatid="10155" lane="1" entrytime="00:01:03.00" />
                <RESULT eventid="1465" points="360" swimtime="00:02:36.96" resultid="4291" heatid="10220" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="357" swimtime="00:01:18.51" resultid="4292" heatid="10239" lane="3" entrytime="00:01:09.00" />
                <RESULT eventid="1369" points="439" swimtime="00:00:38.76" resultid="9471" heatid="10183" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="4293">
              <RESULTS>
                <RESULT eventid="1109" points="521" swimtime="00:02:39.92" resultid="4294" heatid="10121" lane="8" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="474" swimtime="00:21:00.78" resultid="4295" heatid="10296" lane="2" entrytime="00:20:00.00" />
                <RESULT eventid="1195" points="484" swimtime="00:00:33.24" resultid="4296" heatid="10140" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1497" points="462" swimtime="00:05:55.15" resultid="4297" heatid="10231" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="200" swimtime="00:02:48.63" />
                    <SPLIT distance="300" swimtime="00:04:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="498" swimtime="00:05:03.59" resultid="4298" heatid="10292" lane="6" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="200" swimtime="00:02:25.96" />
                    <SPLIT distance="300" swimtime="00:03:45.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-07" firstname="Łukasz" gender="M" lastname="Litwora" nation="POL" athleteid="4299">
              <RESULTS>
                <RESULT eventid="1195" points="376" swimtime="00:00:38.05" resultid="4301" heatid="10139" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1228" points="491" swimtime="00:01:05.19" resultid="8053" heatid="10155" lane="6" entrytime="00:01:03.00" />
                <RESULT eventid="1465" points="374" swimtime="00:02:41.12" resultid="8054" heatid="10222" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="532" swimtime="00:00:28.57" resultid="8055" heatid="10255" lane="3" entrytime="00:00:27.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-07" firstname="Gabriela" gender="F" lastname="Gurak" nation="POL" athleteid="4302">
              <RESULTS>
                <RESULT eventid="1308" points="390" swimtime="00:03:32.30" resultid="4303" heatid="10169" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="504" swimtime="00:00:41.80" resultid="4304" heatid="10182" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1638" points="318" swimtime="00:01:44.54" resultid="4305" heatid="10273" lane="1" entrytime="00:01:29.00" />
                <RESULT eventid="1558" points="441" swimtime="00:00:34.90" resultid="9053" heatid="10244" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-01" firstname="Małgorzata" gender="F" lastname="Głowacka" nation="POL" athleteid="4306">
              <RESULTS>
                <RESULT eventid="1352" points="273" swimtime="00:00:59.25" resultid="4307" heatid="10179" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="1558" points="291" swimtime="00:00:46.78" resultid="4308" heatid="10242" lane="8" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-06-18" firstname="Paweł" gender="M" lastname="Pastuszko" nation="POL" athleteid="4309">
              <RESULTS>
                <RESULT eventid="1162" points="162" swimtime="00:30:02.86" resultid="4310" heatid="10301" lane="3" entrytime="00:30:09.00" />
                <RESULT eventid="1324" points="250" swimtime="00:03:44.83" resultid="4311" heatid="10172" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="249" swimtime="00:00:45.74" resultid="4312" heatid="10184" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="1654" status="DSQ" swimtime="00:01:44.14" resultid="4313" heatid="10276" lane="3" entrytime="00:01:40.00" />
                <RESULT eventid="1686" points="148" status="EXH" swimtime="00:07:43.01" resultid="10311" heatid="10286" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.30" />
                    <SPLIT distance="200" swimtime="00:03:46.18" />
                    <SPLIT distance="300" swimtime="00:05:47.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-23" firstname="Mateusz" gender="M" lastname="Dymiter" nation="POL" athleteid="4314">
              <RESULTS>
                <RESULT eventid="1109" points="499" swimtime="00:02:42.73" resultid="4315" heatid="10119" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="349" swimtime="00:22:52.28" resultid="4316" heatid="10298" lane="7" entrytime="00:23:40.00" />
                <RESULT eventid="1228" points="460" swimtime="00:01:05.51" resultid="4317" heatid="10154" lane="7" entrytime="00:01:05.00" />
                <RESULT eventid="1497" points="421" swimtime="00:06:02.68" resultid="4318" heatid="10230" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="200" swimtime="00:02:52.51" />
                    <SPLIT distance="300" swimtime="00:04:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="404" swimtime="00:05:26.47" resultid="4319" heatid="10291" lane="1" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="200" swimtime="00:02:37.35" />
                    <SPLIT distance="300" swimtime="00:04:02.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-09" firstname="Andrzej" gender="M" lastname="Jagiełło" nation="POL" athleteid="4320">
              <RESULTS>
                <RESULT eventid="1574" points="315" swimtime="00:00:37.25" resultid="4321" heatid="10248" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1077" points="170" swimtime="00:00:50.04" resultid="9052" heatid="10102" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-23" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" athleteid="7968">
              <RESULTS>
                <RESULT eventid="1178" points="547" swimtime="00:00:37.22" resultid="7969" heatid="10129" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1385" points="497" reactiontime="+85" swimtime="00:01:20.09" resultid="7970" heatid="10196" lane="2" entrytime="00:01:28.00" />
                <RESULT eventid="1590" points="475" reactiontime="+89" swimtime="00:02:53.20" resultid="7971" heatid="10260" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+80" swimtime="00:01:59.79" resultid="4324" heatid="10161" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4293" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4272" number="2" />
                    <RELAYPOSITION athleteid="4269" number="3" />
                    <RELAYPOSITION athleteid="4299" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:01:52.15" resultid="4325" heatid="10208" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4299" number="1" />
                    <RELAYPOSITION athleteid="4288" number="2" />
                    <RELAYPOSITION athleteid="4314" number="3" />
                    <RELAYPOSITION athleteid="4293" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+75" swimtime="00:02:40.88" resultid="4326" heatid="10160" lane="2" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4320" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4309" number="2" />
                    <RELAYPOSITION athleteid="4288" number="3" />
                    <RELAYPOSITION athleteid="4278" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:02:11.96" resultid="4327" heatid="10207" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4273" number="1" />
                    <RELAYPOSITION athleteid="4320" number="2" />
                    <RELAYPOSITION athleteid="4278" number="3" />
                    <RELAYPOSITION athleteid="4269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1417" swimtime="00:03:05.64" resultid="4322" heatid="10206" lane="1" entrytime="00:03:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4283" number="1" />
                    <RELAYPOSITION athleteid="4306" number="2" />
                    <RELAYPOSITION athleteid="4266" number="3" />
                    <RELAYPOSITION athleteid="4302" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1244" reactiontime="+116" swimtime="00:03:28.29" resultid="4323" heatid="10159" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:08.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4283" number="1" reactiontime="+116" />
                    <RELAYPOSITION athleteid="4306" number="2" />
                    <RELAYPOSITION athleteid="4302" number="3" />
                    <RELAYPOSITION athleteid="4266" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+83" swimtime="00:02:14.77" resultid="4328" heatid="10269" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4293" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="4302" number="2" />
                    <RELAYPOSITION athleteid="4269" number="3" />
                    <RELAYPOSITION athleteid="7968" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" swimtime="00:02:04.48" resultid="4329" heatid="10123" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4269" number="1" />
                    <RELAYPOSITION athleteid="4266" number="2" />
                    <RELAYPOSITION athleteid="4302" number="3" />
                    <RELAYPOSITION athleteid="4288" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1622" swimtime="00:02:50.77" resultid="4330" heatid="10267" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4266" number="1" />
                    <RELAYPOSITION athleteid="4288" number="2" />
                    <RELAYPOSITION athleteid="4306" number="3" />
                    <RELAYPOSITION athleteid="4278" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" swimtime="00:02:56.20" resultid="4331" heatid="10123" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4283" number="1" />
                    <RELAYPOSITION athleteid="4306" number="2" />
                    <RELAYPOSITION athleteid="4278" number="3" />
                    <RELAYPOSITION athleteid="4314" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MATOR" name="Toruńczyk Masters Toruń" nation="POL" region="KUJ" shortname="Masters Toruń">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Bażyńskich 9/17" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="4352">
              <RESULTS>
                <RESULT eventid="1077" points="385" swimtime="00:00:41.72" resultid="4353" heatid="10102" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1109" points="383" swimtime="00:03:41.78" resultid="4354" heatid="10116" lane="8" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="263" swimtime="00:00:52.17" resultid="4355" heatid="10134" lane="8" entrytime="00:00:53.00" />
                <RESULT eventid="1324" points="392" swimtime="00:04:01.09" resultid="4356" heatid="10171" lane="2" entrytime="00:03:56.00" />
                <RESULT eventid="1369" points="299" swimtime="00:00:51.21" resultid="4357" heatid="10185" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1401" points="248" reactiontime="+102" swimtime="00:01:57.01" resultid="4358" heatid="10199" lane="7" entrytime="00:01:59.00" />
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="4359" heatid="10236" lane="1" entrytime="00:01:49.00" />
                <RESULT eventid="1654" points="350" swimtime="00:01:52.06" resultid="4360" heatid="10275" lane="3" entrytime="00:01:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Sławomir" gender="M" lastname="Predki" nation="POL" athleteid="4361">
              <RESULTS>
                <RESULT eventid="1077" points="723" swimtime="00:00:28.00" resultid="4362" heatid="10110" lane="5" entrytime="00:00:26.49" />
                <RESULT eventid="1109" points="627" swimtime="00:02:26.55" resultid="4363" heatid="10122" lane="4" entrytime="00:02:14.94">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="697" swimtime="00:00:57.98" resultid="4364" heatid="10158" lane="6" entrytime="00:00:57.09" />
                <RESULT eventid="1324" points="660" swimtime="00:02:42.84" resultid="4365" heatid="10177" lane="6" entrytime="00:02:47.46">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="143" swimtime="00:00:55.09" resultid="4366" heatid="10192" lane="3" entrytime="00:00:31.84" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4367" heatid="10231" lane="4" entrytime="00:04:46.97" />
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="4368" heatid="10240" lane="4" entrytime="00:01:00.11" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="4369" heatid="10281" lane="5" entrytime="00:01:11.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="4370">
              <RESULTS>
                <RESULT eventid="1093" points="414" swimtime="00:03:06.37" resultid="4371" heatid="10112" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="328" swimtime="00:12:40.34" resultid="4372" heatid="10293" lane="2" entrytime="00:12:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="200" swimtime="00:03:00.23" />
                    <SPLIT distance="300" swimtime="00:04:39.01" />
                    <SPLIT distance="400" swimtime="00:06:17.70" />
                    <SPLIT distance="500" swimtime="00:07:54.17" />
                    <SPLIT distance="600" swimtime="00:09:29.82" />
                    <SPLIT distance="700" swimtime="00:11:06.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="466" swimtime="00:01:11.97" resultid="4373" heatid="10145" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1308" points="323" swimtime="00:03:41.27" resultid="4374" heatid="10167" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="266" reactiontime="+97" swimtime="00:01:39.56" resultid="4375" heatid="10196" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1449" points="447" swimtime="00:02:42.22" resultid="4376" heatid="10212" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="369" reactiontime="+83" swimtime="00:03:08.97" resultid="4377" heatid="10260" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="351" swimtime="00:05:59.43" resultid="4378" heatid="10284" lane="4" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                    <SPLIT distance="200" swimtime="00:02:58.58" />
                    <SPLIT distance="300" swimtime="00:04:31.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="4379">
              <RESULTS>
                <RESULT eventid="1077" points="471" swimtime="00:00:32.45" resultid="7962" heatid="10106" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1109" points="382" swimtime="00:02:57.33" resultid="4381" heatid="10118" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="308" swimtime="00:03:06.26" resultid="4382" heatid="10165" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="351" swimtime="00:02:38.17" resultid="4383" heatid="10218" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="364" swimtime="00:06:24.61" resultid="4384" heatid="10229" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.12" />
                    <SPLIT distance="200" swimtime="00:03:13.72" />
                    <SPLIT distance="300" swimtime="00:05:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="352" swimtime="00:01:18.87" resultid="4385" heatid="10238" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1686" status="DNS" swimtime="00:00:00.00" resultid="4386" heatid="10289" lane="4" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="4387">
              <RESULTS>
                <RESULT eventid="1228" points="644" swimtime="00:00:59.53" resultid="4388" heatid="10157" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1401" points="622" reactiontime="+71" swimtime="00:01:08.87" resultid="4389" heatid="10204" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1606" points="531" reactiontime="+84" swimtime="00:02:36.99" resultid="4390" heatid="10265" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Marta" gender="F" lastname="Lord" nation="POL" athleteid="4391">
              <RESULTS>
                <RESULT eventid="1178" points="601" swimtime="00:00:36.12" resultid="4392" heatid="10130" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1212" points="516" swimtime="00:01:12.35" resultid="4393" heatid="10145" lane="7" entrytime="00:01:11.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1385" points="623" reactiontime="+85" swimtime="00:01:16.70" resultid="4394" heatid="10197" lane="1" entrytime="00:01:19.00" />
                <RESULT eventid="1449" points="507" swimtime="00:02:37.08" resultid="4395" heatid="10213" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1590" points="590" reactiontime="+90" swimtime="00:02:45.84" resultid="4396" heatid="10260" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Karol" gender="M" lastname="Twarowski" nation="POL" athleteid="4397">
              <RESULTS>
                <RESULT eventid="1077" points="637" swimtime="00:00:29.35" resultid="4398" heatid="10105" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1109" points="695" swimtime="00:02:25.28" resultid="4399" heatid="10120" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="665" swimtime="00:00:58.00" resultid="4400" heatid="10157" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1324" points="592" swimtime="00:02:47.35" resultid="4401" heatid="10170" lane="2" />
                <RESULT eventid="1401" points="545" reactiontime="+100" swimtime="00:01:09.34" resultid="4402" heatid="10203" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="1497" points="650" swimtime="00:05:17.02" resultid="4403" heatid="10227" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="200" swimtime="00:02:33.96" />
                    <SPLIT distance="300" swimtime="00:04:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="268" reactiontime="+114" swimtime="00:03:15.93" resultid="4404" heatid="10266" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="608" swimtime="00:04:44.01" resultid="4405" heatid="10286" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="200" swimtime="00:02:17.99" />
                    <SPLIT distance="300" swimtime="00:03:31.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="4406">
              <RESULTS>
                <RESULT eventid="1109" status="DSQ" swimtime="00:03:42.02" resultid="4407" heatid="10116" lane="1" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="496" swimtime="00:03:42.89" resultid="4408" heatid="10172" lane="2" entrytime="00:03:42.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="493" swimtime="00:00:43.34" resultid="4409" heatid="10186" lane="5" entrytime="00:00:44.20" />
                <RESULT eventid="1654" points="485" swimtime="00:01:40.48" resultid="4410" heatid="10277" lane="1" entrytime="00:01:37.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="4411">
              <RESULTS>
                <RESULT eventid="1077" points="645" swimtime="00:00:35.14" resultid="4412" heatid="10105" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1109" points="487" swimtime="00:03:24.72" resultid="4413" heatid="10117" lane="5" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="603" swimtime="00:01:13.82" resultid="4414" heatid="10150" lane="4" entrytime="00:01:13.50" />
                <RESULT eventid="1369" points="484" swimtime="00:00:43.62" resultid="4415" heatid="10188" lane="1" entrytime="00:00:40.50" />
                <RESULT eventid="1497" points="455" swimtime="00:07:32.72" resultid="4416" heatid="10228" lane="4" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.52" />
                    <SPLIT distance="200" swimtime="00:03:54.18" />
                    <SPLIT distance="300" swimtime="00:05:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="470" swimtime="00:01:30.08" resultid="4417" heatid="10237" lane="6" entrytime="00:01:26.60" />
                <RESULT eventid="1574" points="606" swimtime="00:00:32.24" resultid="4418" heatid="10251" lane="7" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Magdalena" gender="F" lastname="Bolewska" nation="POL" athleteid="4419">
              <RESULTS>
                <RESULT eventid="1061" points="635" swimtime="00:00:33.91" resultid="4420" heatid="10095" lane="4" />
                <RESULT eventid="1093" points="598" swimtime="00:02:48.49" resultid="4421" heatid="10113" lane="6" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="490" swimtime="00:00:38.62" resultid="4422" heatid="10129" lane="5" entrytime="00:00:38.15" />
                <RESULT eventid="1352" points="640" swimtime="00:00:39.54" resultid="4423" heatid="10182" lane="3" entrytime="00:00:37.80" />
                <RESULT eventid="1558" points="617" swimtime="00:00:31.00" resultid="4424" heatid="10245" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1638" points="540" swimtime="00:01:26.81" resultid="4425" heatid="10273" lane="2" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+71" swimtime="00:02:09.55" resultid="4428" heatid="10161" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4387" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4361" number="2" />
                    <RELAYPOSITION athleteid="4411" number="3" />
                    <RELAYPOSITION athleteid="4397" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:01:55.65" resultid="4429" heatid="10208" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4387" number="1" />
                    <RELAYPOSITION athleteid="4411" number="2" />
                    <RELAYPOSITION athleteid="4397" number="3" />
                    <RELAYPOSITION athleteid="4379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+90" swimtime="00:02:10.48" resultid="4426" heatid="10269" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4391" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="4419" number="2" />
                    <RELAYPOSITION athleteid="4397" number="3" />
                    <RELAYPOSITION athleteid="4387" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1125" swimtime="00:01:54.71" resultid="4427" heatid="10125" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4419" number="1" />
                    <RELAYPOSITION athleteid="4391" number="2" />
                    <RELAYPOSITION athleteid="4397" number="3" />
                    <RELAYPOSITION athleteid="4361" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="VIELB" name="Victory Masters Elbląg" nation="POL" shortname="Masters Elbląg">
          <CONTACT city="ELBLĄG" email="lateccy@o2.pl" name="LATECKI GRZEGORZ" street="ŁOKIETKA 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1966-06-06" firstname="ANDRZEJ" gender="M" lastname="PASIECZNY" nation="POL" athleteid="4438">
              <RESULTS>
                <RESULT eventid="1077" points="799" swimtime="00:00:29.51" resultid="7679" heatid="10108" lane="5" entrytime="00:00:30.24" />
                <RESULT eventid="1292" status="DNF" swimtime="00:02:39.80" resultid="7680" heatid="10166" lane="6" entrytime="00:02:25.65">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="747" swimtime="00:02:15.04" resultid="7681" heatid="10223" lane="7" entrytime="00:02:12.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="820" swimtime="00:01:05.53" resultid="7682" heatid="10240" lane="1" entrytime="00:01:03.83" />
                <RESULT eventid="1686" points="741" swimtime="00:04:50.39" resultid="7683" heatid="10292" lane="2" entrytime="00:04:47.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.51" />
                    <SPLIT distance="200" swimtime="00:02:25.56" />
                    <SPLIT distance="300" swimtime="00:03:39.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-18" firstname="TOMASZ" gender="M" lastname="GLEB" nation="POL" athleteid="4444">
              <RESULTS>
                <RESULT eventid="1162" points="483" swimtime="00:22:20.71" resultid="7684" heatid="10297" lane="3" entrytime="00:21:25.01" />
                <RESULT eventid="1228" points="535" swimtime="00:01:07.43" resultid="7685" heatid="10153" lane="7" entrytime="00:01:06.05" />
                <RESULT eventid="1324" points="476" swimtime="00:03:17.10" resultid="7686" heatid="10174" lane="1" entrytime="00:03:20.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="534" swimtime="00:02:31.07" resultid="7687" heatid="10221" lane="8" entrytime="00:02:25.49">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="508" swimtime="00:00:30.74" resultid="7688" heatid="10252" lane="4" entrytime="00:00:29.34" />
                <RESULT eventid="1686" points="515" swimtime="00:05:27.82" resultid="7689" heatid="10290" lane="6" entrytime="00:05:23.17">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="200" swimtime="00:02:39.95" />
                    <SPLIT distance="300" swimtime="00:04:05.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="KAROLINA" gender="F" lastname="KARAŚ" nation="POL" athleteid="4456">
              <RESULTS>
                <RESULT eventid="1141" points="273" swimtime="00:14:15.42" resultid="7690" heatid="10294" lane="8" entrytime="00:16:15.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.30" />
                    <SPLIT distance="200" swimtime="00:03:28.98" />
                    <SPLIT distance="300" swimtime="00:05:18.27" />
                    <SPLIT distance="400" swimtime="00:07:06.23" />
                    <SPLIT distance="500" swimtime="00:08:53.00" />
                    <SPLIT distance="600" swimtime="00:10:40.46" />
                    <SPLIT distance="700" swimtime="00:12:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="229" swimtime="00:01:33.79" resultid="7691" heatid="10142" lane="8" entrytime="00:01:37.25" />
                <RESULT eventid="1449" points="225" swimtime="00:03:21.84" resultid="7692" heatid="10210" lane="3" entrytime="00:03:43.27">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="7693" heatid="10242" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1670" points="273" swimtime="00:06:49.62" resultid="7694" heatid="10283" lane="1" entrytime="00:07:20.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.42" />
                    <SPLIT distance="200" swimtime="00:03:22.91" />
                    <SPLIT distance="300" swimtime="00:05:06.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="GRZEGORZ" gender="M" lastname="LATECKI" nation="POL" athleteid="4462">
              <RESULTS>
                <RESULT eventid="1077" points="830" swimtime="00:00:29.14" resultid="7695" heatid="10109" lane="6" entrytime="00:00:29.80" />
                <RESULT eventid="1228" points="647" swimtime="00:01:03.30" resultid="7696" heatid="10155" lane="5" entrytime="00:01:02.60" />
                <RESULT eventid="1324" points="565" swimtime="00:03:06.21" resultid="7697" heatid="10176" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="455" swimtime="00:00:39.94" resultid="7698" heatid="10190" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1574" points="693" swimtime="00:00:27.72" resultid="7700" heatid="10255" lane="6" entrytime="00:00:27.80" />
                <RESULT eventid="1606" points="578" reactiontime="+84" swimtime="00:02:49.09" resultid="7701" heatid="10265" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="7702">
              <RESULTS>
                <RESULT eventid="1178" points="206" swimtime="00:01:02.72" resultid="7703" heatid="10126" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1212" points="220" swimtime="00:01:53.38" resultid="7704" heatid="10141" lane="6" entrytime="00:02:05.00" />
                <RESULT eventid="1352" points="126" swimtime="00:01:16.55" resultid="7705" heatid="10179" lane="2" entrytime="00:01:07.00" />
                <RESULT eventid="1385" points="183" reactiontime="+98" swimtime="00:02:24.25" resultid="7706" heatid="10193" lane="6" entrytime="00:02:33.00" />
                <RESULT eventid="1558" points="267" swimtime="00:00:48.16" resultid="7707" heatid="10241" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1638" points="178" swimtime="00:02:35.10" resultid="7708" heatid="10271" lane="7" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZUWA" name="AZS Uniwersytet Warszawski" nation="POL" shortname="AZS UW">
          <ATHLETES>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="4476">
              <RESULTS>
                <RESULT eventid="1195" points="441" swimtime="00:00:33.43" resultid="4477" heatid="10132" lane="2" />
                <RESULT eventid="1228" points="596" swimtime="00:00:58.66" resultid="4478" heatid="10158" lane="7" entrytime="00:00:58.30" />
                <RESULT eventid="1465" points="457" swimtime="00:02:19.79" resultid="4479" heatid="10220" lane="5" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="609" swimtime="00:01:03.29" resultid="4480" heatid="10234" lane="5" />
                <RESULT eventid="1574" points="534" swimtime="00:00:27.50" resultid="4481" heatid="10257" lane="3" entrytime="00:00:25.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REWRO" name="Redeco Wrocław" nation="POL">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="4488">
              <RESULTS>
                <RESULT eventid="1077" points="733" swimtime="00:00:30.75" resultid="4489" heatid="10108" lane="3" entrytime="00:00:30.30" />
                <RESULT eventid="1109" points="967" swimtime="00:02:30.23" resultid="4490" heatid="10122" lane="1" entrytime="00:02:29.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="878" swimtime="00:00:31.97" resultid="4491" heatid="10140" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="4492" heatid="10189" lane="5" entrytime="00:00:37.37" />
                <RESULT eventid="1401" points="907" reactiontime="+78" swimtime="00:01:09.39" resultid="4493" heatid="10205" lane="8" entrytime="00:01:08.08" />
                <RESULT eventid="1606" points="985" reactiontime="+75" swimtime="00:02:29.67" resultid="4494" heatid="10266" lane="6" entrytime="00:02:28.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="742" swimtime="00:01:20.38" resultid="4495" heatid="10280" lane="7" entrytime="00:01:19.64" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="4496">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="4497" heatid="10099" lane="3" entrytime="00:00:32.88" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1308" points="790" swimtime="00:02:47.83" resultid="4498" heatid="10169" lane="4" entrytime="00:02:47.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="883" swimtime="00:00:34.68" resultid="4499" heatid="10182" lane="4" entrytime="00:00:34.88" />
                <RESULT eventid="1638" points="811" swimtime="00:01:16.56" resultid="4500" heatid="10273" lane="4" entrytime="00:01:18.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-13" firstname="Kazimiera" gender="F" lastname="Syguła" nation="POL" athleteid="4501">
              <RESULTS>
                <RESULT eventid="1178" points="438" swimtime="00:00:54.16" resultid="4502" heatid="10126" lane="4" entrytime="00:00:57.44" />
                <RESULT eventid="1212" points="293" swimtime="00:01:55.91" resultid="4503" heatid="10141" lane="5" entrytime="00:01:49.07" />
                <RESULT eventid="1385" points="480" reactiontime="+84" swimtime="00:01:58.08" resultid="4504" heatid="10194" lane="7" entrytime="00:01:57.11" />
                <RESULT eventid="1558" points="371" swimtime="00:00:48.41" resultid="4505" heatid="10241" lane="3" entrytime="00:00:47.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-08" firstname="Mariusz" gender="M" lastname="Bazanowski" nation="POL" athleteid="4506">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="4507" heatid="10104" lane="1" entrytime="00:00:37.88" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4508" heatid="10153" lane="6" entrytime="00:01:06.00" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4509" heatid="10221" lane="2" entrytime="00:02:24.00" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="4510" heatid="10253" lane="6" entrytime="00:00:28.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="4511">
              <RESULTS>
                <RESULT eventid="1077" points="465" swimtime="00:00:32.72" resultid="4512" heatid="10106" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1228" points="447" swimtime="00:01:06.12" resultid="4513" heatid="10155" lane="7" entrytime="00:01:03.00" />
                <RESULT eventid="1542" points="282" swimtime="00:01:24.63" resultid="4514" heatid="10237" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="1574" points="476" swimtime="00:00:29.11" resultid="4515" heatid="10254" lane="7" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Wojciech" gender="M" lastname="Sobczak" nation="POL" athleteid="4516">
              <RESULTS>
                <RESULT eventid="1077" points="239" swimtime="00:00:40.70" resultid="4517" heatid="10105" lane="5" entrytime="00:00:34.55" />
                <RESULT eventid="1109" points="272" swimtime="00:03:18.59" resultid="4518" heatid="10118" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="351" swimtime="00:01:11.77" resultid="4519" heatid="10152" lane="3" entrytime="00:01:08.08" />
                <RESULT eventid="1324" points="296" swimtime="00:03:30.71" resultid="4520" heatid="10173" lane="8" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="362" swimtime="00:00:41.33" resultid="4521" heatid="10188" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1497" points="256" swimtime="00:07:12.64" resultid="4522" heatid="10230" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.12" />
                    <SPLIT distance="200" swimtime="00:03:40.68" />
                    <SPLIT distance="300" swimtime="00:05:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="168" swimtime="00:01:40.92" resultid="4523" heatid="10238" lane="4" entrytime="00:01:15.68" />
                <RESULT eventid="1654" points="288" swimtime="00:01:38.16" resultid="4524" heatid="10276" lane="2" entrytime="00:01:40.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-23" firstname="Agata" gender="F" lastname="Sobczak" nation="POL" athleteid="4525">
              <RESULTS>
                <RESULT eventid="1141" points="221" swimtime="00:15:18.75" resultid="4526" heatid="10294" lane="2" entrytime="00:14:14.14">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.46" />
                    <SPLIT distance="200" swimtime="00:03:36.68" />
                    <SPLIT distance="300" swimtime="00:05:32.72" />
                    <SPLIT distance="400" swimtime="00:07:29.25" />
                    <SPLIT distance="500" swimtime="00:09:26.82" />
                    <SPLIT distance="600" swimtime="00:11:25.97" />
                    <SPLIT distance="700" swimtime="00:13:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="229" swimtime="00:01:33.81" resultid="4527" heatid="10143" lane="1" entrytime="00:01:25.24" />
                <RESULT eventid="1449" points="212" swimtime="00:03:25.98" resultid="4528" heatid="10211" lane="4" entrytime="00:03:01.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="155" swimtime="00:01:57.39" resultid="4529" heatid="10232" lane="5" entrytime="00:01:45.00" />
                <RESULT eventid="1670" points="214" swimtime="00:07:24.34" resultid="4530" heatid="10283" lane="7" entrytime="00:07:07.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.66" />
                    <SPLIT distance="200" swimtime="00:03:35.11" />
                    <SPLIT distance="300" swimtime="00:05:32.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-24" firstname="Małgorzata" gender="F" lastname="Garbarek" nation="POL" athleteid="4531">
              <RESULTS>
                <RESULT eventid="1061" points="359" swimtime="00:00:40.56" resultid="4532" heatid="10098" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1212" points="349" swimtime="00:01:22.41" resultid="4533" heatid="10143" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="1352" points="343" swimtime="00:00:47.52" resultid="4534" heatid="10180" lane="4" entrytime="00:00:44.44" />
                <RESULT eventid="1558" points="369" swimtime="00:00:37.03" resultid="4535" heatid="10244" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1638" status="DNS" swimtime="00:00:00.00" resultid="4536" heatid="10272" lane="1" entrytime="00:01:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-13" firstname="Agata" gender="F" lastname="Grochowska" nation="POL" athleteid="4537">
              <RESULTS>
                <RESULT eventid="1061" points="270" swimtime="00:00:45.88" resultid="4538" heatid="10096" lane="3" entrytime="00:00:54.22" />
                <RESULT eventid="1141" points="223" swimtime="00:15:33.16" resultid="4539" heatid="10294" lane="7" entrytime="00:15:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="200" swimtime="00:03:36.23" />
                    <SPLIT distance="300" swimtime="00:05:35.05" />
                    <SPLIT distance="400" swimtime="00:09:37.23" />
                    <SPLIT distance="500" swimtime="00:11:39.81" />
                    <SPLIT distance="600" swimtime="00:13:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="293" swimtime="00:00:47.30" resultid="4540" heatid="10127" lane="3" entrytime="00:00:45.21" />
                <RESULT eventid="1212" points="246" swimtime="00:01:34.09" resultid="4541" heatid="10143" lane="6" entrytime="00:01:20.26" />
                <RESULT eventid="1385" points="256" reactiontime="+78" swimtime="00:01:45.00" resultid="4542" heatid="10195" lane="8" entrytime="00:01:38.00" />
                <RESULT eventid="1449" points="238" swimtime="00:03:29.60" resultid="4543" heatid="10212" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="261" reactiontime="+73" swimtime="00:03:47.36" resultid="4544" heatid="10258" lane="4" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="207" swimtime="00:07:39.28" resultid="4545" heatid="10282" lane="5" entrytime="00:07:58.88">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.49" />
                    <SPLIT distance="200" swimtime="00:03:46.79" />
                    <SPLIT distance="300" swimtime="00:05:46.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Dariusz" gender="M" lastname="Patrzałek" nation="POL" athleteid="4546">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="4547" heatid="10134" lane="6" entrytime="00:00:49.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4548" heatid="10148" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="4549" heatid="10185" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4550" heatid="10200" lane="7" entrytime="00:01:44.44" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="4551" heatid="10247" lane="2" entrytime="00:00:42.22" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="4552" heatid="10275" lane="6" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-28" firstname="Przemysław" gender="M" lastname="Matuszek" nation="POL" athleteid="4553">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="4554" heatid="10109" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4555" heatid="10154" lane="3" entrytime="00:01:05.00" />
                <RESULT eventid="1465" points="361" swimtime="00:02:36.72" resultid="4556" heatid="10220" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="4557" heatid="10239" lane="8" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="4558">
              <RESULTS>
                <RESULT eventid="1061" points="277" swimtime="00:00:44.84" resultid="4559" heatid="10097" lane="4" entrytime="00:00:42.44" />
                <RESULT eventid="1093" points="294" swimtime="00:03:33.78" resultid="4560" heatid="10111" lane="4" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="350" swimtime="00:00:44.40" resultid="4561" heatid="10129" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1212" points="350" swimtime="00:01:21.83" resultid="4562" heatid="10143" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1385" points="261" reactiontime="+62" swimtime="00:01:41.23" resultid="4563" heatid="10194" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="1449" points="276" swimtime="00:03:13.24" resultid="4564" heatid="10211" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="203" swimtime="00:01:49.85" resultid="4565" heatid="10233" lane="8" entrytime="00:01:34.44" />
                <RESULT eventid="1670" points="232" swimtime="00:07:15.82" resultid="4566" heatid="10284" lane="8" entrytime="00:06:34.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.21" />
                    <SPLIT distance="200" swimtime="00:03:27.56" />
                    <SPLIT distance="300" swimtime="00:05:24.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1260" status="DNS" swimtime="00:00:00.00" resultid="4571" heatid="10161" lane="8" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4488" number="1" />
                    <RELAYPOSITION athleteid="4553" number="2" />
                    <RELAYPOSITION athleteid="4516" number="3" />
                    <RELAYPOSITION athleteid="4506" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="4572" heatid="10208" lane="1" entrytime="00:01:59.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4488" number="1" />
                    <RELAYPOSITION athleteid="4511" number="2" />
                    <RELAYPOSITION athleteid="4553" number="3" />
                    <RELAYPOSITION athleteid="4506" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1244" status="DNS" swimtime="00:00:00.00" resultid="4573" heatid="10159" lane="4" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4537" number="1" />
                    <RELAYPOSITION athleteid="4531" number="2" />
                    <RELAYPOSITION athleteid="4496" number="3" />
                    <RELAYPOSITION athleteid="4558" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="4574" heatid="10206" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4537" number="1" />
                    <RELAYPOSITION athleteid="4558" number="2" />
                    <RELAYPOSITION athleteid="4496" number="3" />
                    <RELAYPOSITION athleteid="4531" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:02.16" resultid="4567" heatid="10125" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4531" number="1" />
                    <RELAYPOSITION athleteid="4496" number="2" />
                    <RELAYPOSITION athleteid="4488" number="3" />
                    <RELAYPOSITION athleteid="4553" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="4570" heatid="10125" lane="2" entrytime="00:02:02.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4511" number="1" />
                    <RELAYPOSITION athleteid="4506" number="2" />
                    <RELAYPOSITION athleteid="4501" number="3" />
                    <RELAYPOSITION athleteid="4558" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TAKAS" name="Takas" nation="LTU">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Viktoras Snieska" phone="+37068297778" street="Lentvario g. 19-1" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="yliene" nation="LTU" athleteid="4587">
              <RESULTS>
                <RESULT eventid="1178" points="504" swimtime="00:00:51.68" resultid="4588" heatid="10127" lane="7" entrytime="00:00:49.85" />
                <RESULT eventid="1385" points="424" reactiontime="+89" swimtime="00:02:03.04" resultid="4589" heatid="10194" lane="2" entrytime="00:01:56.00" />
                <RESULT eventid="1590" points="358" reactiontime="+145" swimtime="00:04:44.05" resultid="4590" heatid="10258" lane="3" entrytime="00:04:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="316" swimtime="00:08:40.91" resultid="4591" heatid="10283" lane="8" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:04:17.67" />
                    <SPLIT distance="300" swimtime="00:06:32.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1927-04-21" firstname="Vladas" gender="M" lastname="vimbaras" nation="LTU" athleteid="4592">
              <RESULTS>
                <RESULT eventid="1195" points="212" swimtime="00:01:16.25" resultid="4593" heatid="10132" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1574" points="388" swimtime="00:00:51.47" resultid="4594" heatid="10246" lane="4" entrytime="00:00:50.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-08" firstname="Viktoras" gender="M" lastname="snieska" nation="LTU" athleteid="4595">
              <RESULTS>
                <RESULT eventid="1109" points="635" swimtime="00:03:21.19" resultid="4596" heatid="10116" lane="4" entrytime="00:03:37.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="600" swimtime="00:00:41.81" resultid="4597" heatid="10136" lane="5" entrytime="00:00:40.23" />
                <RESULT eventid="1228" points="652" swimtime="00:01:16.15" resultid="4598" heatid="10151" lane="7" entrytime="00:01:12.76" />
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="4599" heatid="10163" lane="6" entrytime="00:04:24.82" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="4600" heatid="10171" lane="1" entrytime="00:03:58.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:04:01.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="4601" heatid="10186" lane="1" entrytime="00:00:45.41" />
                <RESULT eventid="1401" points="603" reactiontime="+100" swimtime="00:01:34.62" resultid="4602" heatid="10201" lane="1" entrytime="00:01:31.04" />
                <RESULT eventid="1465" points="528" swimtime="00:03:03.91" resultid="4603" heatid="10217" lane="7" entrytime="00:02:51.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4604" heatid="10228" lane="1" entrytime="00:07:41.03" />
                <RESULT eventid="1574" points="633" swimtime="00:00:32.92" resultid="4605" heatid="10249" lane="5" entrytime="00:00:33.40" />
                <RESULT eventid="1606" points="516" reactiontime="+161" swimtime="00:03:37.53" resultid="4606" heatid="10263" lane="3" entrytime="00:03:21.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1686" points="501" swimtime="00:06:51.68" resultid="4607" heatid="10288" lane="8" entrytime="00:06:18.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.17" />
                    <SPLIT distance="200" swimtime="00:03:27.13" />
                    <SPLIT distance="300" swimtime="00:05:10.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-09" firstname="Nijole" gender="F" lastname="macerinskiene" nation="LTU" athleteid="4608">
              <RESULTS>
                <RESULT eventid="1061" points="306" swimtime="00:00:49.77" resultid="4609" heatid="10096" lane="5" entrytime="00:00:52.10" />
                <RESULT eventid="1352" points="380" swimtime="00:00:53.07" resultid="4610" heatid="10179" lane="4" entrytime="00:00:54.30" />
                <RESULT eventid="1558" points="419" swimtime="00:00:41.45" resultid="4611" heatid="10242" lane="7" entrytime="00:00:42.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+92" swimtime="00:03:24.49" resultid="9475" heatid="10268" lane="1" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4587" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="4595" number="2" />
                    <RELAYPOSITION athleteid="4592" number="3" />
                    <RELAYPOSITION athleteid="4608" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" swimtime="00:02:57.90" resultid="9476" heatid="10124" lane="8" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4608" number="1" />
                    <RELAYPOSITION athleteid="4587" number="2" />
                    <RELAYPOSITION athleteid="4595" number="3" />
                    <RELAYPOSITION athleteid="4592" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TRPRA" name="Triva Praha" nation="CZE">
          <CONTACT email="benova.dana@seznam.cz" name="Triva Praha" phone="+420728212656" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Benova" nation="CZE" athleteid="4613">
              <RESULTS>
                <RESULT eventid="1385" points="253" reactiontime="+82" swimtime="00:02:09.54" resultid="4614" heatid="10194" lane="1" entrytime="00:02:03.80" entrycourse="LCM" />
                <RESULT eventid="1449" points="189" swimtime="00:04:22.10" resultid="4615" heatid="10209" lane="5" entrytime="00:04:23.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:08.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="289" reactiontime="+83" swimtime="00:04:40.61" resultid="4616" heatid="10258" lane="6" entrytime="00:04:36.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:20.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="218" swimtime="00:09:14.12" resultid="4617" heatid="10282" lane="6" entrytime="00:08:47.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:11.40" />
                    <SPLIT distance="200" swimtime="00:04:32.29" />
                    <SPLIT distance="300" swimtime="00:06:55.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-10" firstname="Vaclav" gender="M" lastname="Valtr" nation="CZE" athleteid="4618">
              <RESULTS>
                <RESULT eventid="1401" points="613" reactiontime="+76" swimtime="00:01:19.51" resultid="4619" heatid="10203" lane="2" entrytime="00:01:16.50" entrycourse="LCM" />
                <RESULT eventid="1497" points="669" swimtime="00:06:26.26" resultid="4620" heatid="10229" lane="5" entrytime="00:06:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="200" swimtime="00:03:12.21" />
                    <SPLIT distance="300" swimtime="00:04:59.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="599" reactiontime="+91" swimtime="00:02:58.59" resultid="4621" heatid="10265" lane="1" entrytime="00:02:52.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="592" swimtime="00:01:28.47" resultid="4622" heatid="10279" lane="8" entrytime="00:01:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKAT" name="UKS Wodnik 29 Katowice" nation="POL" shortname="Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas" phone="662 297 707" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4624">
              <RESULTS>
                <RESULT eventid="1109" points="548" swimtime="00:03:01.54" resultid="4625" heatid="10119" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="595" swimtime="00:03:11.63" resultid="4626" heatid="10175" lane="3" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="662" swimtime="00:00:36.93" resultid="4627" heatid="10190" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1654" points="621" swimtime="00:01:25.27" resultid="4628" heatid="10279" lane="4" entrytime="00:01:24.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="4629">
              <RESULTS>
                <RESULT eventid="1077" points="763" swimtime="00:00:33.23" resultid="4630" heatid="10106" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1228" points="529" swimtime="00:01:17.10" resultid="4631" heatid="10150" lane="6" entrytime="00:01:14.00" />
                <RESULT eventid="1292" points="352" swimtime="00:03:49.37" resultid="4632" heatid="10164" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="449" swimtime="00:03:04.28" resultid="4633" heatid="10217" lane="8" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="465" swimtime="00:01:30.44" resultid="4634" heatid="10237" lane="2" entrytime="00:01:28.00" />
                <RESULT eventid="1574" points="566" swimtime="00:00:32.99" resultid="4635" heatid="10250" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4636">
              <RESULTS>
                <RESULT eventid="1162" points="512" swimtime="00:21:55.39" resultid="4637" heatid="10297" lane="6" entrytime="00:22:00.00" />
                <RESULT eventid="1195" points="526" swimtime="00:00:35.74" resultid="4638" heatid="10138" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1228" points="523" swimtime="00:01:07.96" resultid="4639" heatid="10155" lane="3" entrytime="00:01:03.00" />
                <RESULT eventid="1401" points="490" reactiontime="+89" swimtime="00:01:22.52" resultid="4640" heatid="10203" lane="1" entrytime="00:01:17.00" />
                <RESULT eventid="1465" points="423" swimtime="00:02:43.25" resultid="4641" heatid="10220" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="534" swimtime="00:00:30.23" resultid="4642" heatid="10253" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1606" points="408" reactiontime="+94" swimtime="00:03:09.99" resultid="4643" heatid="10265" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-05" firstname="Marcin" gender="M" lastname="Szczypiński" nation="POL" athleteid="4644">
              <RESULTS>
                <RESULT eventid="1077" points="889" swimtime="00:00:26.37" resultid="4645" heatid="10110" lane="7" entrytime="00:00:27.80" />
                <RESULT eventid="1162" points="642" swimtime="00:18:40.29" resultid="4646" heatid="10296" lane="3" entrytime="00:19:00.00" />
                <RESULT eventid="1195" points="719" swimtime="00:00:29.19" resultid="4647" heatid="10140" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1228" points="766" swimtime="00:00:55.26" resultid="4648" heatid="10158" lane="5" entrytime="00:00:56.00" />
                <RESULT eventid="1401" points="686" reactiontime="+76" swimtime="00:01:03.74" resultid="4649" heatid="10205" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1465" points="649" swimtime="00:02:07.78" resultid="4650" heatid="10223" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="832" swimtime="00:00:59.04" resultid="4651" heatid="10240" lane="3" entrytime="00:01:01.50" />
                <RESULT eventid="1686" points="666" swimtime="00:04:36.40" resultid="4652" heatid="10292" lane="5" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="200" swimtime="00:02:16.87" />
                    <SPLIT distance="300" swimtime="00:03:28.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="4653">
              <RESULTS>
                <RESULT eventid="1077" points="711" swimtime="00:00:31.46" resultid="4654" heatid="10107" lane="6" entrytime="00:00:31.70" />
                <RESULT eventid="1292" points="427" swimtime="00:03:22.11" resultid="4655" heatid="10165" lane="1" entrytime="00:03:13.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="587" swimtime="00:01:16.85" resultid="4656" heatid="10238" lane="1" entrytime="00:01:17.45" />
                <RESULT eventid="1574" points="732" swimtime="00:00:28.96" resultid="4657" heatid="10253" lane="8" entrytime="00:00:29.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="4658">
              <RESULTS>
                <RESULT eventid="1141" status="DNF" swimtime="00:00:00.00" resultid="4659" heatid="10295" lane="5" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:46.08" />
                    <SPLIT distance="200" swimtime="00:05:55.58" />
                    <SPLIT distance="300" swimtime="00:09:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="579" swimtime="00:01:06.08" resultid="4660" heatid="10126" lane="6" entrytime="00:01:12.00" />
                <RESULT eventid="1212" points="307" swimtime="00:02:35.38" resultid="4661" heatid="10141" lane="7" entrytime="00:02:30.00" />
                <RESULT eventid="1385" points="547" reactiontime="+85" swimtime="00:02:39.64" resultid="4662" heatid="10193" lane="3" entrytime="00:02:30.00" />
                <RESULT eventid="1558" points="383" swimtime="00:01:01.93" resultid="4663" heatid="10241" lane="7" entrytime="00:01:12.00" />
                <RESULT eventid="1670" points="285" swimtime="00:11:48.54" resultid="4664" heatid="10282" lane="7" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:47.54" />
                    <SPLIT distance="200" swimtime="00:05:48.84" />
                    <SPLIT distance="300" swimtime="00:08:54.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-02-02" firstname="Maria" gender="F" lastname="Śmiglewska" nation="POL" athleteid="4665">
              <RESULTS>
                <RESULT eventid="1178" points="206" swimtime="00:01:21.07" resultid="4666" heatid="10126" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1308" points="207" swimtime="00:07:10.78" resultid="4667" heatid="10167" lane="6" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:03:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="158" swimtime="00:01:27.14" resultid="4668" heatid="10179" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="1385" points="181" reactiontime="+127" swimtime="00:03:09.62" resultid="4669" heatid="10193" lane="2" entrytime="00:02:45.00" />
                <RESULT eventid="1638" points="136" swimtime="00:03:35.26" resultid="4670" heatid="10270" lane="4" entrytime="00:03:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-15" firstname="Andrzej" gender="M" lastname="Porszke" nation="POL" athleteid="4673">
              <RESULTS>
                <RESULT eventid="1369" points="300" swimtime="00:00:43.01" resultid="4674" heatid="10184" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1574" points="140" swimtime="00:00:44.58" resultid="4675" heatid="10249" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1654" status="DSQ" swimtime="00:01:39.66" resultid="4676" heatid="10276" lane="6" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+88" swimtime="00:02:22.61" resultid="4677" heatid="10161" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4636" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="4624" number="2" />
                    <RELAYPOSITION athleteid="4629" number="3" />
                    <RELAYPOSITION athleteid="4653" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:02:03.53" resultid="4678" heatid="10207" lane="4" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4653" number="1" />
                    <RELAYPOSITION athleteid="4624" number="2" />
                    <RELAYPOSITION athleteid="4629" number="3" />
                    <RELAYPOSITION athleteid="4636" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UKFOX" name="UKS Foxball" nation="POL">
          <CONTACT city="Rzeszów" name="Nabożny Maciej" street="ks. Jałowego 22" zip="35-010" />
          <ATHLETES>
            <ATHLETE birthdate="1976-11-13" firstname="Tomasz" gender="M" lastname="Marek" nation="POL" athleteid="4687">
              <RESULTS>
                <RESULT eventid="1077" points="241" swimtime="00:00:40.37" resultid="4688" heatid="10107" lane="1" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT eventid="1228" points="326" swimtime="00:01:14.68" resultid="4689" heatid="10152" lane="2" entrytime="00:01:10.00" entrycourse="LCM" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4690" heatid="10219" lane="4" entrytime="00:02:35.00" entrycourse="LCM" />
                <RESULT eventid="1574" points="349" swimtime="00:00:32.87" resultid="4691" heatid="10251" lane="3" entrytime="00:00:30.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-18" firstname="Mateusz" gender="M" lastname="Szal" nation="POL" athleteid="4692">
              <RESULTS>
                <RESULT eventid="1228" points="366" swimtime="00:01:10.65" resultid="4693" heatid="10153" lane="1" entrytime="00:01:07.00" entrycourse="LCM" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4694" heatid="10219" lane="3" entrytime="00:02:35.00" entrycourse="LCM" />
                <RESULT eventid="1574" points="428" swimtime="00:00:30.17" resultid="4695" heatid="10255" lane="2" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1686" points="267" swimtime="00:06:14.63" resultid="4696" heatid="10290" lane="8" entrytime="00:05:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.29" />
                    <SPLIT distance="200" swimtime="00:02:54.56" />
                    <SPLIT distance="300" swimtime="00:04:34.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASBYD" name="Astoria Bydgoszcz" nation="POL">
          <CONTACT email="sikoreczka7@o2.pl" name="Sikorska" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Kawecki" nation="POL" athleteid="4698">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4699" heatid="10119" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="1162" status="DNS" swimtime="00:00:00.00" resultid="4700" heatid="10298" lane="5" entrytime="00:23:00.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4701" heatid="10152" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="4702" heatid="10174" lane="5" entrytime="00:03:15.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4703" heatid="10202" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4704" heatid="10230" lane="8" entrytime="00:06:20.00" />
                <RESULT eventid="1606" status="DNS" swimtime="00:00:00.00" resultid="4705" heatid="10264" lane="5" entrytime="00:02:58.00" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="4706" heatid="10279" lane="3" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" name="TS Olimpia Poznań" nation="POL" region="WIE" shortname="Olimpia Poznań">
          <CONTACT email="zpietraszewski@empi2.pl" name="Pietraszewski Zbigniew" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="4995">
              <RESULTS>
                <RESULT eventid="1093" points="678" swimtime="00:03:16.30" resultid="4996" heatid="10112" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="690" swimtime="00:00:41.92" resultid="4997" heatid="10128" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1308" points="747" swimtime="00:03:29.24" resultid="4998" heatid="10168" lane="3" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1352" points="710" swimtime="00:00:43.11" resultid="4999" heatid="10181" lane="7" entrytime="00:00:44.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1385" points="752" reactiontime="+84" swimtime="00:01:30.13" resultid="5000" heatid="10196" lane="1" entrytime="00:01:30.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1590" points="880" reactiontime="+93" swimtime="00:03:13.59" resultid="5001" heatid="10259" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="712" swimtime="00:01:37.74" resultid="5002" heatid="10272" lane="2" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="5003">
              <RESULTS>
                <RESULT eventid="1212" points="461" swimtime="00:01:32.41" resultid="5004" heatid="10142" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="1352" points="431" swimtime="00:00:51.07" resultid="5005" heatid="10180" lane="8" entrytime="00:00:54.00" />
                <RESULT eventid="1481" points="454" swimtime="00:08:19.43" resultid="5006" heatid="10224" lane="3" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:09.71" />
                    <SPLIT distance="200" swimtime="00:04:19.70" />
                    <SPLIT distance="300" swimtime="00:06:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="611" swimtime="00:00:37.87" resultid="5007" heatid="10242" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1638" points="309" swimtime="00:02:07.80" resultid="5008" heatid="10271" lane="5" entrytime="00:01:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="5009">
              <RESULTS>
                <RESULT eventid="1686" status="DNS" swimtime="00:00:00.00" resultid="5012" heatid="10286" lane="4" entrytime="00:07:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="5013">
              <RESULTS>
                <RESULT eventid="1109" points="545" swimtime="00:03:09.46" resultid="5014" heatid="10118" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="564" swimtime="00:06:48.88" resultid="5017" heatid="10229" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.11" />
                    <SPLIT distance="200" swimtime="00:03:26.22" />
                    <SPLIT distance="300" swimtime="00:05:17.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="503" reactiontime="+91" swimtime="00:03:09.34" resultid="5018" heatid="10264" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="421" swimtime="00:00:42.55" resultid="10302" heatid="10136" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1401" points="421" reactiontime="+89" swimtime="00:01:30.15" resultid="10303" heatid="10200" lane="4" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOPO" name="TP Masters Opole" nation="POL" shortname="Masters Opole">
          <CONTACT email="OPOLBUD@ONET.EU" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="TADEUSZ" gender="M" lastname="WITKOWSKI" nation="POL" athleteid="5045">
              <RESULTS>
                <RESULT eventid="1195" points="470" swimtime="00:00:50.83" resultid="5046" heatid="10134" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1228" points="476" swimtime="00:01:34.78" resultid="5047" heatid="10148" lane="8" entrytime="00:01:36.00" />
                <RESULT eventid="1369" points="355" swimtime="00:00:56.60" resultid="5048" heatid="10184" lane="2" entrytime="00:00:51.00" />
                <RESULT eventid="1401" points="393" reactiontime="+70" swimtime="00:02:00.19" resultid="5049" heatid="10199" lane="6" entrytime="00:01:52.00" />
                <RESULT eventid="1574" points="812" swimtime="00:00:35.14" resultid="5050" heatid="10249" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1606" points="377" reactiontime="+102" swimtime="00:04:20.00" resultid="5051" heatid="10262" lane="2" entrytime="00:04:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEOSI" name="Dęby Osielsko" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1990-09-12" firstname="Adrian" gender="M" lastname="Teodorski" nation="POL" athleteid="5618">
              <RESULTS>
                <RESULT eventid="1077" points="656" swimtime="00:00:28.54" resultid="5620" heatid="10110" lane="3" entrytime="00:00:26.90" />
                <RESULT eventid="1109" points="423" swimtime="00:02:44.47" resultid="5621" heatid="10122" lane="5" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="534" swimtime="00:01:00.84" resultid="5622" heatid="10158" lane="3" entrytime="00:00:56.80" />
                <RESULT eventid="1292" points="379" swimtime="00:02:45.81" resultid="5623" heatid="10166" lane="7" entrytime="00:02:32.15">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="462" swimtime="00:02:19.29" resultid="5624" heatid="10223" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="343" swimtime="00:06:16.99" resultid="5625" heatid="10231" lane="7" entrytime="00:05:24.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="200" swimtime="00:02:58.03" />
                    <SPLIT distance="300" swimtime="00:04:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="584" swimtime="00:01:04.19" resultid="5626" heatid="10240" lane="6" entrytime="00:01:01.50" />
                <RESULT eventid="1574" points="547" swimtime="00:00:27.29" resultid="5627" heatid="10257" lane="5" entrytime="00:00:25.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOLS" name="AZS UWM Masters Olsztyn" nation="POL" shortname="Masters Olsztyn">
          <CONTACT city="Łupstych" email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" phone="501372846" state="WARM-" street="Leśna 1" zip="11-041" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="5629">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1077" points="774" swimtime="00:00:30.58" resultid="5630" heatid="10108" lane="8" entrytime="00:00:31.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1162" points="898" swimtime="00:20:20.71" resultid="5631" heatid="10296" lane="6" entrytime="00:19:50.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1195" points="824" swimtime="00:00:34.03" resultid="5632" heatid="10139" lane="7" entrytime="00:00:34.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1292" points="757" swimtime="00:02:47.03" resultid="5633" heatid="10165" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="724" reactiontime="+87" swimtime="00:01:15.25" resultid="5634" heatid="10204" lane="6" entrytime="00:01:12.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1542" points="757" swimtime="00:01:10.62" resultid="5635" heatid="10239" lane="6" entrytime="00:01:10.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1686" points="872" swimtime="00:04:59.65" resultid="5636" heatid="10292" lane="1" entrytime="00:04:54.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="200" swimtime="00:02:28.07" />
                    <SPLIT distance="300" swimtime="00:03:44.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="5637">
              <RESULTS>
                <RESULT eventid="1061" points="283" swimtime="00:00:43.89" resultid="5638" heatid="10098" lane="1" entrytime="00:00:40.05" />
                <RESULT eventid="1141" points="382" swimtime="00:12:58.85" resultid="5639" heatid="10293" lane="8" entrytime="00:12:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.86" />
                    <SPLIT distance="200" swimtime="00:04:42.14" />
                    <SPLIT distance="300" swimtime="00:06:21.09" />
                    <SPLIT distance="400" swimtime="00:08:00.94" />
                    <SPLIT distance="500" swimtime="00:09:41.56" />
                    <SPLIT distance="600" swimtime="00:11:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="385" swimtime="00:01:19.76" resultid="5640" heatid="10143" lane="4" entrytime="00:01:19.00" />
                <RESULT eventid="1449" points="367" swimtime="00:02:54.93" resultid="5641" heatid="10212" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="292" swimtime="00:01:36.32" resultid="5642" heatid="10232" lane="4" entrytime="00:01:35.00" />
                <RESULT eventid="1670" points="367" swimtime="00:06:14.37" resultid="5643" heatid="10284" lane="2" entrytime="00:06:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="200" swimtime="00:03:04.32" />
                    <SPLIT distance="300" swimtime="00:04:41.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="5644">
              <RESULTS>
                <RESULT eventid="1077" points="648" swimtime="00:00:29.04" resultid="5645" heatid="10102" lane="4" entrytime="00:00:41.50" />
                <RESULT eventid="1109" points="510" swimtime="00:02:36.97" resultid="5646" heatid="10121" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="635" swimtime="00:00:59.81" resultid="5647" heatid="10156" lane="5" entrytime="00:01:01.00" />
                <RESULT eventid="1369" points="525" swimtime="00:00:35.71" resultid="5648" heatid="10190" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1574" points="620" swimtime="00:00:27.14" resultid="5649" heatid="10255" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1686" points="519" swimtime="00:05:05.24" resultid="5650" heatid="10291" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="200" swimtime="00:02:30.30" />
                    <SPLIT distance="300" swimtime="00:03:47.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="5651">
              <RESULTS>
                <RESULT eventid="1141" points="581" swimtime="00:12:18.65" resultid="5652" heatid="10293" lane="7" entrytime="00:12:15.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.00" />
                    <SPLIT distance="200" swimtime="00:02:59.50" />
                    <SPLIT distance="300" swimtime="00:04:33.42" />
                    <SPLIT distance="400" swimtime="00:06:07.25" />
                    <SPLIT distance="500" swimtime="00:07:41.08" />
                    <SPLIT distance="600" swimtime="00:09:14.46" />
                    <SPLIT distance="700" swimtime="00:10:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="577" swimtime="00:01:16.31" resultid="5653" heatid="10144" lane="2" entrytime="00:01:16.50" />
                <RESULT eventid="1308" points="525" swimtime="00:03:32.10" resultid="5654" heatid="10168" lane="2" entrytime="00:03:30.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="575" swimtime="00:06:53.18" resultid="5655" heatid="10225" lane="2" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.33" />
                    <SPLIT distance="200" swimtime="00:03:32.01" />
                    <SPLIT distance="300" swimtime="00:05:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="531" swimtime="00:00:34.76" resultid="5656" heatid="10244" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="1670" points="518" swimtime="00:06:04.64" resultid="5657" heatid="10284" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="200" swimtime="00:03:00.75" />
                    <SPLIT distance="300" swimtime="00:04:34.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="5658">
              <RESULTS>
                <RESULT eventid="1109" points="489" swimtime="00:02:43.34" resultid="5659" heatid="10121" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="455" swimtime="00:00:33.94" resultid="5660" heatid="10139" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1324" points="538" swimtime="00:02:52.76" resultid="5661" heatid="10177" lane="2" entrytime="00:02:47.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="625" swimtime="00:00:34.45" resultid="5662" heatid="10191" lane="6" entrytime="00:00:34.80" />
                <RESULT eventid="1401" points="415" reactiontime="+74" swimtime="00:01:15.92" resultid="5663" heatid="10204" lane="8" entrytime="00:01:15.00" />
                <RESULT eventid="1654" points="558" swimtime="00:01:18.77" resultid="5664" heatid="10281" lane="7" entrytime="00:01:16.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:10.86" resultid="5665" heatid="10123" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5651" number="1" />
                    <RELAYPOSITION athleteid="5637" number="2" />
                    <RELAYPOSITION athleteid="5629" number="3" />
                    <RELAYPOSITION athleteid="5644" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+88" swimtime="00:02:32.39" resultid="5666" heatid="10267" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5629" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5658" number="2" />
                    <RELAYPOSITION athleteid="5637" number="3" />
                    <RELAYPOSITION athleteid="5651" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAKRO" name="Master Krosno" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1966-04-10" firstname="Bogdan" gender="M" lastname="Żebracki" nation="POL" athleteid="5672">
              <RESULTS>
                <RESULT eventid="1162" points="409" swimtime="00:23:38.04" resultid="5674" heatid="10298" lane="2" entrytime="00:23:35.00" />
                <RESULT eventid="1195" points="495" swimtime="00:00:36.48" resultid="5675" heatid="10138" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1324" points="516" swimtime="00:03:11.91" resultid="5677" heatid="10175" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="429" swimtime="00:00:40.73" resultid="5678" heatid="10189" lane="1" entrytime="00:00:38.70" />
                <RESULT eventid="1401" points="501" reactiontime="+97" swimtime="00:01:21.89" resultid="5679" heatid="10202" lane="6" entrytime="00:01:21.00" />
                <RESULT eventid="1606" points="390" reactiontime="+104" swimtime="00:03:12.76" resultid="5681" heatid="10264" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="485" swimtime="00:01:27.48" resultid="5688" heatid="10278" lane="4" entrytime="00:01:26.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" name="MKP BOBRY Dębica" nation="POL" shortname="BOBRY Dębica">
          <CONTACT name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1967-11-09" firstname="Elżbieta" gender="F" lastname="Nowak-Bereś" nation="POL" athleteid="5030">
              <RESULTS>
                <RESULT eventid="1061" points="244" swimtime="00:00:48.77" resultid="5031" heatid="10096" lane="4" entrytime="00:00:48.98" />
                <RESULT eventid="1352" points="418" swimtime="00:00:48.25" resultid="5032" heatid="10180" lane="7" entrytime="00:00:51.95" />
                <RESULT eventid="1558" points="241" swimtime="00:00:45.21" resultid="5033" heatid="10241" lane="4" entrytime="00:00:46.05" />
                <RESULT eventid="1638" status="DSQ" swimtime="00:01:59.53" resultid="5034" heatid="10271" lane="3" entrytime="00:01:57.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-04" firstname="Zenon" gender="M" lastname="Dul" nation="POL" athleteid="5682">
              <RESULTS>
                <RESULT eventid="1077" points="258" swimtime="00:00:44.09" resultid="5684" heatid="10102" lane="6" entrytime="00:00:42.51" />
                <RESULT eventid="1369" points="252" swimtime="00:00:52.51" resultid="5685" heatid="10185" lane="3" entrytime="00:00:47.22" />
                <RESULT eventid="1324" points="216" swimtime="00:04:34.31" resultid="5686" heatid="10170" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="315" swimtime="00:00:38.36" resultid="5687" heatid="10248" lane="6" entrytime="00:00:36.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-25" firstname="Stanisław" gender="M" lastname="Skop" nation="POL" athleteid="7955">
              <RESULTS>
                <RESULT eventid="1109" points="375" swimtime="00:02:51.16" resultid="7956" heatid="10119" lane="7" entrytime="00:02:59.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="355" swimtime="00:00:35.94" resultid="7957" heatid="10139" lane="2" entrytime="00:00:33.87" />
                <RESULT eventid="1324" points="430" swimtime="00:02:58.64" resultid="7958" heatid="10175" lane="4" entrytime="00:03:05.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="623" swimtime="00:00:33.16" resultid="7959" heatid="10192" lane="7" entrytime="00:00:33.26" />
                <RESULT eventid="1574" status="DNS" swimtime="00:00:00.00" resultid="7960" heatid="10253" lane="3" entrytime="00:00:28.55" />
                <RESULT eventid="1654" points="475" swimtime="00:01:19.61" resultid="7961" heatid="10281" lane="1" entrytime="00:01:17.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-15" firstname="Tomasz" gender="M" lastname="Dąbrowski" nation="POL" athleteid="8071" />
            <ATHLETE birthdate="1987-07-07" firstname="Olga" gender="F" lastname="Siembab" nation="POL" athleteid="8177">
              <RESULTS>
                <RESULT eventid="1141" points="256" swimtime="00:14:33.85" resultid="8178" heatid="10293" lane="1" entrytime="00:12:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.07" />
                    <SPLIT distance="200" swimtime="00:03:18.04" />
                    <SPLIT distance="300" swimtime="00:05:12.77" />
                    <SPLIT distance="400" swimtime="00:07:07.51" />
                    <SPLIT distance="500" swimtime="00:09:01.00" />
                    <SPLIT distance="600" swimtime="00:10:52.50" />
                    <SPLIT distance="700" swimtime="00:12:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="303" swimtime="00:00:45.33" resultid="8179" heatid="10128" lane="6" entrytime="00:00:42.30" />
                <RESULT eventid="1385" points="257" reactiontime="+86" swimtime="00:01:39.74" resultid="8180" heatid="10195" lane="4" entrytime="00:01:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" athleteid="8181">
              <RESULTS>
                <RESULT eventid="1077" points="520" swimtime="00:00:31.25" resultid="8182" heatid="10107" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1162" points="455" swimtime="00:21:19.39" resultid="8183" heatid="10297" lane="4" entrytime="00:20:30.00" />
                <RESULT eventid="1574" points="542" swimtime="00:00:28.38" resultid="8185" heatid="10255" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1686" points="477" swimtime="00:05:14.10" resultid="8186" heatid="10291" lane="8" entrytime="00:05:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="200" swimtime="00:02:33.69" />
                    <SPLIT distance="300" swimtime="00:03:54.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:22.71" resultid="8140" heatid="10124" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5030" number="1" />
                    <RELAYPOSITION athleteid="8071" number="2" />
                    <RELAYPOSITION athleteid="8177" number="3" />
                    <RELAYPOSITION athleteid="8181" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+84" swimtime="00:02:38.48" resultid="8141" heatid="10268" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8177" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="5030" number="2" />
                    <RELAYPOSITION athleteid="8181" number="3" />
                    <RELAYPOSITION athleteid="8071" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00608" name="Wodnik MOSiR Krosno" nation="POL" region="PDK" shortname="Wodnik Krosno">
          <CONTACT city="Krosno" name="Wodnik MOSiR Krosno" phone="013 43 20480" state="PODKA" street="Bursaki 41" zip="38-400" />
        </CLUB>
        <CLUB type="CLUB" code="KOKRA" name="Masters Korona Kraków" nation="POL" region="KR" shortname="Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" street="Kalwaryjska" />
          <ATHLETES>
            <ATHLETE birthdate="1933-04-07" firstname="Tadeusz" gender="M" lastname="Banach" nation="POL" athleteid="5705">
              <RESULTS>
                <RESULT eventid="1195" points="102" swimtime="00:01:27.58" resultid="5706" heatid="10132" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1574" points="77" swimtime="00:01:17.84" resultid="5707" heatid="10246" lane="5" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-04-24" firstname="Krzysztof" gender="M" lastname="Chołda" nation="POL" athleteid="5708">
              <RESULTS>
                <RESULT eventid="1162" points="406" swimtime="00:23:41.10" resultid="5709" heatid="10298" lane="3" entrytime="00:23:25.00" />
                <RESULT eventid="1228" points="481" swimtime="00:01:09.88" resultid="5710" heatid="10149" lane="4" entrytime="00:01:16.00" />
                <RESULT eventid="1369" points="425" swimtime="00:00:40.83" resultid="5711" heatid="10187" lane="6" entrytime="00:00:42.25" />
                <RESULT eventid="1574" points="408" swimtime="00:00:33.06" resultid="5712" heatid="10251" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1654" points="383" swimtime="00:01:34.61" resultid="5713" heatid="10277" lane="2" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="Data" nation="POL" athleteid="5714">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="5715" heatid="10149" lane="5" entrytime="00:01:18.00" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="5716" heatid="10173" lane="7" entrytime="00:03:35.00" />
                <RESULT eventid="1369" points="359" swimtime="00:00:45.27" resultid="5717" heatid="10185" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1465" points="322" swimtime="00:03:01.27" resultid="5718" heatid="10217" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="391" swimtime="00:01:39.44" resultid="5719" heatid="10277" lane="7" entrytime="00:01:37.00" />
                <RESULT eventid="1686" points="317" swimtime="00:06:33.52" resultid="5720" heatid="10288" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.33" />
                    <SPLIT distance="200" swimtime="00:03:06.17" />
                    <SPLIT distance="300" swimtime="00:04:52.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-07" firstname="Robert" gender="M" lastname="Grela" nation="POL" athleteid="5721">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:31.33" resultid="5722" heatid="10109" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1292" points="586" swimtime="00:02:49.45" resultid="5723" heatid="10166" lane="8" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="519" reactiontime="+78" swimtime="00:01:20.94" resultid="5724" heatid="10203" lane="6" entrytime="00:01:16.00" />
                <RESULT eventid="1542" points="665" swimtime="00:01:10.27" resultid="5725" heatid="10239" lane="5" entrytime="00:01:07.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Wojciech" gender="M" lastname="Hoffman" nation="POL" athleteid="5726">
              <RESULTS>
                <RESULT eventid="1162" points="427" swimtime="00:21:46.60" resultid="5727" heatid="10296" lane="7" entrytime="00:20:00.00" />
                <RESULT eventid="1228" points="438" swimtime="00:01:07.71" resultid="5728" heatid="10154" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1465" points="465" swimtime="00:02:29.91" resultid="5729" heatid="10220" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="427" swimtime="00:00:30.74" resultid="5730" heatid="10252" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1686" points="421" swimtime="00:05:27.42" resultid="5731" heatid="10290" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="200" swimtime="00:02:39.17" />
                    <SPLIT distance="300" swimtime="00:04:04.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="5732">
              <RESULTS>
                <RESULT eventid="1061" points="426" swimtime="00:00:39.39" resultid="5733" heatid="10098" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1093" points="335" swimtime="00:03:32.69" resultid="5734" heatid="10111" lane="6" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="400" swimtime="00:00:42.65" resultid="5735" heatid="10128" lane="2" entrytime="00:00:42.70" />
                <RESULT eventid="1385" points="377" reactiontime="+99" swimtime="00:01:32.31" resultid="5736" heatid="10195" lane="1" entrytime="00:01:38.00" />
                <RESULT eventid="1481" points="334" swimtime="00:07:38.50" resultid="5737" heatid="10225" lane="7" entrytime="00:07:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:03:51.11" />
                    <SPLIT distance="300" swimtime="00:05:59.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="364" reactiontime="+101" swimtime="00:03:23.58" resultid="5738" heatid="10259" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="307" swimtime="00:06:43.14" resultid="5739" heatid="10283" lane="2" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.00" />
                    <SPLIT distance="200" swimtime="00:03:16.70" />
                    <SPLIT distance="300" swimtime="00:05:02.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-15" firstname="Monika" gender="F" lastname="Jaworska" nation="POL" athleteid="5740">
              <RESULTS>
                <RESULT eventid="1061" points="522" swimtime="00:00:34.27" resultid="5741" heatid="10099" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1093" points="376" swimtime="00:03:12.40" resultid="5742" heatid="10112" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="373" swimtime="00:01:17.52" resultid="5743" heatid="10145" lane="8" entrytime="00:01:12.00" />
                <RESULT eventid="1352" points="321" swimtime="00:00:47.90" resultid="5744" heatid="10181" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1525" points="342" swimtime="00:01:27.68" resultid="5745" heatid="10233" lane="6" entrytime="00:01:23.00" />
                <RESULT eventid="1558" points="383" swimtime="00:00:35.26" resultid="5746" heatid="10245" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-20" firstname="Joanna" gender="F" lastname="Kieszek" nation="POL" athleteid="5747">
              <RESULTS>
                <RESULT eventid="1061" points="479" swimtime="00:00:35.27" resultid="5748" heatid="10099" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1212" points="550" swimtime="00:01:08.11" resultid="5749" heatid="10146" lane="2" entrytime="00:01:07.00" />
                <RESULT eventid="1449" points="489" swimtime="00:02:37.39" resultid="5750" heatid="10213" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="596" swimtime="00:00:30.42" resultid="5751" heatid="10245" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1093" points="386" swimtime="00:03:10.80" resultid="7713" heatid="10113" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="401" swimtime="00:00:44.46" resultid="7714" heatid="10181" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1670" points="348" swimtime="00:06:00.43" resultid="7715" heatid="10285" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.61" />
                    <SPLIT distance="200" swimtime="00:02:52.41" />
                    <SPLIT distance="300" swimtime="00:04:26.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="5752">
              <RESULTS>
                <RESULT eventid="1401" points="148" reactiontime="+61" swimtime="00:02:39.78" resultid="5756" heatid="10198" lane="6" entrytime="00:02:30.00" />
                <RESULT eventid="1465" points="207" swimtime="00:04:21.40" resultid="5757" heatid="10215" lane="6" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="251" swimtime="00:00:47.78" resultid="5758" heatid="10247" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1606" points="163" reactiontime="+79" swimtime="00:05:39.07" resultid="5759" heatid="10261" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:48.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="143" swimtime="00:05:55.21" resultid="5753" heatid="10114" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="184" swimtime="00:01:07.19" resultid="5754" heatid="10132" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1228" points="235" swimtime="00:01:48.54" resultid="5755" heatid="10147" lane="5" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="5760">
              <RESULTS>
                <RESULT eventid="1178" points="702" swimtime="00:00:37.54" resultid="5761" heatid="10127" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="600" swimtime="00:01:15.31" resultid="5762" heatid="10145" lane="1" entrytime="00:01:12.00" />
                <RESULT eventid="1352" points="692" swimtime="00:00:40.79" resultid="5763" heatid="10180" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1558" points="635" swimtime="00:00:32.76" resultid="5764" heatid="10244" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="5765">
              <RESULTS>
                <RESULT eventid="1093" points="335" swimtime="00:03:24.24" resultid="5766" heatid="10111" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="502" swimtime="00:03:18.54" resultid="5767" heatid="10168" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="491" swimtime="00:00:43.21" resultid="5768" heatid="10181" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1638" points="416" swimtime="00:01:34.65" resultid="5769" heatid="10272" lane="3" entrytime="00:01:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="5770">
              <RESULTS>
                <RESULT eventid="1077" points="548" swimtime="00:00:30.99" resultid="5771" heatid="10108" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1228" points="604" swimtime="00:00:59.83" resultid="5772" heatid="10157" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1465" points="475" swimtime="00:02:21.81" resultid="5773" heatid="10222" lane="6" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="646" swimtime="00:00:26.30" resultid="5774" heatid="10256" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1686" points="434" swimtime="00:05:18.75" resultid="5775" heatid="10290" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="200" swimtime="00:02:37.30" />
                    <SPLIT distance="300" swimtime="00:03:58.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="5776">
              <RESULTS>
                <RESULT eventid="1061" points="463" swimtime="00:00:43.37" resultid="5777" heatid="10095" lane="3" />
                <RESULT eventid="1093" points="520" swimtime="00:03:34.41" resultid="5778" heatid="10111" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="588" swimtime="00:00:44.22" resultid="5779" heatid="10128" lane="8" entrytime="00:00:43.67" />
                <RESULT eventid="1276" points="471" swimtime="00:03:58.94" resultid="5780" heatid="10162" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="530" reactiontime="+100" swimtime="00:01:41.28" resultid="5781" heatid="10195" lane="3" entrytime="00:01:33.45" />
                <RESULT eventid="1481" points="491" swimtime="00:07:48.50" resultid="5782" heatid="10224" lane="4" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.78" />
                    <SPLIT distance="200" swimtime="00:03:56.66" />
                    <SPLIT distance="300" swimtime="00:06:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="638" swimtime="00:00:36.03" resultid="5783" heatid="10243" lane="4" entrytime="00:00:35.54" />
                <RESULT eventid="1670" points="488" swimtime="00:07:03.37" resultid="5784" heatid="10284" lane="1" entrytime="00:06:30.54">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.93" />
                    <SPLIT distance="200" swimtime="00:03:26.63" />
                    <SPLIT distance="300" swimtime="00:05:16.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="5785">
              <RESULTS>
                <RESULT eventid="1061" points="568" swimtime="00:00:39.81" resultid="5786" heatid="10095" lane="5" />
                <RESULT eventid="1141" points="465" swimtime="00:13:33.44" resultid="5787" heatid="10295" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="200" swimtime="00:03:11.60" />
                    <SPLIT distance="300" swimtime="00:04:56.05" />
                    <SPLIT distance="400" swimtime="00:06:40.96" />
                    <SPLIT distance="500" swimtime="00:08:25.97" />
                    <SPLIT distance="600" swimtime="00:10:10.63" />
                    <SPLIT distance="700" swimtime="00:11:55.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="5803">
              <RESULTS>
                <RESULT eventid="1061" points="122" swimtime="00:01:19.08" resultid="5804" heatid="10096" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1093" points="211" swimtime="00:05:30.57" resultid="5805" heatid="10111" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="207" swimtime="00:02:10.03" resultid="5806" heatid="10141" lane="2" entrytime="00:02:06.00" />
                <RESULT eventid="1308" points="257" swimtime="00:05:40.21" resultid="5807" heatid="10167" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1385" points="193" reactiontime="+65" swimtime="00:02:39.98" resultid="5808" heatid="10193" lane="5" entrytime="00:02:28.00" />
                <RESULT eventid="1449" points="155" swimtime="00:05:15.41" resultid="5809" heatid="10209" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:19.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="263" swimtime="00:02:31.66" resultid="5810" heatid="10271" lane="2" entrytime="00:02:15.00" />
                <RESULT eventid="1670" points="132" swimtime="00:11:35.68" resultid="5811" heatid="10282" lane="2" entrytime="00:09:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:45.06" />
                    <SPLIT distance="200" swimtime="00:05:47.04" />
                    <SPLIT distance="300" swimtime="00:08:49.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="5812">
              <RESULTS>
                <RESULT eventid="1093" points="545" swimtime="00:02:53.75" resultid="5813" heatid="10112" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="611" swimtime="00:00:35.87" resultid="5814" heatid="10130" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1212" points="510" swimtime="00:01:11.89" resultid="5815" heatid="10145" lane="2" entrytime="00:01:10.00" />
                <RESULT eventid="1385" points="548" reactiontime="+72" swimtime="00:01:17.54" resultid="5816" heatid="10197" lane="6" entrytime="00:01:17.00" />
                <RESULT eventid="1590" points="494" reactiontime="+73" swimtime="00:02:50.89" resultid="5817" heatid="10260" lane="7" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="446" swimtime="00:05:48.02" resultid="5818" heatid="10284" lane="6" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.81" />
                    <SPLIT distance="200" swimtime="00:02:52.10" />
                    <SPLIT distance="300" swimtime="00:04:23.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="5819">
              <RESULTS>
                <RESULT eventid="1077" points="764" swimtime="00:00:30.33" resultid="5820" heatid="10106" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1195" points="607" swimtime="00:00:36.16" resultid="5821" heatid="10137" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="5822" heatid="10152" lane="5" entrytime="00:01:08.00" />
                <RESULT eventid="1369" points="584" swimtime="00:00:38.51" resultid="5823" heatid="10187" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1401" points="563" reactiontime="+95" swimtime="00:01:21.36" resultid="5824" heatid="10203" lane="8" entrytime="00:01:19.00" />
                <RESULT eventid="1542" status="DSQ" swimtime="00:01:22.74" resultid="5825" heatid="10238" lane="5" entrytime="00:01:16.00" />
                <RESULT eventid="1606" status="DNS" swimtime="00:00:00.00" resultid="5826" heatid="10264" lane="2" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="5827">
              <RESULTS>
                <RESULT eventid="1195" points="141" swimtime="00:00:52.70" resultid="5828" heatid="10133" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1401" points="119" reactiontime="+86" swimtime="00:01:59.47" resultid="5829" heatid="10199" lane="8" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="5830">
              <RESULTS>
                <RESULT eventid="1061" points="537" swimtime="00:00:37.51" resultid="5831" heatid="10099" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="5832">
              <RESULTS>
                <RESULT eventid="1308" points="723" swimtime="00:03:18.79" resultid="5833" heatid="10169" lane="8" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" status="DSQ" swimtime="00:00:42.05" resultid="5834" heatid="10181" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1638" points="730" swimtime="00:01:32.54" resultid="5835" heatid="10273" lane="8" entrytime="00:01:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="5836">
              <RESULTS>
                <RESULT eventid="1162" points="333" swimtime="00:25:17.62" resultid="5837" heatid="10299" lane="5" entrytime="00:25:00.00" />
                <RESULT eventid="1228" points="402" swimtime="00:01:14.20" resultid="5838" heatid="10150" lane="8" entrytime="00:01:16.00" />
                <RESULT eventid="1324" points="278" swimtime="00:03:55.75" resultid="5839" heatid="10172" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="413" swimtime="00:02:44.51" resultid="5840" heatid="10217" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="358" swimtime="00:00:34.54" resultid="5841" heatid="10250" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1686" points="384" swimtime="00:06:01.44" resultid="5842" heatid="10289" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.74" />
                    <SPLIT distance="200" swimtime="00:02:55.94" />
                    <SPLIT distance="300" swimtime="00:04:31.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-17" firstname="Kinga" gender="F" lastname="Sowa" nation="POL" athleteid="5843">
              <RESULTS>
                <RESULT eventid="1178" points="628" swimtime="00:00:34.77" resultid="5844" heatid="10129" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1212" points="550" swimtime="00:01:08.13" resultid="5845" heatid="10145" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1385" points="614" reactiontime="+76" swimtime="00:01:15.35" resultid="5846" heatid="10196" lane="4" entrytime="00:01:22.00" />
                <RESULT eventid="1558" points="624" swimtime="00:00:29.96" resultid="5847" heatid="10245" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-05" firstname="Aleksandra" gender="F" lastname="Jamrozik" nation="POL" athleteid="5848">
              <RESULTS>
                <RESULT eventid="1093" points="581" swimtime="00:02:46.42" resultid="5849" heatid="10113" lane="3" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="532" swimtime="00:00:36.76" resultid="5850" heatid="10130" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1212" points="478" swimtime="00:01:11.35" resultid="5851" heatid="10146" lane="1" entrytime="00:01:08.00" />
                <RESULT eventid="1385" points="520" reactiontime="+76" swimtime="00:01:19.67" resultid="5852" heatid="10197" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1449" points="511" swimtime="00:02:35.15" resultid="5853" heatid="10213" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="484" reactiontime="+75" swimtime="00:02:52.68" resultid="5854" heatid="10260" lane="5" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1670" points="442" swimtime="00:05:32.85" resultid="5855" heatid="10285" lane="7" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.12" />
                    <SPLIT distance="200" swimtime="00:02:41.44" />
                    <SPLIT distance="300" swimtime="00:04:07.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-15" firstname="Klara" gender="F" lastname="Laudańska" nation="POL" athleteid="5856">
              <RESULTS>
                <RESULT eventid="1061" points="177" swimtime="00:00:52.81" resultid="5857" heatid="10096" lane="7" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="5858">
              <RESULTS>
                <RESULT eventid="1077" points="427" swimtime="00:00:35.39" resultid="5859" heatid="10108" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1162" points="541" swimtime="00:20:52.69" resultid="5860" heatid="10296" lane="8" entrytime="00:20:20.00" />
                <RESULT eventid="1292" points="563" swimtime="00:02:37.96" resultid="5861" heatid="10166" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="598" swimtime="00:05:48.19" resultid="5862" heatid="10230" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="200" swimtime="00:02:49.10" />
                    <SPLIT distance="300" swimtime="00:04:29.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-10-10" firstname="Marcin" gender="M" lastname="Wasylewski" nation="POL" athleteid="5863">
              <RESULTS>
                <RESULT eventid="1077" points="253" swimtime="00:00:42.15" resultid="5864" heatid="10102" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-01" firstname="Konrad" gender="M" lastname="Latuszek" nation="POL" athleteid="5865">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5866" heatid="10120" lane="7" entrytime="00:02:45.00" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="5867" heatid="10176" lane="7" entrytime="00:03:05.00" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="5868" heatid="10190" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1654" status="DNS" swimtime="00:00:00.00" resultid="5869" heatid="10280" lane="3" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-01" firstname="Karolina" gender="F" lastname="Zadrożna" nation="POL" athleteid="5870">
              <RESULTS>
                <RESULT eventid="1141" points="513" swimtime="00:10:55.25" resultid="5871" heatid="10293" lane="5" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="200" swimtime="00:02:34.26" />
                    <SPLIT distance="300" swimtime="00:03:56.94" />
                    <SPLIT distance="400" swimtime="00:05:20.96" />
                    <SPLIT distance="500" swimtime="00:06:45.71" />
                    <SPLIT distance="600" swimtime="00:08:09.50" />
                    <SPLIT distance="700" swimtime="00:09:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="544" swimtime="00:01:08.37" resultid="5872" heatid="10141" lane="1" />
                <RESULT eventid="1276" points="251" swimtime="00:03:35.00" resultid="5873" heatid="10162" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="308" swimtime="00:00:48.54" resultid="5874" heatid="10178" lane="3" />
                <RESULT eventid="1449" points="581" swimtime="00:02:28.60" resultid="5875" heatid="10213" lane="3" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1525" points="336" swimtime="00:01:28.23" resultid="5876" heatid="10232" lane="7" />
                <RESULT eventid="1670" points="520" swimtime="00:05:15.32" resultid="5877" heatid="10285" lane="4" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="200" swimtime="00:02:35.34" />
                    <SPLIT distance="300" swimtime="00:03:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-03" firstname="Patrycja" gender="F" lastname="Urbaniak" nation="POL" athleteid="5878">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="5879" heatid="10146" lane="7" entrytime="00:01:07.00" />
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="5880" heatid="10233" lane="4" entrytime="00:01:16.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="5881">
              <RESULTS>
                <RESULT eventid="1178" points="168" swimtime="00:00:56.94" resultid="5882" heatid="10127" lane="8" entrytime="00:00:57.00" />
                <RESULT eventid="1308" points="174" swimtime="00:04:52.26" resultid="5883" heatid="10167" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:20.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="195" swimtime="00:00:58.58" resultid="5884" heatid="10179" lane="6" entrytime="00:00:59.71" />
                <RESULT eventid="1385" points="137" reactiontime="+88" swimtime="00:02:09.06" resultid="5885" heatid="10194" lane="8" entrytime="00:02:07.00" />
                <RESULT eventid="1590" points="142" reactiontime="+111" swimtime="00:04:38.54" resultid="5886" heatid="10258" lane="2" entrytime="00:04:45.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1638" points="166" swimtime="00:02:16.66" resultid="5887" heatid="10271" lane="6" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Robert" gender="M" lastname="Trzos" nation="POL" athleteid="5958">
              <RESULTS>
                <RESULT eventid="1324" points="447" swimtime="00:03:05.42" resultid="5959" heatid="10176" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="7716">
              <RESULTS>
                <RESULT eventid="1109" points="461" swimtime="00:03:43.87" resultid="7717" heatid="10116" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="445" swimtime="00:28:07.47" resultid="7718" heatid="10299" lane="8" entrytime="00:26:15.00" />
                <RESULT eventid="1228" points="632" swimtime="00:01:16.93" resultid="7719" heatid="10150" lane="5" entrytime="00:01:14.00" />
                <RESULT eventid="1292" status="DSQ" swimtime="00:04:56.21" resultid="7720" heatid="10164" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:06.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="479" swimtime="00:03:09.98" resultid="7721" heatid="10217" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="348" swimtime="00:08:51.33" resultid="7722" heatid="10227" lane="4" entrytime="00:07:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:08.01" />
                    <SPLIT distance="200" swimtime="00:04:34.69" />
                    <SPLIT distance="300" swimtime="00:06:58.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="298" swimtime="00:01:53.85" resultid="7723" heatid="10236" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1686" points="473" swimtime="00:06:59.67" resultid="7724" heatid="10287" lane="7" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.11" />
                    <SPLIT distance="200" swimtime="00:03:35.64" />
                    <SPLIT distance="300" swimtime="00:05:22.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+77" swimtime="00:02:27.92" resultid="5897" heatid="10161" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5770" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5708" number="2" />
                    <RELAYPOSITION athleteid="5858" number="3" />
                    <RELAYPOSITION athleteid="5836" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:02:02.59" resultid="5898" heatid="10208" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5858" number="1" />
                    <RELAYPOSITION athleteid="5708" number="2" />
                    <RELAYPOSITION athleteid="5836" number="3" />
                    <RELAYPOSITION athleteid="5770" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Masters Korona Kraków D" number="2">
              <RESULTS>
                <RESULT eventid="1260" reactiontime="+76" swimtime="00:02:20.55" resultid="5899" heatid="10161" lane="2" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5726" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5819" number="2" />
                    <RELAYPOSITION athleteid="5721" number="3" />
                    <RELAYPOSITION athleteid="7716" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1433" swimtime="00:02:05.72" resultid="5900" heatid="10208" lane="2" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5721" number="2" />
                    <RELAYPOSITION athleteid="5819" number="3" />
                    <RELAYPOSITION athleteid="5726" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kraków 0" number="1">
              <RESULTS>
                <RESULT eventid="1244" reactiontime="+87" swimtime="00:02:32.01" resultid="5901" heatid="10159" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5848" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="5870" number="2" />
                    <RELAYPOSITION athleteid="5747" number="3" />
                    <RELAYPOSITION athleteid="5878" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1417" swimtime="00:02:07.15" resultid="7739" heatid="10206" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5747" number="1" />
                    <RELAYPOSITION athleteid="5870" number="2" />
                    <RELAYPOSITION athleteid="5848" number="3" />
                    <RELAYPOSITION athleteid="5740" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Masters Korona Kraków C" number="2">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1244" reactiontime="+73" swimtime="00:02:27.75" resultid="5903" heatid="10159" lane="6" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5812" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5832" number="2" />
                    <RELAYPOSITION athleteid="5830" number="3" />
                    <RELAYPOSITION athleteid="5760" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1417" swimtime="00:02:13.58" resultid="5904" heatid="10206" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5760" number="1" />
                    <RELAYPOSITION athleteid="5830" number="2" />
                    <RELAYPOSITION athleteid="5812" number="3" />
                    <RELAYPOSITION athleteid="5832" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+104" swimtime="00:02:30.06" resultid="5889" heatid="10269" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5732" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="5765" number="2" />
                    <RELAYPOSITION athleteid="5770" number="3" />
                    <RELAYPOSITION athleteid="5836" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" status="DSQ" swimtime="00:01:59.57" resultid="7725" heatid="10125" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5760" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="5770" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="5812" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="5726" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:12.91" resultid="5892" heatid="10125" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5858" number="1" />
                    <RELAYPOSITION athleteid="5765" number="2" />
                    <RELAYPOSITION athleteid="5830" number="3" />
                    <RELAYPOSITION athleteid="5708" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+103" swimtime="00:02:16.71" resultid="5893" heatid="10269" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5812" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="5819" number="2" />
                    <RELAYPOSITION athleteid="5721" number="3" />
                    <RELAYPOSITION athleteid="5760" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Masters Korona Kraków D" number="3">
              <RESULTS>
                <RESULT eventid="1125" swimtime="00:02:09.96" resultid="5894" heatid="10124" lane="4" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5819" number="1" />
                    <RELAYPOSITION athleteid="5832" number="2" />
                    <RELAYPOSITION athleteid="5785" number="3" />
                    <RELAYPOSITION athleteid="5721" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" reactiontime="+77" swimtime="00:02:29.56" resultid="5895" heatid="10268" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5726" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5832" number="2" />
                    <RELAYPOSITION athleteid="5830" number="3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Korona Kraków E" number="4">
              <RESULTS>
                <RESULT eventid="1622" reactiontime="+104" swimtime="00:03:29.16" resultid="5896" heatid="10268" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5803" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="5708" number="2" />
                    <RELAYPOSITION athleteid="5776" number="3" />
                    <RELAYPOSITION athleteid="5752" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Masters Korona Kraków 0" number="5">
              <RESULTS>
                <RESULT eventid="1622" status="DSQ" swimtime="00:00:00.00" resultid="5890" heatid="10269" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5848" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="5714" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="5747" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="5705" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1125" status="EXH" swimtime="00:02:12.09" resultid="5891" heatid="10125" lane="5" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5958" number="1" />
                    <RELAYPOSITION athleteid="5747" number="2" />
                    <RELAYPOSITION athleteid="5848" number="3" />
                    <RELAYPOSITION athleteid="5836" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" name="Sraż Miejska Miasta Kraków" nation="POL" region="KR" shortname="Sraż Miejska Kraków">
          <CONTACT city="Kraków" name="Jawień Krzysztof" phone="505593911" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-11" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="5928">
              <RESULTS>
                <RESULT eventid="1162" points="339" swimtime="00:24:23.48" resultid="5929" heatid="10297" lane="2" entrytime="00:22:00.00" />
                <RESULT eventid="1228" points="497" swimtime="00:01:07.44" resultid="5930" heatid="10147" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="1324" points="543" swimtime="00:03:04.23" resultid="5931" heatid="10177" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="491" swimtime="00:00:37.39" resultid="5932" heatid="10191" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1465" points="443" swimtime="00:02:35.24" resultid="5933" heatid="10221" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="543" swimtime="00:00:29.92" resultid="5934" heatid="10255" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1654" points="572" swimtime="00:01:20.91" resultid="5935" heatid="10280" lane="5" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" name="Ursynów Masters" nation="POL" region="MAZ">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1970-01-23" firstname="MICHAŁ" gender="M" lastname="RYBARCZYK" nation="POL" athleteid="5937">
              <RESULTS>
                <RESULT eventid="1077" points="506" swimtime="00:00:33.45" resultid="5938" heatid="10106" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1195" points="174" swimtime="00:00:50.12" resultid="5939" heatid="10135" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1228" points="495" swimtime="00:01:07.49" resultid="5940" heatid="10154" lane="6" entrytime="00:01:05.00" />
                <RESULT eventid="1401" points="174" reactiontime="+81" swimtime="00:01:48.60" resultid="5941" heatid="10200" lane="2" entrytime="00:01:40.00" />
                <RESULT eventid="1465" points="429" swimtime="00:02:36.90" resultid="5942" heatid="10220" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="492" swimtime="00:00:30.92" resultid="5943" heatid="10253" lane="2" entrytime="00:00:28.99" />
                <RESULT eventid="1686" points="394" swimtime="00:05:42.58" resultid="5944" heatid="10289" lane="2" entrytime="00:05:49.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="200" swimtime="00:02:47.58" />
                    <SPLIT distance="300" swimtime="00:04:17.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="RYSZARD" gender="M" lastname="RYBARCZYK" nation="POL" athleteid="5945">
              <RESULTS>
                <RESULT eventid="1195" points="335" swimtime="00:00:55.03" resultid="5946" heatid="10133" lane="4" entrytime="00:00:53.00" />
                <RESULT eventid="1324" points="477" swimtime="00:04:09.40" resultid="5947" heatid="10171" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="594" swimtime="00:00:45.47" resultid="5948" heatid="10185" lane="6" entrytime="00:00:47.55" />
                <RESULT eventid="1465" points="185" swimtime="00:04:31.52" resultid="5949" heatid="10215" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="437" swimtime="00:00:39.71" resultid="5950" heatid="10247" lane="7" entrytime="00:00:43.51" />
                <RESULT eventid="1654" points="540" swimtime="00:01:47.47" resultid="5951" heatid="10275" lane="7" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="MICHAŁ" gender="M" lastname="NOWAk" nation="POL" athleteid="5952">
              <RESULTS>
                <RESULT eventid="1109" points="619" swimtime="00:03:08.97" resultid="5953" heatid="10118" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="708" swimtime="00:03:18.03" resultid="5954" heatid="10175" lane="6" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="671" swimtime="00:00:39.12" resultid="5955" heatid="10190" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1497" points="534" swimtime="00:07:09.08" resultid="5956" heatid="10228" lane="5" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.07" />
                    <SPLIT distance="200" swimtime="00:03:41.17" />
                    <SPLIT distance="300" swimtime="00:05:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="729" swimtime="00:01:27.74" resultid="5957" heatid="10279" lane="7" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KPKOZ" name="Klub Pływacki Koziegłowy" nation="POL" region="WIE" shortname="KP Koziegłowy">
          <CONTACT city="Koziegłowy" email="ewaszala59@wp.pl" name="Ewa Szała" street="os. Leśne 13/21" zip="62-028" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="5969">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1093" points="657" swimtime="00:03:07.59" resultid="5970" heatid="10112" lane="7" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="573" swimtime="00:12:38.42" resultid="5971" heatid="10294" lane="4" entrytime="00:12:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="200" swimtime="00:03:00.22" />
                    <SPLIT distance="300" swimtime="00:04:36.44" />
                    <SPLIT distance="400" swimtime="00:06:12.08" />
                    <SPLIT distance="500" swimtime="00:09:25.99" />
                    <SPLIT distance="600" swimtime="00:11:04.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="579" swimtime="00:00:41.49" resultid="5972" heatid="10128" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1212" points="520" swimtime="00:01:20.87" resultid="5973" heatid="10144" lane="7" entrytime="00:01:17.00" />
                <RESULT eventid="1385" points="658" reactiontime="+95" swimtime="00:01:28.79" resultid="5974" heatid="10196" lane="3" entrytime="00:01:27.00" />
                <RESULT eventid="1481" points="612" swimtime="00:06:52.02" resultid="5975" heatid="10225" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.11" />
                    <SPLIT distance="200" swimtime="00:03:23.36" />
                    <SPLIT distance="300" swimtime="00:05:21.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1590" points="718" reactiontime="+88" swimtime="00:03:11.08" resultid="5976" heatid="10259" lane="4" entrytime="00:03:08.00" />
                <RESULT eventid="1670" points="565" swimtime="00:06:13.79" resultid="5977" heatid="10284" lane="3" entrytime="00:05:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="200" swimtime="00:03:03.21" />
                    <SPLIT distance="300" swimtime="00:04:39.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" name="Steef Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wroclaw" email="ste1@wp.pl" name="Skrzypek Stefan" street="Szewska 18" zip="50-132" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="5979">
              <RESULTS>
                <RESULT eventid="1162" points="529" swimtime="00:24:16.27" resultid="5980" heatid="10299" lane="4" entrytime="00:24:15.00" />
                <RESULT eventid="1292" points="365" swimtime="00:03:32.93" resultid="5981" heatid="10164" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="495" swimtime="00:02:46.57" resultid="5982" heatid="10218" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" points="323" swimtime="00:01:33.75" resultid="5983" heatid="10237" lane="3" entrytime="00:01:26.00" />
                <RESULT eventid="1686" points="506" swimtime="00:05:59.18" resultid="5984" heatid="10289" lane="3" entrytime="00:05:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.70" />
                    <SPLIT distance="200" swimtime="00:02:58.20" />
                    <SPLIT distance="300" swimtime="00:04:27.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKKON" name="IKS Konstancin-Jeziorna" nation="POL">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="5986">
              <RESULTS>
                <RESULT eventid="1228" points="640" swimtime="00:01:01.98" resultid="5987" heatid="10156" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="1324" points="568" swimtime="00:03:01.45" resultid="5988" heatid="10176" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="426" swimtime="00:00:39.20" resultid="5989" heatid="10189" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1465" points="603" swimtime="00:02:20.08" resultid="5990" heatid="10222" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="685" swimtime="00:00:27.69" resultid="5991" heatid="10253" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1686" points="543" swimtime="00:05:07.82" resultid="5992" heatid="10290" lane="5" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="300" swimtime="00:03:51.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POWAR" name="Śródmiejski UKS Polna Warszawa" nation="POL" shortname="Polna Warszawa">
          <CONTACT name="Przybylski Piotr" phone="501704665" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="7945">
              <RESULTS>
                <RESULT eventid="1109" points="361" swimtime="00:02:56.02" resultid="7946" heatid="10119" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="569" swimtime="00:00:34.76" resultid="7947" heatid="10190" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1574" points="519" swimtime="00:00:28.79" resultid="7948" heatid="10254" lane="2" entrytime="00:00:28.36" />
                <RESULT eventid="1654" points="468" swimtime="00:01:21.47" resultid="7949" heatid="10279" lane="6" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZWRO" name="AZS Wrocław" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1959-02-07" firstname="Piotr" gender="M" lastname="Figiel" nation="POL" athleteid="7950">
              <RESULTS>
                <RESULT eventid="1195" points="401" swimtime="00:00:41.52" resultid="7953" heatid="10137" lane="4" entrytime="00:00:37.19" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="7954" heatid="10201" lane="4" entrytime="00:01:27.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SZMAS" name="SzTP Masters" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="8143">
              <RESULTS>
                <RESULT eventid="1195" points="363" swimtime="00:00:57.43" resultid="8145" heatid="10133" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1228" points="360" swimtime="00:01:48.69" resultid="8146" heatid="10147" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="1401" points="384" reactiontime="+120" swimtime="00:02:07.85" resultid="8147" heatid="10198" lane="5" entrytime="00:02:08.00" />
                <RESULT eventid="1465" points="507" swimtime="00:04:01.46" resultid="8148" heatid="10215" lane="7" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1606" points="334" reactiontime="+126" swimtime="00:04:55.95" resultid="8149" heatid="10262" lane="8" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1654" points="497" swimtime="00:02:14.99" resultid="8150" heatid="10275" lane="1" entrytime="00:02:06.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POOST" name="Pływalnia Oceanik Ostrzeszów" nation="POL" shortname="PO Ostrzeszów">
          <CONTACT name="Burghardt" phone="660945504" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-21" firstname="Nina" gender="F" lastname="Burghardt" nation="POL" athleteid="8152">
              <RESULTS>
                <RESULT eventid="1178" points="667" swimtime="00:00:34.84" resultid="8153" heatid="10130" lane="5" entrytime="00:00:34.20" />
                <RESULT eventid="1212" points="503" swimtime="00:01:12.24" resultid="8154" heatid="10146" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1352" points="624" swimtime="00:00:39.89" resultid="8155" heatid="10182" lane="2" entrytime="00:00:38.50" />
                <RESULT eventid="1385" points="556" reactiontime="+75" swimtime="00:01:17.17" resultid="8156" heatid="10197" lane="7" entrytime="00:01:18.50" />
                <RESULT eventid="1558" points="546" swimtime="00:00:32.29" resultid="8157" heatid="10245" lane="2" entrytime="00:00:30.10" />
                <RESULT eventid="1638" points="511" swimtime="00:01:28.41" resultid="8158" heatid="10273" lane="3" entrytime="00:01:23.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPIA" name="MKS Piaseczno" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1949-04-10" firstname="Andrzej" gender="M" lastname="Rubaszkiewicz" nation="POL" athleteid="8159">
              <RESULTS>
                <RESULT eventid="1077" points="696" swimtime="00:00:34.27" resultid="8161" heatid="10106" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1195" points="705" swimtime="00:00:37.57" resultid="8162" heatid="10138" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1369" status="DNS" swimtime="00:00:00.00" resultid="8163" heatid="10188" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1574" status="DSQ" swimtime="00:00:29.94" resultid="8164" heatid="10252" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1401" points="555" reactiontime="+104" swimtime="00:01:29.51" resultid="8165" heatid="10201" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1228" points="746" swimtime="00:01:08.76" resultid="8166" heatid="10152" lane="4" entrytime="00:01:08.00" />
                <RESULT eventid="1465" points="607" swimtime="00:02:46.70" resultid="8167" heatid="10219" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1542" status="DNS" swimtime="00:00:00.00" resultid="8168" heatid="10237" lane="1" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOCZE" name="MOSiR Częstochowa" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="2252">
              <RESULTS>
                <RESULT eventid="1195" points="230" swimtime="00:00:45.73" resultid="2253" heatid="10135" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1401" points="247" reactiontime="+100" swimtime="00:01:36.75" resultid="2254" heatid="10200" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1606" points="264" reactiontime="+105" swimtime="00:03:31.02" resultid="2255" heatid="10263" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIKON" name="Niezrzeszony KONIN" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1993-12-09" firstname="Norbert" gender="M" lastname="Cezak" nation="POL" athleteid="4430">
              <RESULTS>
                <RESULT eventid="1228" status="DSQ" swimtime="00:01:03.47" resultid="4431" heatid="10158" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="1324" points="442" swimtime="00:02:56.94" resultid="4432" heatid="10177" lane="3" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="458" swimtime="00:00:36.73" resultid="4433" heatid="10191" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1465" points="371" swimtime="00:02:29.78" resultid="4434" heatid="10221" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1574" points="527" swimtime="00:00:27.62" resultid="4435" heatid="10257" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1654" points="457" swimtime="00:01:20.68" resultid="4436" heatid="10281" lane="6" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1709" code="1" course="LCM" gender="M" name="Minima " type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:30:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1711" code="1" course="LCM" gender="F" name="Minima " type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:22:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SiKReT Gliwice" version="11.42512">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Gliwice" name="Letnie Mistrzostwa Polski w Pływaniu Masters" course="LCM" hostclub="SiKReT Gliwice" hostclub.url="http://www.sikret-plywanie.pl" nation="POL" organizer="Samorząd Miasta Gliwice, MZUK Gliwice, PZP,SLOZP,SiKReT Gliwice" reservecount="2" result.url="http://www.megatiming.pl" startmethod="1" timing="AUTOMATIC">
      <AGEDATE value="2016-06-10" type="YEAR" />
      <POOL name="Olimpijczyk Gliwice" lanemax="9" />
      <POINTTABLE pointtableid="3009" name="FINA Point Scoring" version="2016" />
      <CONTACT email="wisniowicz@interia.pl" name="Wojciech Wiśniowicz" phone="500193225" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="11000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="15000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2016-06-10" daytime="15:45" endtime="21:28" name="BLOK I" number="1" warmupfrom="14:30">
          <EVENTS>
            <EVENT eventid="1062" daytime="16:00" gender="F" number="1" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10913" />
                    <RANKING order="2" place="2" resultid="11086" />
                    <RANKING order="3" place="3" resultid="10497" />
                    <RANKING order="4" place="4" resultid="10482" />
                    <RANKING order="5" place="5" resultid="9984" />
                    <RANKING order="6" place="-1" resultid="10133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12101" />
                    <RANKING order="2" place="2" resultid="10092" />
                    <RANKING order="3" place="3" resultid="10126" />
                    <RANKING order="4" place="4" resultid="12766" />
                    <RANKING order="5" place="5" resultid="9834" />
                    <RANKING order="6" place="-1" resultid="12176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12759" />
                    <RANKING order="2" place="2" resultid="11656" />
                    <RANKING order="3" place="3" resultid="10518" />
                    <RANKING order="4" place="4" resultid="12356" />
                    <RANKING order="5" place="5" resultid="10276" />
                    <RANKING order="6" place="6" resultid="10153" />
                    <RANKING order="7" place="7" resultid="11665" />
                    <RANKING order="8" place="-1" resultid="10342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11064" />
                    <RANKING order="2" place="2" resultid="12426" />
                    <RANKING order="3" place="3" resultid="12435" />
                    <RANKING order="4" place="4" resultid="11836" />
                    <RANKING order="5" place="5" resultid="11734" />
                    <RANKING order="6" place="6" resultid="9655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9553" />
                    <RANKING order="2" place="2" resultid="11514" />
                    <RANKING order="3" place="3" resultid="12238" />
                    <RANKING order="4" place="4" resultid="11945" />
                    <RANKING order="5" place="5" resultid="10454" />
                    <RANKING order="6" place="6" resultid="11478" />
                    <RANKING order="7" place="7" resultid="10769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11389" />
                    <RANKING order="2" place="2" resultid="12231" />
                    <RANKING order="3" place="3" resultid="9913" />
                    <RANKING order="4" place="4" resultid="11583" />
                    <RANKING order="5" place="5" resultid="10774" />
                    <RANKING order="6" place="6" resultid="10415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11393" />
                    <RANKING order="2" place="2" resultid="9513" />
                    <RANKING order="3" place="3" resultid="9505" />
                    <RANKING order="4" place="4" resultid="11307" />
                    <RANKING order="5" place="-1" resultid="11991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11458" />
                    <RANKING order="2" place="2" resultid="11285" />
                    <RANKING order="3" place="3" resultid="12095" />
                    <RANKING order="4" place="4" resultid="11439" />
                    <RANKING order="5" place="5" resultid="9670" />
                    <RANKING order="6" place="6" resultid="12245" />
                    <RANKING order="7" place="7" resultid="9662" />
                    <RANKING order="8" place="8" resultid="11370" />
                    <RANKING order="9" place="9" resultid="10467" />
                    <RANKING order="10" place="10" resultid="9967" />
                    <RANKING order="11" place="-1" resultid="11467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9498" />
                    <RANKING order="2" place="2" resultid="10406" />
                    <RANKING order="3" place="3" resultid="9849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10289" />
                    <RANKING order="2" place="2" resultid="12123" />
                    <RANKING order="3" place="3" resultid="9950" />
                    <RANKING order="4" place="-1" resultid="10724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1076" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1077" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1078" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1063" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13896" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13897" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13898" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13899" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13900" daytime="16:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13901" daytime="16:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13902" daytime="16:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="17:40" gender="X" number="5" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12486" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12821" />
                    <RANKING order="2" place="2" resultid="11540" />
                    <RANKING order="3" place="3" resultid="11905" />
                    <RANKING order="4" place="4" resultid="10546" />
                    <RANKING order="5" place="5" resultid="10358" />
                    <RANKING order="6" place="6" resultid="11750" />
                    <RANKING order="7" place="7" resultid="10359" />
                    <RANKING order="8" place="8" resultid="10829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11480" />
                    <RANKING order="2" place="2" resultid="9565" />
                    <RANKING order="3" place="3" resultid="11904" />
                    <RANKING order="4" place="4" resultid="12281" />
                    <RANKING order="5" place="-1" resultid="12120" />
                    <RANKING order="6" place="-1" resultid="12283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11345" />
                    <RANKING order="2" place="2" resultid="9699" />
                    <RANKING order="3" place="3" resultid="10545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9567" />
                    <RANKING order="2" place="2" resultid="11486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9982" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13932" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13933" daytime="17:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13934" daytime="17:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="17:50" gender="F" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12102" />
                    <RANKING order="2" place="2" resultid="10885" />
                    <RANKING order="3" place="3" resultid="11675" />
                    <RANKING order="4" place="4" resultid="12253" />
                    <RANKING order="5" place="-1" resultid="9835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10519" />
                    <RANKING order="2" place="2" resultid="11666" />
                    <RANKING order="3" place="3" resultid="12774" />
                    <RANKING order="4" place="4" resultid="11929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10086" />
                    <RANKING order="2" place="2" resultid="11828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10729" />
                    <RANKING order="2" place="2" resultid="10100" />
                    <RANKING order="3" place="3" resultid="11515" />
                    <RANKING order="4" place="4" resultid="11946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11291" />
                    <RANKING order="2" place="2" resultid="9841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12096" />
                    <RANKING order="2" place="2" resultid="11105" />
                    <RANKING order="3" place="3" resultid="11459" />
                    <RANKING order="4" place="4" resultid="11371" />
                    <RANKING order="5" place="-1" resultid="9968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1160" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1161" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1162" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1163" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1164" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13935" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13936" daytime="18:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13937" daytime="18:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="16:55" gender="M" number="4" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12361" />
                    <RANKING order="2" place="2" resultid="12465" />
                    <RANKING order="3" place="3" resultid="10879" />
                    <RANKING order="4" place="-1" resultid="9731" />
                    <RANKING order="5" place="-1" resultid="10941" />
                    <RANKING order="6" place="-1" resultid="11637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12406" />
                    <RANKING order="2" place="2" resultid="9535" />
                    <RANKING order="3" place="3" resultid="12182" />
                    <RANKING order="4" place="4" resultid="11560" />
                    <RANKING order="5" place="5" resultid="10107" />
                    <RANKING order="6" place="6" resultid="10923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12796" />
                    <RANKING order="2" place="2" resultid="11025" />
                    <RANKING order="3" place="3" resultid="11709" />
                    <RANKING order="4" place="4" resultid="10301" />
                    <RANKING order="5" place="5" resultid="10147" />
                    <RANKING order="6" place="6" resultid="10988" />
                    <RANKING order="7" place="7" resultid="12787" />
                    <RANKING order="8" place="8" resultid="10212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11298" />
                    <RANKING order="2" place="2" resultid="9607" />
                    <RANKING order="3" place="3" resultid="10961" />
                    <RANKING order="4" place="4" resultid="10954" />
                    <RANKING order="5" place="5" resultid="11719" />
                    <RANKING order="6" place="6" resultid="11074" />
                    <RANKING order="7" place="7" resultid="11330" />
                    <RANKING order="8" place="8" resultid="12368" />
                    <RANKING order="9" place="9" resultid="9522" />
                    <RANKING order="10" place="10" resultid="11617" />
                    <RANKING order="11" place="11" resultid="10678" />
                    <RANKING order="12" place="12" resultid="9687" />
                    <RANKING order="13" place="13" resultid="10969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11624" />
                    <RANKING order="2" place="2" resultid="11848" />
                    <RANKING order="3" place="3" resultid="10316" />
                    <RANKING order="4" place="4" resultid="11592" />
                    <RANKING order="5" place="5" resultid="11857" />
                    <RANKING order="6" place="6" resultid="11527" />
                    <RANKING order="7" place="7" resultid="10981" />
                    <RANKING order="8" place="8" resultid="10740" />
                    <RANKING order="9" place="9" resultid="10389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11684" />
                    <RANKING order="2" place="2" resultid="10339" />
                    <RANKING order="3" place="3" resultid="10427" />
                    <RANKING order="4" place="4" resultid="11894" />
                    <RANKING order="5" place="5" resultid="11176" />
                    <RANKING order="6" place="6" resultid="10869" />
                    <RANKING order="7" place="7" resultid="9906" />
                    <RANKING order="8" place="8" resultid="11506" />
                    <RANKING order="9" place="9" resultid="12265" />
                    <RANKING order="10" place="10" resultid="10528" />
                    <RANKING order="11" place="11" resultid="12213" />
                    <RANKING order="12" place="-1" resultid="11700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9828" />
                    <RANKING order="2" place="2" resultid="11013" />
                    <RANKING order="3" place="3" resultid="10221" />
                    <RANKING order="4" place="4" resultid="9714" />
                    <RANKING order="5" place="5" resultid="12154" />
                    <RANKING order="6" place="6" resultid="12112" />
                    <RANKING order="7" place="7" resultid="12323" />
                    <RANKING order="8" place="8" resultid="11324" />
                    <RANKING order="9" place="9" resultid="9897" />
                    <RANKING order="10" place="-1" resultid="10394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9490" />
                    <RANKING order="2" place="2" resultid="11608" />
                    <RANKING order="3" place="3" resultid="9638" />
                    <RANKING order="4" place="4" resultid="12146" />
                    <RANKING order="5" place="5" resultid="11807" />
                    <RANKING order="6" place="6" resultid="9620" />
                    <RANKING order="7" place="7" resultid="11362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10206" />
                    <RANKING order="2" place="2" resultid="9770" />
                    <RANKING order="3" place="3" resultid="12193" />
                    <RANKING order="4" place="4" resultid="12138" />
                    <RANKING order="5" place="5" resultid="9721" />
                    <RANKING order="6" place="6" resultid="11007" />
                    <RANKING order="7" place="7" resultid="9649" />
                    <RANKING order="8" place="8" resultid="9863" />
                    <RANKING order="9" place="9" resultid="11572" />
                    <RANKING order="10" place="10" resultid="11816" />
                    <RANKING order="11" place="11" resultid="10050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9528" />
                    <RANKING order="2" place="2" resultid="11408" />
                    <RANKING order="3" place="3" resultid="10815" />
                    <RANKING order="4" place="4" resultid="12416" />
                    <RANKING order="5" place="5" resultid="10000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9593" />
                    <RANKING order="2" place="2" resultid="9888" />
                    <RANKING order="3" place="3" resultid="11443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9976" />
                    <RANKING order="2" place="-1" resultid="9879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1127" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1129" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13922" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13923" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13924" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13925" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13926" daytime="17:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13927" daytime="17:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13928" daytime="17:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13929" daytime="17:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="13930" daytime="17:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="13931" daytime="17:35" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="16:35" gender="F" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10139" />
                    <RANKING order="2" place="2" resultid="11087" />
                    <RANKING order="3" place="3" resultid="10914" />
                    <RANKING order="4" place="4" resultid="10483" />
                    <RANKING order="5" place="-1" resultid="10134" />
                    <RANKING order="6" place="-1" resultid="10498" />
                    <RANKING order="7" place="-1" resultid="10931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10884" />
                    <RANKING order="2" place="2" resultid="11674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11657" />
                    <RANKING order="2" place="2" resultid="10023" />
                    <RANKING order="3" place="3" resultid="11928" />
                    <RANKING order="4" place="4" resultid="10343" />
                    <RANKING order="5" place="5" resultid="10311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11065" />
                    <RANKING order="2" place="2" resultid="12427" />
                    <RANKING order="3" place="3" resultid="11886" />
                    <RANKING order="4" place="4" resultid="12436" />
                    <RANKING order="5" place="-1" resultid="10460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9554" />
                    <RANKING order="2" place="2" resultid="11727" />
                    <RANKING order="3" place="3" resultid="11479" />
                    <RANKING order="4" place="4" resultid="11823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9542" />
                    <RANKING order="2" place="2" resultid="11584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11308" />
                    <RANKING order="2" place="2" resultid="9840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11104" />
                    <RANKING order="2" place="2" resultid="10763" />
                    <RANKING order="3" place="3" resultid="11440" />
                    <RANKING order="4" place="4" resultid="12246" />
                    <RANKING order="5" place="5" resultid="9671" />
                    <RANKING order="6" place="6" resultid="10468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10407" />
                    <RANKING order="2" place="2" resultid="9959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1110" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1111" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1112" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13918" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13919" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13920" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13921" daytime="16:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="16:10" gender="M" number="2" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12170" />
                    <RANKING order="2" place="2" resultid="12464" />
                    <RANKING order="3" place="3" resultid="10446" />
                    <RANKING order="4" place="4" resultid="11690" />
                    <RANKING order="5" place="-1" resultid="9730" />
                    <RANKING order="6" place="-1" resultid="10940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12443" />
                    <RANKING order="2" place="2" resultid="9534" />
                    <RANKING order="3" place="3" resultid="10890" />
                    <RANKING order="4" place="4" resultid="10295" />
                    <RANKING order="5" place="5" resultid="12181" />
                    <RANKING order="6" place="6" resultid="10491" />
                    <RANKING order="7" place="7" resultid="12450" />
                    <RANKING order="8" place="8" resultid="10874" />
                    <RANKING order="9" place="9" resultid="10106" />
                    <RANKING order="10" place="10" resultid="10785" />
                    <RANKING order="11" place="11" resultid="10688" />
                    <RANKING order="12" place="12" resultid="12332" />
                    <RANKING order="13" place="13" resultid="10780" />
                    <RANKING order="14" place="14" resultid="9616" />
                    <RANKING order="15" place="-1" resultid="10922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12781" />
                    <RANKING order="2" place="2" resultid="12795" />
                    <RANKING order="3" place="3" resultid="12786" />
                    <RANKING order="4" place="4" resultid="11429" />
                    <RANKING order="5" place="5" resultid="12188" />
                    <RANKING order="6" place="6" resultid="11024" />
                    <RANKING order="7" place="7" resultid="10146" />
                    <RANKING order="8" place="8" resultid="11997" />
                    <RANKING order="9" place="9" resultid="12166" />
                    <RANKING order="10" place="10" resultid="10030" />
                    <RANKING order="11" place="11" resultid="10120" />
                    <RANKING order="12" place="12" resultid="12341" />
                    <RANKING order="13" place="13" resultid="9918" />
                    <RANKING order="14" place="14" resultid="10211" />
                    <RANKING order="15" place="15" resultid="11472" />
                    <RANKING order="16" place="-1" resultid="10709" />
                    <RANKING order="17" place="-1" resultid="11570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9606" />
                    <RANKING order="2" place="2" resultid="10347" />
                    <RANKING order="3" place="3" resultid="11650" />
                    <RANKING order="4" place="4" resultid="12367" />
                    <RANKING order="5" place="5" resultid="10535" />
                    <RANKING order="6" place="6" resultid="12350" />
                    <RANKING order="7" place="7" resultid="11318" />
                    <RANKING order="8" place="8" resultid="10976" />
                    <RANKING order="9" place="9" resultid="11329" />
                    <RANKING order="10" place="10" resultid="11718" />
                    <RANKING order="11" place="11" resultid="9686" />
                    <RANKING order="12" place="12" resultid="9858" />
                    <RANKING order="13" place="13" resultid="10038" />
                    <RANKING order="14" place="14" resultid="10968" />
                    <RANKING order="15" place="15" resultid="12272" />
                    <RANKING order="16" place="16" resultid="11616" />
                    <RANKING order="17" place="17" resultid="10439" />
                    <RANKING order="18" place="-1" resultid="10960" />
                    <RANKING order="19" place="-1" resultid="10949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11535" />
                    <RANKING order="2" place="2" resultid="10671" />
                    <RANKING order="3" place="3" resultid="12315" />
                    <RANKING order="4" place="4" resultid="11847" />
                    <RANKING order="5" place="5" resultid="11623" />
                    <RANKING order="6" place="6" resultid="12277" />
                    <RANKING order="7" place="7" resultid="11591" />
                    <RANKING order="8" place="8" resultid="9693" />
                    <RANKING order="9" place="9" resultid="11522" />
                    <RANKING order="10" place="10" resultid="11865" />
                    <RANKING order="11" place="11" resultid="10683" />
                    <RANKING order="12" place="12" resultid="11856" />
                    <RANKING order="13" place="13" resultid="10712" />
                    <RANKING order="14" place="14" resultid="10115" />
                    <RANKING order="15" place="15" resultid="11875" />
                    <RANKING order="16" place="16" resultid="10760" />
                    <RANKING order="17" place="17" resultid="9935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11699" />
                    <RANKING order="2" place="2" resultid="12755" />
                    <RANKING order="3" place="3" resultid="10338" />
                    <RANKING order="4" place="4" resultid="11683" />
                    <RANKING order="5" place="5" resultid="10426" />
                    <RANKING order="6" place="6" resultid="10868" />
                    <RANKING order="7" place="7" resultid="11056" />
                    <RANKING order="8" place="8" resultid="11171" />
                    <RANKING order="9" place="9" resultid="11600" />
                    <RANKING order="10" place="10" resultid="10527" />
                    <RANKING order="11" place="11" resultid="12198" />
                    <RANKING order="12" place="12" resultid="12212" />
                    <RANKING order="13" place="13" resultid="10270" />
                    <RANKING order="14" place="14" resultid="12447" />
                    <RANKING order="15" place="15" resultid="10435" />
                    <RANKING order="16" place="16" resultid="10752" />
                    <RANKING order="17" place="-1" resultid="11900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10228" />
                    <RANKING order="2" place="2" resultid="9827" />
                    <RANKING order="3" place="3" resultid="11012" />
                    <RANKING order="4" place="4" resultid="10220" />
                    <RANKING order="5" place="5" resultid="9713" />
                    <RANKING order="6" place="6" resultid="11278" />
                    <RANKING order="7" place="7" resultid="11962" />
                    <RANKING order="8" place="8" resultid="11400" />
                    <RANKING order="9" place="9" resultid="9896" />
                    <RANKING order="10" place="10" resultid="9679" />
                    <RANKING order="11" place="11" resultid="10803" />
                    <RANKING order="12" place="12" resultid="10263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11554" />
                    <RANKING order="2" place="2" resultid="9489" />
                    <RANKING order="3" place="3" resultid="11979" />
                    <RANKING order="4" place="4" resultid="11607" />
                    <RANKING order="5" place="5" resultid="10719" />
                    <RANKING order="6" place="6" resultid="9751" />
                    <RANKING order="7" place="7" resultid="12456" />
                    <RANKING order="8" place="8" resultid="9923" />
                    <RANKING order="9" place="9" resultid="12107" />
                    <RANKING order="10" place="10" resultid="11361" />
                    <RANKING order="11" place="11" resultid="10235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9601" />
                    <RANKING order="2" place="2" resultid="11006" />
                    <RANKING order="3" place="3" resultid="9408" />
                    <RANKING order="4" place="4" resultid="10015" />
                    <RANKING order="5" place="5" resultid="11954" />
                    <RANKING order="6" place="6" resultid="9648" />
                    <RANKING order="7" place="7" resultid="9937" />
                    <RANKING order="8" place="8" resultid="9695" />
                    <RANKING order="9" place="9" resultid="11543" />
                    <RANKING order="10" place="10" resultid="10505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9527" />
                    <RANKING order="2" place="2" resultid="10249" />
                    <RANKING order="3" place="3" resultid="11407" />
                    <RANKING order="4" place="4" resultid="12132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9592" />
                    <RANKING order="2" place="2" resultid="10182" />
                    <RANKING order="3" place="3" resultid="9398" />
                    <RANKING order="4" place="4" resultid="12206" />
                    <RANKING order="5" place="5" resultid="10008" />
                    <RANKING order="6" place="6" resultid="11442" />
                    <RANKING order="7" place="7" resultid="11377" />
                    <RANKING order="8" place="8" resultid="9887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11017" />
                    <RANKING order="2" place="2" resultid="9975" />
                    <RANKING order="3" place="3" resultid="11971" />
                    <RANKING order="4" place="4" resultid="11382" />
                    <RANKING order="5" place="5" resultid="9992" />
                    <RANKING order="6" place="6" resultid="9878" />
                    <RANKING order="7" place="7" resultid="9997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10511" />
                    <RANKING order="2" place="2" resultid="12387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1095" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13903" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13904" daytime="16:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13905" daytime="16:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13906" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13907" daytime="16:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13908" daytime="16:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13909" daytime="16:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13910" daytime="16:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="13911" daytime="16:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="13912" daytime="16:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="13913" daytime="16:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="13914" daytime="16:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="13915" daytime="16:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="13916" daytime="16:30" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="13917" daytime="16:35" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="18:35" gender="M" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12396" />
                    <RANKING order="2" place="2" resultid="9428" />
                    <RANKING order="3" place="3" resultid="10544" />
                    <RANKING order="4" place="-1" resultid="11691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12407" />
                    <RANKING order="2" place="2" resultid="11561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11710" />
                    <RANKING order="2" place="-1" resultid="12342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11299" />
                    <RANKING order="2" place="2" resultid="10200" />
                    <RANKING order="3" place="-1" resultid="10440" />
                    <RANKING order="4" place="-1" resultid="10536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12316" />
                    <RANKING order="2" place="2" resultid="11082" />
                    <RANKING order="3" place="3" resultid="11455" />
                    <RANKING order="4" place="4" resultid="9612" />
                    <RANKING order="5" place="5" resultid="10317" />
                    <RANKING order="6" place="6" resultid="11548" />
                    <RANKING order="7" place="7" resultid="10327" />
                    <RANKING order="8" place="-1" resultid="11876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9391" />
                    <RANKING order="2" place="2" resultid="9626" />
                    <RANKING order="3" place="-1" resultid="10340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11279" />
                    <RANKING order="2" place="2" resultid="11963" />
                    <RANKING order="3" place="3" resultid="12324" />
                    <RANKING order="4" place="4" resultid="11432" />
                    <RANKING order="5" place="5" resultid="11271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11555" />
                    <RANKING order="2" place="2" resultid="9639" />
                    <RANKING order="3" place="3" resultid="12457" />
                    <RANKING order="4" place="4" resultid="11808" />
                    <RANKING order="5" place="5" resultid="9621" />
                    <RANKING order="6" place="6" resultid="9752" />
                    <RANKING order="7" place="-1" resultid="9628" />
                    <RANKING order="8" place="-1" resultid="10236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11112" />
                    <RANKING order="2" place="2" resultid="10016" />
                    <RANKING order="3" place="3" resultid="9864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10250" />
                    <RANKING order="2" place="-1" resultid="12417" />
                    <RANKING order="3" place="-1" resultid="9350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9399" />
                    <RANKING order="2" place="2" resultid="10183" />
                    <RANKING order="3" place="-1" resultid="9417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9356" />
                    <RANKING order="2" place="2" resultid="11383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1181" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13938" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13939" daytime="18:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13940" daytime="19:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13941" daytime="19:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13942" daytime="20:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13943" daytime="20:40" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-06-11" daytime="09:00" endtime="12:24" name="BLOK II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1187" daytime="09:00" gender="F" number="8" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11801" />
                    <RANKING order="2" place="2" resultid="10915" />
                    <RANKING order="3" place="3" resultid="11088" />
                    <RANKING order="4" place="4" resultid="10933" />
                    <RANKING order="5" place="5" resultid="9985" />
                    <RANKING order="6" place="-1" resultid="10135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10401" />
                    <RANKING order="2" place="2" resultid="11676" />
                    <RANKING order="3" place="3" resultid="10127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11658" />
                    <RANKING order="2" place="2" resultid="10520" />
                    <RANKING order="3" place="3" resultid="9630" />
                    <RANKING order="4" place="4" resultid="11532" />
                    <RANKING order="5" place="5" resultid="10154" />
                    <RANKING order="6" place="6" resultid="11930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10081" />
                    <RANKING order="2" place="2" resultid="11066" />
                    <RANKING order="3" place="3" resultid="11829" />
                    <RANKING order="4" place="4" resultid="11837" />
                    <RANKING order="5" place="5" resultid="11735" />
                    <RANKING order="6" place="-1" resultid="11887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9555" />
                    <RANKING order="2" place="2" resultid="11728" />
                    <RANKING order="3" place="3" resultid="10455" />
                    <RANKING order="4" place="4" resultid="12239" />
                    <RANKING order="5" place="5" resultid="10770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12306" />
                    <RANKING order="2" place="2" resultid="10903" />
                    <RANKING order="3" place="3" resultid="12232" />
                    <RANKING order="4" place="4" resultid="10416" />
                    <RANKING order="5" place="-1" resultid="12080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11394" />
                    <RANKING order="2" place="2" resultid="9506" />
                    <RANKING order="3" place="3" resultid="11292" />
                    <RANKING order="4" place="4" resultid="11309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11052" />
                    <RANKING order="2" place="2" resultid="9672" />
                    <RANKING order="3" place="3" resultid="12247" />
                    <RANKING order="4" place="4" resultid="10469" />
                    <RANKING order="5" place="5" resultid="10717" />
                    <RANKING order="6" place="6" resultid="9969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9499" />
                    <RANKING order="2" place="2" resultid="10408" />
                    <RANKING order="3" place="3" resultid="9960" />
                    <RANKING order="4" place="4" resultid="9851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10290" />
                    <RANKING order="2" place="2" resultid="12125" />
                    <RANKING order="3" place="3" resultid="9951" />
                    <RANKING order="4" place="4" resultid="11644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1200" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1202" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1203" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1204" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13944" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13945" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13946" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13947" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13948" daytime="09:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="11:10" gender="F" number="14" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10521" />
                    <RANKING order="2" place="2" resultid="11668" />
                    <RANKING order="3" place="3" resultid="11931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11067" />
                    <RANKING order="2" place="2" resultid="12429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1330" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9507" />
                    <RANKING order="2" place="2" resultid="9843" />
                    <RANKING order="3" place="3" resultid="11310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1332" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11106" />
                    <RANKING order="2" place="2" resultid="11372" />
                    <RANKING order="3" place="3" resultid="9664" />
                    <RANKING order="4" place="-1" resultid="11461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1335" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1336" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1338" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1339" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1340" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13990" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13991" daytime="11:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="09:25" gender="F" number="10" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10421" />
                    <RANKING order="2" place="2" resultid="10499" />
                    <RANKING order="3" place="3" resultid="10484" />
                    <RANKING order="4" place="4" resultid="10916" />
                    <RANKING order="5" place="5" resultid="10934" />
                    <RANKING order="6" place="6" resultid="10285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10093" />
                    <RANKING order="2" place="2" resultid="12767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12760" />
                    <RANKING order="2" place="2" resultid="10024" />
                    <RANKING order="3" place="3" resultid="10277" />
                    <RANKING order="4" place="4" resultid="12775" />
                    <RANKING order="5" place="5" resultid="11744" />
                    <RANKING order="6" place="6" resultid="10312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11888" />
                    <RANKING order="2" place="2" resultid="12437" />
                    <RANKING order="3" place="3" resultid="11830" />
                    <RANKING order="4" place="4" resultid="9656" />
                    <RANKING order="5" place="-1" resultid="10461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10730" />
                    <RANKING order="2" place="2" resultid="11947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11585" />
                    <RANKING order="2" place="2" resultid="11938" />
                    <RANKING order="3" place="3" resultid="10775" />
                    <RANKING order="4" place="4" resultid="10417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11468" />
                    <RANKING order="2" place="2" resultid="11286" />
                    <RANKING order="3" place="3" resultid="9663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10706" />
                    <RANKING order="2" place="2" resultid="11418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1238" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13959" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13960" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13961" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13962" daytime="09:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1341" daytime="11:20" gender="M" number="15" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1342" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1343" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12409" />
                    <RANKING order="2" place="2" resultid="10109" />
                    <RANKING order="3" place="3" resultid="11562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12798" />
                    <RANKING order="2" place="2" resultid="11712" />
                    <RANKING order="3" place="3" resultid="10990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11301" />
                    <RANKING order="2" place="2" resultid="11721" />
                    <RANKING order="3" place="3" resultid="10680" />
                    <RANKING order="4" place="4" resultid="10039" />
                    <RANKING order="5" place="5" resultid="11619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11456" />
                    <RANKING order="2" place="2" resultid="9613" />
                    <RANKING order="3" place="3" resultid="10713" />
                    <RANKING order="4" place="4" resultid="10741" />
                    <RANKING order="5" place="-1" resultid="11878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9393" />
                    <RANKING order="2" place="2" resultid="11508" />
                    <RANKING order="3" place="3" resultid="11602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11965" />
                    <RANKING order="2" place="2" resultid="11272" />
                    <RANKING order="3" place="3" resultid="12326" />
                    <RANKING order="4" place="4" resultid="10396" />
                    <RANKING order="5" place="5" resultid="10808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9492" />
                    <RANKING order="2" place="2" resultid="9640" />
                    <RANKING order="3" place="3" resultid="12148" />
                    <RANKING order="4" place="4" resultid="11364" />
                    <RANKING order="5" place="5" resultid="9754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9723" />
                    <RANKING order="2" place="2" resultid="11113" />
                    <RANKING order="3" place="3" resultid="11956" />
                    <RANKING order="4" place="4" resultid="9866" />
                    <RANKING order="5" place="-1" resultid="12140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9530" />
                    <RANKING order="2" place="2" resultid="11410" />
                    <RANKING order="3" place="3" resultid="10002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1353" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1355" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1356" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1357" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13992" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13993" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13994" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13995" daytime="11:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="09:45" gender="M" number="11" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12362" />
                    <RANKING order="2" place="2" resultid="12467" />
                    <RANKING order="3" place="3" resultid="11639" />
                    <RANKING order="4" place="4" resultid="11097" />
                    <RANKING order="5" place="-1" resultid="9733" />
                    <RANKING order="6" place="-1" resultid="10880" />
                    <RANKING order="7" place="-1" resultid="12400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12408" />
                    <RANKING order="2" place="2" resultid="11474" />
                    <RANKING order="3" place="3" resultid="10195" />
                    <RANKING order="4" place="4" resultid="10925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10303" />
                    <RANKING order="2" place="2" resultid="10351" />
                    <RANKING order="3" place="3" resultid="10031" />
                    <RANKING order="4" place="4" resultid="12072" />
                    <RANKING order="5" place="-1" resultid="12472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11300" />
                    <RANKING order="2" place="2" resultid="11331" />
                    <RANKING order="3" place="3" resultid="10955" />
                    <RANKING order="4" place="4" resultid="11618" />
                    <RANKING order="5" place="5" resultid="11076" />
                    <RANKING order="6" place="6" resultid="12084" />
                    <RANKING order="7" place="-1" resultid="10281" />
                    <RANKING order="8" place="-1" resultid="10971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10672" />
                    <RANKING order="2" place="2" resultid="11859" />
                    <RANKING order="3" place="3" resultid="11450" />
                    <RANKING order="4" place="4" resultid="10077" />
                    <RANKING order="5" place="5" resultid="11528" />
                    <RANKING order="6" place="6" resultid="10390" />
                    <RANKING order="7" place="-1" resultid="12260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9740" />
                    <RANKING order="2" place="2" resultid="10898" />
                    <RANKING order="3" place="3" resultid="11895" />
                    <RANKING order="4" place="4" resultid="11507" />
                    <RANKING order="5" place="5" resultid="10073" />
                    <RANKING order="6" place="6" resultid="9760" />
                    <RANKING order="7" place="7" resultid="9392" />
                    <RANKING order="8" place="8" resultid="10753" />
                    <RANKING order="9" place="-1" resultid="9908" />
                    <RANKING order="10" place="-1" resultid="10428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12113" />
                    <RANKING order="2" place="2" resultid="11325" />
                    <RANKING order="3" place="3" resultid="12155" />
                    <RANKING order="4" place="4" resultid="10264" />
                    <RANKING order="5" place="5" resultid="10791" />
                    <RANKING order="6" place="6" resultid="9898" />
                    <RANKING order="7" place="-1" resultid="10229" />
                    <RANKING order="8" place="-1" resultid="9548" />
                    <RANKING order="9" place="-1" resultid="10395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11980" />
                    <RANKING order="2" place="2" resultid="12147" />
                    <RANKING order="3" place="3" resultid="11046" />
                    <RANKING order="4" place="4" resultid="9485" />
                    <RANKING order="5" place="5" resultid="11363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12194" />
                    <RANKING order="2" place="2" resultid="9947" />
                    <RANKING order="3" place="3" resultid="11030" />
                    <RANKING order="4" place="4" resultid="11817" />
                    <RANKING order="5" place="5" resultid="10811" />
                    <RANKING order="6" place="6" resultid="9765" />
                    <RANKING order="7" place="-1" resultid="9722" />
                    <RANKING order="8" place="-1" resultid="11573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9481" />
                    <RANKING order="2" place="2" resultid="12419" />
                    <RANKING order="3" place="3" resultid="12064" />
                    <RANKING order="4" place="4" resultid="10541" />
                    <RANKING order="5" place="5" resultid="10001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9594" />
                    <RANKING order="2" place="2" resultid="10010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10703" />
                    <RANKING order="2" place="2" resultid="11973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1255" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13963" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13964" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13965" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13966" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13967" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13968" daytime="10:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13969" daytime="10:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13970" daytime="10:20" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1381" daytime="11:45" gender="M" number="17" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1382" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1383" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10361" />
                    <RANKING order="2" place="2" resultid="10548" />
                    <RANKING order="3" place="3" resultid="10995" />
                    <RANKING order="4" place="4" resultid="12375" />
                    <RANKING order="5" place="5" resultid="10162" />
                    <RANKING order="6" place="6" resultid="10693" />
                    <RANKING order="7" place="-1" resultid="11346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1384" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10360" />
                    <RANKING order="2" place="2" resultid="11631" />
                    <RANKING order="3" place="3" resultid="11910" />
                    <RANKING order="4" place="4" resultid="12285" />
                    <RANKING order="5" place="5" resultid="11482" />
                    <RANKING order="6" place="6" resultid="9701" />
                    <RANKING order="7" place="7" resultid="10550" />
                    <RANKING order="8" place="-1" resultid="9561" />
                    <RANKING order="9" place="-1" resultid="11911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11347" />
                    <RANKING order="2" place="2" resultid="12160" />
                    <RANKING order="3" place="3" resultid="12220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9563" />
                    <RANKING order="2" place="2" resultid="10828" />
                    <RANKING order="3" place="3" resultid="10552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11483" />
                    <RANKING order="2" place="2" resultid="10062" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13997" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13998" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13999" daytime="11:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:25" gender="F" number="12" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10422" />
                    <RANKING order="2" place="2" resultid="11802" />
                    <RANKING order="3" place="3" resultid="11089" />
                    <RANKING order="4" place="4" resultid="10140" />
                    <RANKING order="5" place="5" resultid="10500" />
                    <RANKING order="6" place="6" resultid="9986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12103" />
                    <RANKING order="2" place="2" resultid="10128" />
                    <RANKING order="3" place="3" resultid="11677" />
                    <RANKING order="4" place="4" resultid="12768" />
                    <RANKING order="5" place="5" resultid="12254" />
                    <RANKING order="6" place="6" resultid="9836" />
                    <RANKING order="7" place="-1" resultid="12177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12761" />
                    <RANKING order="2" place="2" resultid="12377" />
                    <RANKING order="3" place="3" resultid="12357" />
                    <RANKING order="4" place="4" resultid="11667" />
                    <RANKING order="5" place="5" resultid="10155" />
                    <RANKING order="6" place="6" resultid="10306" />
                    <RANKING order="7" place="7" resultid="11745" />
                    <RANKING order="8" place="8" resultid="10344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12428" />
                    <RANKING order="2" place="2" resultid="10087" />
                    <RANKING order="3" place="3" resultid="11838" />
                    <RANKING order="4" place="4" resultid="12438" />
                    <RANKING order="5" place="5" resultid="10258" />
                    <RANKING order="6" place="6" resultid="11736" />
                    <RANKING order="7" place="7" resultid="9657" />
                    <RANKING order="8" place="-1" resultid="10462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9556" />
                    <RANKING order="2" place="2" resultid="11516" />
                    <RANKING order="3" place="3" resultid="11729" />
                    <RANKING order="4" place="4" resultid="11948" />
                    <RANKING order="5" place="5" resultid="12240" />
                    <RANKING order="6" place="6" resultid="10101" />
                    <RANKING order="7" place="7" resultid="10456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11338" />
                    <RANKING order="2" place="2" resultid="11390" />
                    <RANKING order="3" place="3" resultid="12233" />
                    <RANKING order="4" place="4" resultid="10776" />
                    <RANKING order="5" place="5" resultid="11939" />
                    <RANKING order="6" place="-1" resultid="12081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11395" />
                    <RANKING order="2" place="2" resultid="10907" />
                    <RANKING order="3" place="3" resultid="9514" />
                    <RANKING order="4" place="4" resultid="11293" />
                    <RANKING order="5" place="5" resultid="9842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11460" />
                    <RANKING order="2" place="2" resultid="12097" />
                    <RANKING order="3" place="3" resultid="12248" />
                    <RANKING order="4" place="4" resultid="9673" />
                    <RANKING order="5" place="5" resultid="10470" />
                    <RANKING order="6" place="-1" resultid="9970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9500" />
                    <RANKING order="2" place="2" resultid="10409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12126" />
                    <RANKING order="2" place="2" resultid="10291" />
                    <RANKING order="3" place="-1" resultid="10334" />
                    <RANKING order="4" place="-1" resultid="10725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1269" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1270" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1271" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1272" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13971" daytime="10:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13972" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13973" daytime="10:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13974" daytime="10:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13975" daytime="10:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13976" daytime="10:40" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="11:40" gender="F" number="16" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1375" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11908" />
                    <RANKING order="2" place="2" resultid="10362" />
                    <RANKING order="3" place="3" resultid="10553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9569" />
                    <RANKING order="2" place="2" resultid="12287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11481" />
                    <RANKING order="2" place="2" resultid="11348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1380" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13996" daytime="11:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="09:10" gender="M" number="9" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11638" />
                    <RANKING order="2" place="2" resultid="12466" />
                    <RANKING order="3" place="3" resultid="11096" />
                    <RANKING order="4" place="4" resultid="10942" />
                    <RANKING order="5" place="5" resultid="10447" />
                    <RANKING order="6" place="6" resultid="11692" />
                    <RANKING order="7" place="-1" resultid="9732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10476" />
                    <RANKING order="2" place="2" resultid="12451" />
                    <RANKING order="3" place="3" resultid="12076" />
                    <RANKING order="4" place="4" resultid="10924" />
                    <RANKING order="5" place="5" resultid="10781" />
                    <RANKING order="6" place="6" resultid="9617" />
                    <RANKING order="7" place="-1" resultid="10689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12797" />
                    <RANKING order="2" place="2" resultid="10989" />
                    <RANKING order="3" place="3" resultid="12788" />
                    <RANKING order="4" place="4" resultid="12167" />
                    <RANKING order="5" place="5" resultid="10213" />
                    <RANKING order="6" place="-1" resultid="12343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11651" />
                    <RANKING order="2" place="2" resultid="10348" />
                    <RANKING order="3" place="3" resultid="11319" />
                    <RANKING order="4" place="4" resultid="9523" />
                    <RANKING order="5" place="5" resultid="11075" />
                    <RANKING order="6" place="6" resultid="11759" />
                    <RANKING order="7" place="7" resultid="12337" />
                    <RANKING order="8" place="8" resultid="12369" />
                    <RANKING order="9" place="9" resultid="10679" />
                    <RANKING order="10" place="10" resultid="12351" />
                    <RANKING order="11" place="11" resultid="11435" />
                    <RANKING order="12" place="12" resultid="10441" />
                    <RANKING order="13" place="-1" resultid="9688" />
                    <RANKING order="14" place="-1" resultid="10950" />
                    <RANKING order="15" place="-1" resultid="10970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11536" />
                    <RANKING order="2" place="2" resultid="11593" />
                    <RANKING order="3" place="3" resultid="11523" />
                    <RANKING order="4" place="4" resultid="11625" />
                    <RANKING order="5" place="5" resultid="11849" />
                    <RANKING order="6" place="6" resultid="9519" />
                    <RANKING order="7" place="7" resultid="11866" />
                    <RANKING order="8" place="8" resultid="9426" />
                    <RANKING order="9" place="9" resultid="11858" />
                    <RANKING order="10" place="10" resultid="10684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12302" />
                    <RANKING order="2" place="2" resultid="11701" />
                    <RANKING order="3" place="3" resultid="12266" />
                    <RANKING order="4" place="4" resultid="9907" />
                    <RANKING order="5" place="5" resultid="11601" />
                    <RANKING order="6" place="6" resultid="11901" />
                    <RANKING order="7" place="7" resultid="12214" />
                    <RANKING order="8" place="8" resultid="10271" />
                    <RANKING order="9" place="9" resultid="10436" />
                    <RANKING order="10" place="10" resultid="12199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11014" />
                    <RANKING order="2" place="2" resultid="11280" />
                    <RANKING order="3" place="3" resultid="9829" />
                    <RANKING order="4" place="4" resultid="10222" />
                    <RANKING order="5" place="5" resultid="11401" />
                    <RANKING order="6" place="6" resultid="10797" />
                    <RANKING order="7" place="7" resultid="9680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9491" />
                    <RANKING order="2" place="2" resultid="11609" />
                    <RANKING order="3" place="3" resultid="10894" />
                    <RANKING order="4" place="4" resultid="11045" />
                    <RANKING order="5" place="5" resultid="9753" />
                    <RANKING order="6" place="6" resultid="10720" />
                    <RANKING order="7" place="7" resultid="12108" />
                    <RANKING order="8" place="8" resultid="10237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9771" />
                    <RANKING order="2" place="2" resultid="9650" />
                    <RANKING order="3" place="3" resultid="9409" />
                    <RANKING order="4" place="4" resultid="11955" />
                    <RANKING order="5" place="5" resultid="9939" />
                    <RANKING order="6" place="6" resultid="12139" />
                    <RANKING order="7" place="7" resultid="9696" />
                    <RANKING order="8" place="8" resultid="9865" />
                    <RANKING order="9" place="9" resultid="9764" />
                    <RANKING order="10" place="10" resultid="10051" />
                    <RANKING order="11" place="11" resultid="9474" />
                    <RANKING order="12" place="12" resultid="10506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10251" />
                    <RANKING order="2" place="2" resultid="12133" />
                    <RANKING order="3" place="3" resultid="12418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10184" />
                    <RANKING order="2" place="2" resultid="9400" />
                    <RANKING order="3" place="3" resultid="10009" />
                    <RANKING order="4" place="4" resultid="12207" />
                    <RANKING order="5" place="5" resultid="11378" />
                    <RANKING order="6" place="6" resultid="9889" />
                    <RANKING order="7" place="7" resultid="11444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9977" />
                    <RANKING order="2" place="2" resultid="11972" />
                    <RANKING order="3" place="3" resultid="9880" />
                    <RANKING order="4" place="4" resultid="9872" />
                    <RANKING order="5" place="-1" resultid="11018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1221" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13949" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13950" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13951" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13952" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13953" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13954" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13955" daytime="09:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13956" daytime="09:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="13957" daytime="09:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="13958" daytime="09:25" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="10:40" gender="M" number="13" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10943" />
                    <RANKING order="2" place="2" resultid="12171" />
                    <RANKING order="3" place="3" resultid="10448" />
                    <RANKING order="4" place="4" resultid="11693" />
                    <RANKING order="5" place="-1" resultid="12401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12444" />
                    <RANKING order="2" place="2" resultid="9536" />
                    <RANKING order="3" place="3" resultid="10875" />
                    <RANKING order="4" place="4" resultid="12183" />
                    <RANKING order="5" place="5" resultid="10492" />
                    <RANKING order="6" place="6" resultid="12452" />
                    <RANKING order="7" place="7" resultid="12077" />
                    <RANKING order="8" place="8" resultid="10108" />
                    <RANKING order="9" place="9" resultid="10690" />
                    <RANKING order="10" place="10" resultid="10786" />
                    <RANKING order="11" place="11" resultid="12333" />
                    <RANKING order="12" place="12" resultid="9618" />
                    <RANKING order="13" place="-1" resultid="10296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11998" />
                    <RANKING order="2" place="2" resultid="10355" />
                    <RANKING order="3" place="3" resultid="12782" />
                    <RANKING order="4" place="4" resultid="10148" />
                    <RANKING order="5" place="5" resultid="12789" />
                    <RANKING order="6" place="6" resultid="11430" />
                    <RANKING order="7" place="7" resultid="12189" />
                    <RANKING order="8" place="8" resultid="12344" />
                    <RANKING order="9" place="9" resultid="10121" />
                    <RANKING order="10" place="10" resultid="10214" />
                    <RANKING order="11" place="11" resultid="9919" />
                    <RANKING order="12" place="-1" resultid="10032" />
                    <RANKING order="13" place="-1" resultid="11711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9608" />
                    <RANKING order="2" place="2" resultid="12370" />
                    <RANKING order="3" place="3" resultid="10537" />
                    <RANKING order="4" place="4" resultid="10962" />
                    <RANKING order="5" place="5" resultid="12352" />
                    <RANKING order="6" place="6" resultid="11332" />
                    <RANKING order="7" place="7" resultid="10201" />
                    <RANKING order="8" place="8" resultid="11760" />
                    <RANKING order="9" place="9" resultid="10977" />
                    <RANKING order="10" place="10" resultid="9859" />
                    <RANKING order="11" place="11" resultid="12273" />
                    <RANKING order="12" place="12" resultid="12085" />
                    <RANKING order="13" place="13" resultid="10442" />
                    <RANKING order="14" place="14" resultid="11436" />
                    <RANKING order="15" place="-1" resultid="11314" />
                    <RANKING order="16" place="-1" resultid="11720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11537" />
                    <RANKING order="2" place="2" resultid="11626" />
                    <RANKING order="3" place="3" resultid="12317" />
                    <RANKING order="4" place="4" resultid="11850" />
                    <RANKING order="5" place="5" resultid="10673" />
                    <RANKING order="6" place="6" resultid="11594" />
                    <RANKING order="7" place="7" resultid="11867" />
                    <RANKING order="8" place="8" resultid="10328" />
                    <RANKING order="9" place="9" resultid="11549" />
                    <RANKING order="10" place="10" resultid="11425" />
                    <RANKING order="11" place="11" resultid="12278" />
                    <RANKING order="12" place="12" resultid="10685" />
                    <RANKING order="13" place="13" resultid="11877" />
                    <RANKING order="14" place="14" resultid="10116" />
                    <RANKING order="15" place="15" resultid="10761" />
                    <RANKING order="16" place="16" resultid="9747" />
                    <RANKING order="17" place="-1" resultid="10983" />
                    <RANKING order="18" place="-1" resultid="11883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10179" />
                    <RANKING order="2" place="2" resultid="11702" />
                    <RANKING order="3" place="3" resultid="11685" />
                    <RANKING order="4" place="4" resultid="11057" />
                    <RANKING order="5" place="5" resultid="10429" />
                    <RANKING order="6" place="6" resultid="10870" />
                    <RANKING order="7" place="7" resultid="12756" />
                    <RANKING order="8" place="8" resultid="11172" />
                    <RANKING order="9" place="9" resultid="11177" />
                    <RANKING order="10" place="10" resultid="10529" />
                    <RANKING order="11" place="11" resultid="12200" />
                    <RANKING order="12" place="12" resultid="12215" />
                    <RANKING order="13" place="13" resultid="12448" />
                    <RANKING order="14" place="14" resultid="10754" />
                    <RANKING order="15" place="-1" resultid="10272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10230" />
                    <RANKING order="2" place="2" resultid="11015" />
                    <RANKING order="3" place="3" resultid="11342" />
                    <RANKING order="4" place="4" resultid="10223" />
                    <RANKING order="5" place="5" resultid="9715" />
                    <RANKING order="6" place="6" resultid="12114" />
                    <RANKING order="7" place="7" resultid="11964" />
                    <RANKING order="8" place="8" resultid="12325" />
                    <RANKING order="9" place="9" resultid="9899" />
                    <RANKING order="10" place="10" resultid="9681" />
                    <RANKING order="11" place="11" resultid="10798" />
                    <RANKING order="12" place="12" resultid="10792" />
                    <RANKING order="13" place="13" resultid="10804" />
                    <RANKING order="14" place="-1" resultid="9830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10191" />
                    <RANKING order="2" place="2" resultid="11556" />
                    <RANKING order="3" place="3" resultid="11610" />
                    <RANKING order="4" place="4" resultid="12458" />
                    <RANKING order="5" place="5" resultid="9622" />
                    <RANKING order="6" place="6" resultid="10238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10207" />
                    <RANKING order="2" place="2" resultid="9602" />
                    <RANKING order="3" place="3" resultid="11008" />
                    <RANKING order="4" place="4" resultid="9410" />
                    <RANKING order="5" place="5" resultid="10017" />
                    <RANKING order="6" place="6" resultid="9697" />
                    <RANKING order="7" place="7" resultid="9940" />
                    <RANKING order="8" place="8" resultid="9475" />
                    <RANKING order="9" place="9" resultid="10507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10252" />
                    <RANKING order="2" place="2" resultid="11409" />
                    <RANKING order="3" place="3" resultid="10816" />
                    <RANKING order="4" place="4" resultid="9351" />
                    <RANKING order="5" place="5" resultid="12065" />
                    <RANKING order="6" place="6" resultid="10542" />
                    <RANKING order="7" place="-1" resultid="9529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9595" />
                    <RANKING order="2" place="2" resultid="10185" />
                    <RANKING order="3" place="3" resultid="9401" />
                    <RANKING order="4" place="4" resultid="11445" />
                    <RANKING order="5" place="5" resultid="9890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9357" />
                    <RANKING order="2" place="2" resultid="9978" />
                    <RANKING order="3" place="3" resultid="11384" />
                    <RANKING order="4" place="4" resultid="9873" />
                    <RANKING order="5" place="-1" resultid="9993" />
                    <RANKING order="6" place="-1" resultid="11019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10514" />
                    <RANKING order="2" place="2" resultid="12390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1289" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13977" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13978" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13979" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13980" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13981" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13982" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13983" daytime="10:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13984" daytime="11:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="13985" daytime="11:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="13986" daytime="11:00" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="13987" daytime="11:05" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="13988" daytime="11:05" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="13989" daytime="11:10" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-06-11" daytime="16:00" endtime="20:21" name="BLOK III" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1508" daytime="17:50" gender="M" number="25" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1509" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12469" />
                    <RANKING order="2" place="2" resultid="12173" />
                    <RANKING order="3" place="3" resultid="9430" />
                    <RANKING order="4" place="4" resultid="10945" />
                    <RANKING order="5" place="5" resultid="10450" />
                    <RANKING order="6" place="6" resultid="11695" />
                    <RANKING order="7" place="7" resultid="10881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9538" />
                    <RANKING order="2" place="2" resultid="12411" />
                    <RANKING order="3" place="3" resultid="12185" />
                    <RANKING order="4" place="4" resultid="10876" />
                    <RANKING order="5" place="5" resultid="10197" />
                    <RANKING order="6" place="6" resultid="10111" />
                    <RANKING order="7" place="7" resultid="12461" />
                    <RANKING order="8" place="-1" resultid="10494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10356" />
                    <RANKING order="2" place="2" resultid="11713" />
                    <RANKING order="3" place="3" resultid="12791" />
                    <RANKING order="4" place="4" resultid="10034" />
                    <RANKING order="5" place="5" resultid="10216" />
                    <RANKING order="6" place="6" resultid="9920" />
                    <RANKING order="7" place="-1" resultid="12346" />
                    <RANKING order="8" place="-1" resultid="10993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11302" />
                    <RANKING order="2" place="2" resultid="10964" />
                    <RANKING order="3" place="3" resultid="10203" />
                    <RANKING order="4" place="4" resultid="10538" />
                    <RANKING order="5" place="5" resultid="12354" />
                    <RANKING order="6" place="6" resultid="12372" />
                    <RANKING order="7" place="7" resultid="10040" />
                    <RANKING order="8" place="-1" resultid="11321" />
                    <RANKING order="9" place="-1" resultid="12275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12319" />
                    <RANKING order="2" place="2" resultid="11852" />
                    <RANKING order="3" place="3" resultid="11083" />
                    <RANKING order="4" place="4" resultid="10330" />
                    <RANKING order="5" place="5" resultid="11550" />
                    <RANKING order="6" place="6" resultid="11869" />
                    <RANKING order="7" place="7" resultid="11879" />
                    <RANKING order="8" place="8" resultid="12262" />
                    <RANKING order="9" place="9" resultid="10117" />
                    <RANKING order="10" place="10" resultid="9748" />
                    <RANKING order="11" place="11" resultid="11577" />
                    <RANKING order="12" place="-1" resultid="10675" />
                    <RANKING order="13" place="-1" resultid="11580" />
                    <RANKING order="14" place="-1" resultid="12280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10180" />
                    <RANKING order="2" place="2" resultid="11686" />
                    <RANKING order="3" place="3" resultid="10872" />
                    <RANKING order="4" place="4" resultid="10900" />
                    <RANKING order="5" place="5" resultid="10531" />
                    <RANKING order="6" place="-1" resultid="9423" />
                    <RANKING order="7" place="-1" resultid="10274" />
                    <RANKING order="8" place="-1" resultid="12202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10225" />
                    <RANKING order="2" place="2" resultid="11343" />
                    <RANKING order="3" place="3" resultid="9717" />
                    <RANKING order="4" place="4" resultid="12157" />
                    <RANKING order="5" place="5" resultid="12327" />
                    <RANKING order="6" place="6" resultid="11967" />
                    <RANKING order="7" place="7" resultid="11274" />
                    <RANKING order="8" place="8" resultid="10800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10192" />
                    <RANKING order="2" place="2" resultid="11557" />
                    <RANKING order="3" place="3" resultid="12459" />
                    <RANKING order="4" place="4" resultid="9623" />
                    <RANKING order="5" place="5" resultid="10239" />
                    <RANKING order="6" place="-1" resultid="9494" />
                    <RANKING order="7" place="-1" resultid="11048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9604" />
                    <RANKING order="2" place="2" resultid="9724" />
                    <RANKING order="3" place="3" resultid="11114" />
                    <RANKING order="4" place="4" resultid="10019" />
                    <RANKING order="5" place="5" resultid="9412" />
                    <RANKING order="6" place="6" resultid="11958" />
                    <RANKING order="7" place="7" resultid="9477" />
                    <RANKING order="8" place="-1" resultid="9942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10254" />
                    <RANKING order="2" place="2" resultid="10817" />
                    <RANKING order="3" place="3" resultid="11411" />
                    <RANKING order="4" place="4" resultid="9352" />
                    <RANKING order="5" place="5" resultid="10003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9418" />
                    <RANKING order="2" place="2" resultid="9597" />
                    <RANKING order="3" place="3" resultid="10187" />
                    <RANKING order="4" place="4" resultid="11447" />
                    <RANKING order="5" place="5" resultid="9892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9358" />
                    <RANKING order="2" place="2" resultid="11385" />
                    <RANKING order="3" place="3" resultid="9875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1522" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10515" />
                    <RANKING order="2" place="2" resultid="12392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1524" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14044" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14045" daytime="18:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14046" daytime="18:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14047" daytime="18:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14048" daytime="18:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14049" daytime="18:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14050" daytime="18:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14051" daytime="18:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14052" daytime="18:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14053" daytime="18:30" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1474" daytime="17:10" gender="M" number="23" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1475" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11099" />
                    <RANKING order="2" place="2" resultid="9429" />
                    <RANKING order="3" place="3" resultid="9735" />
                    <RANKING order="4" place="-1" resultid="12402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10477" />
                    <RANKING order="2" place="2" resultid="12454" />
                    <RANKING order="3" place="3" resultid="10782" />
                    <RANKING order="4" place="4" resultid="10927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12800" />
                    <RANKING order="2" place="2" resultid="11742" />
                    <RANKING order="3" place="3" resultid="10992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11653" />
                    <RANKING order="2" place="2" resultid="11320" />
                    <RANKING order="3" place="3" resultid="9524" />
                    <RANKING order="4" place="4" resultid="12338" />
                    <RANKING order="5" place="5" resultid="11762" />
                    <RANKING order="6" place="6" resultid="10681" />
                    <RANKING order="7" place="-1" resultid="9690" />
                    <RANKING order="8" place="-1" resultid="10443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11538" />
                    <RANKING order="2" place="2" resultid="11596" />
                    <RANKING order="3" place="3" resultid="10984" />
                    <RANKING order="4" place="-1" resultid="9520" />
                    <RANKING order="5" place="-1" resultid="11525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12303" />
                    <RANKING order="2" place="2" resultid="11704" />
                    <RANKING order="3" place="3" resultid="9909" />
                    <RANKING order="4" place="4" resultid="12268" />
                    <RANKING order="5" place="5" resultid="12217" />
                    <RANKING order="6" place="6" resultid="10437" />
                    <RANKING order="7" place="-1" resultid="12757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10224" />
                    <RANKING order="2" place="2" resultid="11281" />
                    <RANKING order="3" place="3" resultid="11966" />
                    <RANKING order="4" place="4" resultid="11403" />
                    <RANKING order="5" place="5" resultid="10799" />
                    <RANKING order="6" place="6" resultid="9683" />
                    <RANKING order="7" place="7" resultid="10794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11925" />
                    <RANKING order="2" place="2" resultid="11611" />
                    <RANKING order="3" place="3" resultid="10895" />
                    <RANKING order="4" place="4" resultid="11047" />
                    <RANKING order="5" place="5" resultid="10721" />
                    <RANKING order="6" place="6" resultid="11809" />
                    <RANKING order="7" place="-1" resultid="9755" />
                    <RANKING order="8" place="-1" resultid="10737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10208" />
                    <RANKING order="2" place="2" resultid="9772" />
                    <RANKING order="3" place="3" resultid="12141" />
                    <RANKING order="4" place="4" resultid="9698" />
                    <RANKING order="5" place="5" resultid="9941" />
                    <RANKING order="6" place="6" resultid="10508" />
                    <RANKING order="7" place="7" resultid="9476" />
                    <RANKING order="8" place="-1" resultid="9867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10253" />
                    <RANKING order="2" place="2" resultid="12134" />
                    <RANKING order="3" place="3" resultid="12067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10186" />
                    <RANKING order="2" place="2" resultid="9403" />
                    <RANKING order="3" place="3" resultid="11379" />
                    <RANKING order="4" place="4" resultid="10012" />
                    <RANKING order="5" place="5" resultid="12209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11975" />
                    <RANKING order="2" place="2" resultid="9994" />
                    <RANKING order="3" place="3" resultid="9874" />
                    <RANKING order="4" place="-1" resultid="11020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1489" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1490" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14032" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14033" daytime="17:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14034" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14035" daytime="17:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14036" daytime="17:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14037" daytime="17:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14038" daytime="17:30" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1548" daytime="18:40" gender="M" number="27" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1549" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1550" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10363" />
                    <RANKING order="2" place="2" resultid="10163" />
                    <RANKING order="3" place="3" resultid="10996" />
                    <RANKING order="4" place="4" resultid="10366" />
                    <RANKING order="5" place="-1" resultid="10549" />
                    <RANKING order="6" place="-1" resultid="10692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12376" />
                    <RANKING order="2" place="2" resultid="11912" />
                    <RANKING order="3" place="3" resultid="12286" />
                    <RANKING order="4" place="4" resultid="9702" />
                    <RANKING order="5" place="5" resultid="10551" />
                    <RANKING order="6" place="-1" resultid="9562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9564" />
                    <RANKING order="2" place="2" resultid="11485" />
                    <RANKING order="3" place="3" resultid="10827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10063" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14055" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14056" daytime="18:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="17:00" gender="F" number="22" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1458" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10936" />
                    <RANKING order="2" place="-1" resultid="10136" />
                    <RANKING order="3" place="-1" resultid="11804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11678" />
                    <RANKING order="2" place="2" resultid="10402" />
                    <RANKING order="3" place="3" resultid="12255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11659" />
                    <RANKING order="2" place="2" resultid="10522" />
                    <RANKING order="3" place="3" resultid="9631" />
                    <RANKING order="4" place="4" resultid="11932" />
                    <RANKING order="5" place="-1" resultid="11533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10082" />
                    <RANKING order="2" place="2" resultid="11831" />
                    <RANKING order="3" place="3" resultid="10259" />
                    <RANKING order="4" place="4" resultid="11738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9558" />
                    <RANKING order="2" place="2" resultid="11731" />
                    <RANKING order="3" place="3" resultid="10457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10904" />
                    <RANKING order="2" place="2" resultid="12307" />
                    <RANKING order="3" place="3" resultid="10418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9509" />
                    <RANKING order="2" place="2" resultid="11294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11107" />
                    <RANKING order="2" place="2" resultid="11053" />
                    <RANKING order="3" place="3" resultid="11470" />
                    <RANKING order="4" place="4" resultid="9674" />
                    <RANKING order="5" place="5" resultid="10472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9963" />
                    <RANKING order="2" place="2" resultid="10411" />
                    <RANKING order="3" place="3" resultid="9854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10292" />
                    <RANKING order="2" place="2" resultid="9952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1469" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1471" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1472" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1473" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14028" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14029" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14030" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14031" daytime="17:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="16:15" gender="M" number="19" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1407" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12363" />
                    <RANKING order="2" place="2" resultid="12468" />
                    <RANKING order="3" place="3" resultid="10944" />
                    <RANKING order="4" place="4" resultid="10449" />
                    <RANKING order="5" place="5" resultid="11098" />
                    <RANKING order="6" place="-1" resultid="9734" />
                    <RANKING order="7" place="-1" resultid="11640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12410" />
                    <RANKING order="2" place="2" resultid="11475" />
                    <RANKING order="3" place="3" resultid="10196" />
                    <RANKING order="4" place="4" resultid="10787" />
                    <RANKING order="5" place="5" resultid="10926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10352" />
                    <RANKING order="2" place="2" resultid="10033" />
                    <RANKING order="3" place="3" resultid="12783" />
                    <RANKING order="4" place="4" resultid="10304" />
                    <RANKING order="5" place="5" resultid="12073" />
                    <RANKING order="6" place="-1" resultid="10991" />
                    <RANKING order="7" place="-1" resultid="12473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11333" />
                    <RANKING order="2" place="2" resultid="10282" />
                    <RANKING order="3" place="3" resultid="10956" />
                    <RANKING order="4" place="4" resultid="11722" />
                    <RANKING order="5" place="5" resultid="12086" />
                    <RANKING order="6" place="-1" resultid="10972" />
                    <RANKING order="7" place="-1" resultid="11077" />
                    <RANKING order="8" place="-1" resultid="11620" />
                    <RANKING order="9" place="-1" resultid="11994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11627" />
                    <RANKING order="2" place="2" resultid="11860" />
                    <RANKING order="3" place="3" resultid="11451" />
                    <RANKING order="4" place="4" resultid="10329" />
                    <RANKING order="5" place="5" resultid="10078" />
                    <RANKING order="6" place="6" resultid="12261" />
                    <RANKING order="7" place="7" resultid="10391" />
                    <RANKING order="8" place="-1" resultid="10674" />
                    <RANKING order="9" place="-1" resultid="11529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10899" />
                    <RANKING order="2" place="2" resultid="9741" />
                    <RANKING order="3" place="3" resultid="10430" />
                    <RANKING order="4" place="4" resultid="11896" />
                    <RANKING order="5" place="5" resultid="11509" />
                    <RANKING order="6" place="6" resultid="9761" />
                    <RANKING order="7" place="7" resultid="11902" />
                    <RANKING order="8" place="8" resultid="10074" />
                    <RANKING order="9" place="9" resultid="11178" />
                    <RANKING order="10" place="10" resultid="10871" />
                    <RANKING order="11" place="11" resultid="9394" />
                    <RANKING order="12" place="12" resultid="10273" />
                    <RANKING order="13" place="13" resultid="10755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10231" />
                    <RANKING order="2" place="2" resultid="12156" />
                    <RANKING order="3" place="3" resultid="12115" />
                    <RANKING order="4" place="4" resultid="11326" />
                    <RANKING order="5" place="5" resultid="9682" />
                    <RANKING order="6" place="6" resultid="10397" />
                    <RANKING order="7" place="7" resultid="10793" />
                    <RANKING order="8" place="8" resultid="10265" />
                    <RANKING order="9" place="-1" resultid="9549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11981" />
                    <RANKING order="2" place="2" resultid="12149" />
                    <RANKING order="3" place="3" resultid="12109" />
                    <RANKING order="4" place="4" resultid="9486" />
                    <RANKING order="5" place="5" resultid="11365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12195" />
                    <RANKING order="2" place="2" resultid="9946" />
                    <RANKING order="3" place="3" resultid="11031" />
                    <RANKING order="4" place="4" resultid="11574" />
                    <RANKING order="5" place="5" resultid="11818" />
                    <RANKING order="6" place="6" resultid="9411" />
                    <RANKING order="7" place="7" resultid="10052" />
                    <RANKING order="8" place="8" resultid="10812" />
                    <RANKING order="9" place="9" resultid="9766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9482" />
                    <RANKING order="2" place="2" resultid="12420" />
                    <RANKING order="3" place="3" resultid="12066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12208" />
                    <RANKING order="2" place="2" resultid="10011" />
                    <RANKING order="3" place="3" resultid="9891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10704" />
                    <RANKING order="2" place="2" resultid="9979" />
                    <RANKING order="3" place="3" resultid="11974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1422" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14005" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14006" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14007" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14008" daytime="16:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14009" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14010" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14011" daytime="16:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14012" daytime="16:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14013" daytime="16:35" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="17:30" gender="F" number="24" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10424" />
                    <RANKING order="2" place="2" resultid="11091" />
                    <RANKING order="3" place="3" resultid="10918" />
                    <RANKING order="4" place="4" resultid="10502" />
                    <RANKING order="5" place="5" resultid="10486" />
                    <RANKING order="6" place="6" resultid="9987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10095" />
                    <RANKING order="2" place="2" resultid="11679" />
                    <RANKING order="3" place="3" resultid="12770" />
                    <RANKING order="4" place="4" resultid="9837" />
                    <RANKING order="5" place="-1" resultid="10130" />
                    <RANKING order="6" place="-1" resultid="11844" />
                    <RANKING order="7" place="-1" resultid="12105" />
                    <RANKING order="8" place="-1" resultid="12178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12763" />
                    <RANKING order="2" place="2" resultid="11660" />
                    <RANKING order="3" place="3" resultid="10523" />
                    <RANKING order="4" place="4" resultid="11670" />
                    <RANKING order="5" place="5" resultid="12777" />
                    <RANKING order="6" place="6" resultid="10308" />
                    <RANKING order="7" place="7" resultid="11747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10088" />
                    <RANKING order="2" place="2" resultid="11832" />
                    <RANKING order="3" place="3" resultid="11840" />
                    <RANKING order="4" place="4" resultid="10260" />
                    <RANKING order="5" place="5" resultid="9659" />
                    <RANKING order="6" place="-1" resultid="10464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10732" />
                    <RANKING order="2" place="2" resultid="11518" />
                    <RANKING order="3" place="3" resultid="10102" />
                    <RANKING order="4" place="4" resultid="11949" />
                    <RANKING order="5" place="5" resultid="12242" />
                    <RANKING order="6" place="-1" resultid="11824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11339" />
                    <RANKING order="2" place="2" resultid="12235" />
                    <RANKING order="3" place="3" resultid="11941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10909" />
                    <RANKING order="2" place="2" resultid="10245" />
                    <RANKING order="3" place="-1" resultid="9844" />
                    <RANKING order="4" place="-1" resultid="9516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11463" />
                    <RANKING order="2" place="2" resultid="9675" />
                    <RANKING order="3" place="3" resultid="12250" />
                    <RANKING order="4" place="-1" resultid="12098" />
                    <RANKING order="5" place="-1" resultid="9971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10335" />
                    <RANKING order="2" place="-1" resultid="10726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1504" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1505" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1506" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1507" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14039" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14040" daytime="17:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14041" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14042" daytime="17:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14043" daytime="17:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="18:35" gender="F" number="26" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1542" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1543" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11909" />
                    <RANKING order="2" place="2" resultid="10554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1544" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9570" />
                    <RANKING order="2" place="2" resultid="12288" />
                    <RANKING order="3" place="3" resultid="10364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1545" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1547" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14054" daytime="18:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="19:05" gender="M" number="29" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1579" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12397" />
                    <RANKING order="2" place="2" resultid="12364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11563" />
                    <RANKING order="2" place="2" resultid="10478" />
                    <RANKING order="3" place="-1" resultid="10298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11026" />
                    <RANKING order="2" place="2" resultid="11714" />
                    <RANKING order="3" place="3" resultid="10150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11303" />
                    <RANKING order="2" place="2" resultid="11723" />
                    <RANKING order="3" place="3" resultid="10041" />
                    <RANKING order="4" place="-1" resultid="11621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9614" />
                    <RANKING order="2" place="2" resultid="11880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9742" />
                    <RANKING order="2" place="2" resultid="11687" />
                    <RANKING order="3" place="3" resultid="11897" />
                    <RANKING order="4" place="4" resultid="10431" />
                    <RANKING order="5" place="5" resultid="11510" />
                    <RANKING order="6" place="6" resultid="9395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9832" />
                    <RANKING order="2" place="2" resultid="12328" />
                    <RANKING order="3" place="3" resultid="9901" />
                    <RANKING order="4" place="4" resultid="10266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11612" />
                    <RANKING order="2" place="2" resultid="9642" />
                    <RANKING order="3" place="3" resultid="9756" />
                    <RANKING order="4" place="4" resultid="11366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12142" />
                    <RANKING order="2" place="2" resultid="9725" />
                    <RANKING order="3" place="3" resultid="9868" />
                    <RANKING order="4" place="4" resultid="11115" />
                    <RANKING order="5" place="-1" resultid="9773" />
                    <RANKING order="6" place="-1" resultid="11813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11412" />
                    <RANKING order="2" place="2" resultid="10004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1592" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1593" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1594" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14059" daytime="19:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14060" daytime="19:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14061" daytime="19:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14062" daytime="19:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1388" daytime="16:00" gender="F" number="18" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10423" />
                    <RANKING order="2" place="2" resultid="9710" />
                    <RANKING order="3" place="3" resultid="10917" />
                    <RANKING order="4" place="4" resultid="10501" />
                    <RANKING order="5" place="5" resultid="10286" />
                    <RANKING order="6" place="-1" resultid="11803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10094" />
                    <RANKING order="2" place="2" resultid="10129" />
                    <RANKING order="3" place="3" resultid="12769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12762" />
                    <RANKING order="2" place="2" resultid="10025" />
                    <RANKING order="3" place="3" resultid="10278" />
                    <RANKING order="4" place="4" resultid="11746" />
                    <RANKING order="5" place="5" resultid="10156" />
                    <RANKING order="6" place="6" resultid="12776" />
                    <RANKING order="7" place="7" resultid="10313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12439" />
                    <RANKING order="2" place="2" resultid="11889" />
                    <RANKING order="3" place="3" resultid="9658" />
                    <RANKING order="4" place="4" resultid="11737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10731" />
                    <RANKING order="2" place="2" resultid="12241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9544" />
                    <RANKING order="2" place="2" resultid="9914" />
                    <RANKING order="3" place="3" resultid="12234" />
                    <RANKING order="4" place="4" resultid="11586" />
                    <RANKING order="5" place="5" resultid="11940" />
                    <RANKING order="6" place="-1" resultid="12082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11396" />
                    <RANKING order="2" place="2" resultid="10244" />
                    <RANKING order="3" place="3" resultid="9515" />
                    <RANKING order="4" place="4" resultid="10908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11469" />
                    <RANKING order="2" place="2" resultid="11287" />
                    <RANKING order="3" place="3" resultid="10764" />
                    <RANKING order="4" place="4" resultid="12249" />
                    <RANKING order="5" place="5" resultid="9665" />
                    <RANKING order="6" place="6" resultid="10471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12311" />
                    <RANKING order="2" place="2" resultid="11646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1402" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1404" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1405" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14000" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14001" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14002" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14003" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14004" daytime="16:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1555" daytime="18:45" gender="F" number="28" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1562" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10142" />
                    <RANKING order="2" place="2" resultid="10487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10886" />
                    <RANKING order="2" place="2" resultid="10403" />
                    <RANKING order="3" place="3" resultid="12256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10026" />
                    <RANKING order="2" place="2" resultid="11933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11069" />
                    <RANKING order="2" place="2" resultid="12431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1567" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11311" />
                    <RANKING order="2" place="2" resultid="9845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11108" />
                    <RANKING order="2" place="2" resultid="9666" />
                    <RANKING order="3" place="3" resultid="11373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1571" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1572" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1573" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1574" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1575" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1576" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1577" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14057" daytime="18:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14058" daytime="18:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1423" daytime="16:40" gender="F" number="20" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10141" />
                    <RANKING order="2" place="2" resultid="11090" />
                    <RANKING order="3" place="3" resultid="10935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12378" />
                    <RANKING order="2" place="2" resultid="12358" />
                    <RANKING order="3" place="3" resultid="11669" />
                    <RANKING order="4" place="4" resultid="10307" />
                    <RANKING order="5" place="-1" resultid="10345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11068" />
                    <RANKING order="2" place="2" resultid="12430" />
                    <RANKING order="3" place="3" resultid="12440" />
                    <RANKING order="4" place="4" resultid="11839" />
                    <RANKING order="5" place="5" resultid="11890" />
                    <RANKING order="6" place="-1" resultid="10463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9557" />
                    <RANKING order="2" place="2" resultid="11517" />
                    <RANKING order="3" place="3" resultid="11730" />
                    <RANKING order="4" place="4" resultid="10771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11391" />
                    <RANKING order="2" place="2" resultid="9545" />
                    <RANKING order="3" place="3" resultid="10777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11397" />
                    <RANKING order="2" place="2" resultid="9508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11462" />
                    <RANKING order="2" place="2" resultid="11288" />
                    <RANKING order="3" place="3" resultid="10765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9501" />
                    <RANKING order="2" place="2" resultid="9962" />
                    <RANKING order="3" place="-1" resultid="10410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1436" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1437" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1438" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1439" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14014" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14015" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14016" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14017" daytime="16:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1440" daytime="16:45" gender="M" number="21" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1441" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12172" />
                    <RANKING order="2" place="2" resultid="11694" />
                    <RANKING order="3" place="-1" resultid="11641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10297" />
                    <RANKING order="2" place="2" resultid="9537" />
                    <RANKING order="3" place="3" resultid="10891" />
                    <RANKING order="4" place="4" resultid="12445" />
                    <RANKING order="5" place="5" resultid="12453" />
                    <RANKING order="6" place="6" resultid="12078" />
                    <RANKING order="7" place="7" resultid="12184" />
                    <RANKING order="8" place="8" resultid="10110" />
                    <RANKING order="9" place="9" resultid="10788" />
                    <RANKING order="10" place="10" resultid="12334" />
                    <RANKING order="11" place="-1" resultid="10493" />
                    <RANKING order="12" place="-1" resultid="10691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12799" />
                    <RANKING order="2" place="2" resultid="12790" />
                    <RANKING order="3" place="3" resultid="11741" />
                    <RANKING order="4" place="4" resultid="10149" />
                    <RANKING order="5" place="5" resultid="12345" />
                    <RANKING order="6" place="6" resultid="12074" />
                    <RANKING order="7" place="7" resultid="10122" />
                    <RANKING order="8" place="-1" resultid="10215" />
                    <RANKING order="9" place="-1" resultid="11999" />
                    <RANKING order="10" place="-1" resultid="12190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11652" />
                    <RANKING order="2" place="2" resultid="9609" />
                    <RANKING order="3" place="3" resultid="11078" />
                    <RANKING order="4" place="4" resultid="10963" />
                    <RANKING order="5" place="5" resultid="12371" />
                    <RANKING order="6" place="6" resultid="10957" />
                    <RANKING order="7" place="7" resultid="11761" />
                    <RANKING order="8" place="8" resultid="12353" />
                    <RANKING order="9" place="9" resultid="9689" />
                    <RANKING order="10" place="10" resultid="11334" />
                    <RANKING order="11" place="11" resultid="9860" />
                    <RANKING order="12" place="12" resultid="10978" />
                    <RANKING order="13" place="13" resultid="10202" />
                    <RANKING order="14" place="14" resultid="12274" />
                    <RANKING order="15" place="15" resultid="12087" />
                    <RANKING order="16" place="-1" resultid="10349" />
                    <RANKING order="17" place="-1" resultid="11315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12318" />
                    <RANKING order="2" place="2" resultid="11628" />
                    <RANKING order="3" place="3" resultid="11851" />
                    <RANKING order="4" place="4" resultid="11524" />
                    <RANKING order="5" place="5" resultid="11595" />
                    <RANKING order="6" place="6" resultid="12279" />
                    <RANKING order="7" place="7" resultid="11426" />
                    <RANKING order="8" place="8" resultid="10714" />
                    <RANKING order="9" place="9" resultid="11868" />
                    <RANKING order="10" place="10" resultid="10686" />
                    <RANKING order="11" place="11" resultid="10742" />
                    <RANKING order="12" place="12" resultid="11884" />
                    <RANKING order="13" place="-1" resultid="11861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11703" />
                    <RANKING order="2" place="2" resultid="11058" />
                    <RANKING order="3" place="3" resultid="11173" />
                    <RANKING order="4" place="4" resultid="11603" />
                    <RANKING order="5" place="5" resultid="11179" />
                    <RANKING order="6" place="6" resultid="11872" />
                    <RANKING order="7" place="7" resultid="10530" />
                    <RANKING order="8" place="8" resultid="12201" />
                    <RANKING order="9" place="9" resultid="12216" />
                    <RANKING order="10" place="10" resultid="10756" />
                    <RANKING order="11" place="-1" resultid="12267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9831" />
                    <RANKING order="2" place="2" resultid="10232" />
                    <RANKING order="3" place="3" resultid="9716" />
                    <RANKING order="4" place="4" resultid="11402" />
                    <RANKING order="5" place="5" resultid="9900" />
                    <RANKING order="6" place="6" resultid="11273" />
                    <RANKING order="7" place="7" resultid="10805" />
                    <RANKING order="8" place="-1" resultid="9550" />
                    <RANKING order="9" place="-1" resultid="12116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9493" />
                    <RANKING order="2" place="2" resultid="9924" />
                    <RANKING order="3" place="3" resultid="12150" />
                    <RANKING order="4" place="4" resultid="9641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11957" />
                    <RANKING order="2" place="2" resultid="9603" />
                    <RANKING order="3" place="3" resultid="11009" />
                    <RANKING order="4" place="4" resultid="10018" />
                    <RANKING order="5" place="5" resultid="11819" />
                    <RANKING order="6" place="6" resultid="10053" />
                    <RANKING order="7" place="7" resultid="9767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9531" />
                    <RANKING order="2" place="2" resultid="12421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9596" />
                    <RANKING order="2" place="2" resultid="9402" />
                    <RANKING order="3" place="3" resultid="11446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1455" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1456" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14018" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14019" daytime="16:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14020" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14021" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14022" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14023" daytime="16:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14024" daytime="16:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14025" daytime="16:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14026" daytime="17:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14027" daytime="17:00" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-06-12" daytime="09:00" endtime="13:21" name="BLOK IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1613" daytime="09:10" gender="M" number="31" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1614" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9539" />
                    <RANKING order="2" place="2" resultid="10299" />
                    <RANKING order="3" place="3" resultid="10112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12801" />
                    <RANKING order="2" place="2" resultid="11715" />
                    <RANKING order="3" place="3" resultid="12792" />
                    <RANKING order="4" place="4" resultid="10123" />
                    <RANKING order="5" place="-1" resultid="12347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11304" />
                    <RANKING order="2" place="2" resultid="9610" />
                    <RANKING order="3" place="3" resultid="11724" />
                    <RANKING order="4" place="4" resultid="10042" />
                    <RANKING order="5" place="-1" resultid="11316" />
                    <RANKING order="6" place="-1" resultid="11335" />
                    <RANKING order="7" place="-1" resultid="12373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11629" />
                    <RANKING order="2" place="2" resultid="12320" />
                    <RANKING order="3" place="3" resultid="11853" />
                    <RANKING order="4" place="4" resultid="10715" />
                    <RANKING order="5" place="5" resultid="11870" />
                    <RANKING order="6" place="6" resultid="10743" />
                    <RANKING order="7" place="-1" resultid="10318" />
                    <RANKING order="8" place="-1" resultid="10985" />
                    <RANKING order="9" place="-1" resultid="11862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11705" />
                    <RANKING order="2" place="2" resultid="11059" />
                    <RANKING order="3" place="3" resultid="9396" />
                    <RANKING order="4" place="4" resultid="11511" />
                    <RANKING order="5" place="5" resultid="12203" />
                    <RANKING order="6" place="-1" resultid="11604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9718" />
                    <RANKING order="2" place="2" resultid="11404" />
                    <RANKING order="3" place="3" resultid="12158" />
                    <RANKING order="4" place="4" resultid="11968" />
                    <RANKING order="5" place="5" resultid="12329" />
                    <RANKING order="6" place="6" resultid="11275" />
                    <RANKING order="7" place="7" resultid="9902" />
                    <RANKING order="8" place="8" resultid="10267" />
                    <RANKING order="9" place="-1" resultid="10398" />
                    <RANKING order="10" place="-1" resultid="10806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9495" />
                    <RANKING order="2" place="2" resultid="9643" />
                    <RANKING order="3" place="3" resultid="12151" />
                    <RANKING order="4" place="4" resultid="9757" />
                    <RANKING order="5" place="5" resultid="11367" />
                    <RANKING order="6" place="6" resultid="10240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9726" />
                    <RANKING order="2" place="2" resultid="11010" />
                    <RANKING order="3" place="3" resultid="11959" />
                    <RANKING order="4" place="4" resultid="9869" />
                    <RANKING order="5" place="5" resultid="11116" />
                    <RANKING order="6" place="6" resultid="11820" />
                    <RANKING order="7" place="7" resultid="9768" />
                    <RANKING order="8" place="-1" resultid="10020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9532" />
                    <RANKING order="2" place="2" resultid="11413" />
                    <RANKING order="3" place="3" resultid="10005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1627" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1628" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1629" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14066" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14067" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14068" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14069" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14070" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14071" daytime="09:25" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1647" daytime="09:45" gender="M" number="33" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1648" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12404" />
                    <RANKING order="2" place="2" resultid="9431" />
                    <RANKING order="3" place="3" resultid="11100" />
                    <RANKING order="4" place="4" resultid="10451" />
                    <RANKING order="5" place="-1" resultid="9736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10479" />
                    <RANKING order="2" place="2" resultid="10783" />
                    <RANKING order="3" place="3" resultid="10928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12802" />
                    <RANKING order="2" place="-1" resultid="11027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11654" />
                    <RANKING order="2" place="2" resultid="11322" />
                    <RANKING order="3" place="3" resultid="9525" />
                    <RANKING order="4" place="4" resultid="12339" />
                    <RANKING order="5" place="5" resultid="10973" />
                    <RANKING order="6" place="6" resultid="11437" />
                    <RANKING order="7" place="-1" resultid="10745" />
                    <RANKING order="8" place="-1" resultid="11763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11597" />
                    <RANKING order="2" place="2" resultid="11084" />
                    <RANKING order="3" place="-1" resultid="11427" />
                    <RANKING order="4" place="-1" resultid="11452" />
                    <RANKING order="5" place="-1" resultid="11539" />
                    <RANKING order="6" place="-1" resultid="11551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12304" />
                    <RANKING order="2" place="2" resultid="9910" />
                    <RANKING order="3" place="3" resultid="12270" />
                    <RANKING order="4" place="4" resultid="11605" />
                    <RANKING order="5" place="-1" resultid="11706" />
                    <RANKING order="6" place="-1" resultid="12218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10226" />
                    <RANKING order="2" place="2" resultid="11282" />
                    <RANKING order="3" place="3" resultid="10801" />
                    <RANKING order="4" place="4" resultid="10795" />
                    <RANKING order="5" place="5" resultid="11276" />
                    <RANKING order="6" place="6" resultid="10809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11926" />
                    <RANKING order="2" place="2" resultid="11613" />
                    <RANKING order="3" place="3" resultid="10896" />
                    <RANKING order="4" place="4" resultid="11810" />
                    <RANKING order="5" place="-1" resultid="9758" />
                    <RANKING order="6" place="-1" resultid="10722" />
                    <RANKING order="7" place="-1" resultid="11049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10209" />
                    <RANKING order="2" place="2" resultid="9774" />
                    <RANKING order="3" place="3" resultid="12143" />
                    <RANKING order="4" place="4" resultid="9870" />
                    <RANKING order="5" place="5" resultid="9478" />
                    <RANKING order="6" place="6" resultid="10509" />
                    <RANKING order="7" place="-1" resultid="9651" />
                    <RANKING order="8" place="-1" resultid="9943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10255" />
                    <RANKING order="2" place="2" resultid="12135" />
                    <RANKING order="3" place="3" resultid="12068" />
                    <RANKING order="4" place="4" resultid="10006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10188" />
                    <RANKING order="2" place="2" resultid="9404" />
                    <RANKING order="3" place="3" resultid="11380" />
                    <RANKING order="4" place="4" resultid="9893" />
                    <RANKING order="5" place="-1" resultid="11448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11976" />
                    <RANKING order="2" place="2" resultid="9885" />
                    <RANKING order="3" place="3" resultid="9876" />
                    <RANKING order="4" place="-1" resultid="9995" />
                    <RANKING order="5" place="-1" resultid="11021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1661" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1662" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1663" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14076" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14077" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14078" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14079" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14080" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14081" daytime="10:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14082" daytime="10:15" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="09:00" gender="F" number="30" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1597" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10143" />
                    <RANKING order="2" place="2" resultid="11092" />
                    <RANKING order="3" place="3" resultid="10937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10887" />
                    <RANKING order="2" place="2" resultid="11845" />
                    <RANKING order="3" place="-1" resultid="12257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10027" />
                    <RANKING order="2" place="2" resultid="12359" />
                    <RANKING order="3" place="3" resultid="11934" />
                    <RANKING order="4" place="4" resultid="11671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11070" />
                    <RANKING order="2" place="2" resultid="12432" />
                    <RANKING order="3" place="3" resultid="11841" />
                    <RANKING order="4" place="-1" resultid="11891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9559" />
                    <RANKING order="2" place="2" resultid="11519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9546" />
                    <RANKING order="2" place="2" resultid="12308" />
                    <RANKING order="3" place="3" resultid="11588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9510" />
                    <RANKING order="2" place="2" resultid="9846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11464" />
                    <RANKING order="2" place="2" resultid="11374" />
                    <RANKING order="3" place="3" resultid="9667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10412" />
                    <RANKING order="2" place="2" resultid="9964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1610" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1611" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1612" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14063" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14064" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14065" daytime="09:05" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1630" daytime="09:25" gender="F" number="32" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1631" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10938" />
                    <RANKING order="2" place="2" resultid="10488" />
                    <RANKING order="3" place="-1" resultid="10137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11680" />
                    <RANKING order="2" place="2" resultid="10404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11661" />
                    <RANKING order="2" place="2" resultid="10524" />
                    <RANKING order="3" place="3" resultid="9632" />
                    <RANKING order="4" place="4" resultid="11935" />
                    <RANKING order="5" place="5" resultid="12778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11833" />
                    <RANKING order="2" place="2" resultid="10083" />
                    <RANKING order="3" place="3" resultid="10261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9560" />
                    <RANKING order="2" place="2" resultid="11732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12309" />
                    <RANKING order="2" place="2" resultid="10905" />
                    <RANKING order="3" place="3" resultid="10419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9511" />
                    <RANKING order="2" place="2" resultid="11295" />
                    <RANKING order="3" place="3" resultid="11312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11109" />
                    <RANKING order="2" place="2" resultid="11054" />
                    <RANKING order="3" place="3" resultid="9676" />
                    <RANKING order="4" place="4" resultid="11375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10413" />
                    <RANKING order="2" place="2" resultid="9965" />
                    <RANKING order="3" place="3" resultid="9855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10293" />
                    <RANKING order="2" place="-1" resultid="10727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1642" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1644" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1645" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1646" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14072" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14073" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14074" daytime="09:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14075" daytime="09:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1744" daytime="11:30" gender="M" number="38" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1745" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12398" />
                    <RANKING order="2" place="2" resultid="12174" />
                    <RANKING order="3" place="3" resultid="9432" />
                    <RANKING order="4" place="4" resultid="10452" />
                    <RANKING order="5" place="5" resultid="11697" />
                    <RANKING order="6" place="6" resultid="10882" />
                    <RANKING order="7" place="-1" resultid="10947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1746" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12413" />
                    <RANKING order="2" place="2" resultid="11564" />
                    <RANKING order="3" place="3" resultid="12186" />
                    <RANKING order="4" place="4" resultid="10480" />
                    <RANKING order="5" place="5" resultid="10113" />
                    <RANKING order="6" place="6" resultid="12462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1747" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11716" />
                    <RANKING order="2" place="2" resultid="10357" />
                    <RANKING order="3" place="3" resultid="10151" />
                    <RANKING order="4" place="4" resultid="10218" />
                    <RANKING order="5" place="5" resultid="9921" />
                    <RANKING order="6" place="-1" resultid="10036" />
                    <RANKING order="7" place="-1" resultid="11028" />
                    <RANKING order="8" place="-1" resultid="12348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1748" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11305" />
                    <RANKING order="2" place="2" resultid="10204" />
                    <RANKING order="3" place="3" resultid="10966" />
                    <RANKING order="4" place="4" resultid="10539" />
                    <RANKING order="5" place="5" resultid="9691" />
                    <RANKING order="6" place="-1" resultid="10043" />
                    <RANKING order="7" place="-1" resultid="11080" />
                    <RANKING order="8" place="-1" resultid="11725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1749" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12321" />
                    <RANKING order="2" place="2" resultid="11168" />
                    <RANKING order="3" place="3" resultid="11552" />
                    <RANKING order="4" place="4" resultid="9646" />
                    <RANKING order="5" place="5" resultid="11881" />
                    <RANKING order="6" place="6" resultid="10986" />
                    <RANKING order="7" place="7" resultid="10118" />
                    <RANKING order="8" place="8" resultid="9749" />
                    <RANKING order="9" place="9" resultid="11578" />
                    <RANKING order="10" place="-1" resultid="10319" />
                    <RANKING order="11" place="-1" resultid="10676" />
                    <RANKING order="12" place="-1" resultid="11581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1750" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9744" />
                    <RANKING order="2" place="2" resultid="11688" />
                    <RANKING order="3" place="3" resultid="10433" />
                    <RANKING order="4" place="4" resultid="10533" />
                    <RANKING order="5" place="5" resultid="12204" />
                    <RANKING order="6" place="6" resultid="9424" />
                    <RANKING order="7" place="7" resultid="10758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11344" />
                    <RANKING order="2" place="2" resultid="11283" />
                    <RANKING order="3" place="3" resultid="11969" />
                    <RANKING order="4" place="4" resultid="12330" />
                    <RANKING order="5" place="5" resultid="11433" />
                    <RANKING order="6" place="-1" resultid="12118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10193" />
                    <RANKING order="2" place="2" resultid="9644" />
                    <RANKING order="3" place="3" resultid="12460" />
                    <RANKING order="4" place="4" resultid="9624" />
                    <RANKING order="5" place="5" resultid="10241" />
                    <RANKING order="6" place="-1" resultid="9496" />
                    <RANKING order="7" place="-1" resultid="11558" />
                    <RANKING order="8" place="-1" resultid="11614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9727" />
                    <RANKING order="2" place="2" resultid="11117" />
                    <RANKING order="3" place="3" resultid="10021" />
                    <RANKING order="4" place="4" resultid="11960" />
                    <RANKING order="5" place="5" resultid="9652" />
                    <RANKING order="6" place="6" resultid="11545" />
                    <RANKING order="7" place="7" resultid="9479" />
                    <RANKING order="8" place="-1" resultid="9414" />
                    <RANKING order="9" place="-1" resultid="11814" />
                    <RANKING order="10" place="-1" resultid="12144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10256" />
                    <RANKING order="2" place="2" resultid="10818" />
                    <RANKING order="3" place="3" resultid="11414" />
                    <RANKING order="4" place="4" resultid="9353" />
                    <RANKING order="5" place="-1" resultid="12069" />
                    <RANKING order="6" place="-1" resultid="12136" />
                    <RANKING order="7" place="-1" resultid="12423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9420" />
                    <RANKING order="2" place="2" resultid="9405" />
                    <RANKING order="3" place="3" resultid="10189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9359" />
                    <RANKING order="2" place="2" resultid="11387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1758" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1760" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14106" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14107" daytime="11:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14108" daytime="11:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14109" daytime="12:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14110" daytime="12:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14111" daytime="12:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14112" daytime="12:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14113" daytime="12:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14114" daytime="12:35" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1681" daytime="10:25" gender="M" number="35" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1682" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12365" />
                    <RANKING order="2" place="2" resultid="10946" />
                    <RANKING order="3" place="3" resultid="11101" />
                    <RANKING order="4" place="4" resultid="11696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12485" />
                    <RANKING order="2" place="2" resultid="11476" />
                    <RANKING order="3" place="3" resultid="12412" />
                    <RANKING order="4" place="4" resultid="9540" />
                    <RANKING order="5" place="5" resultid="10495" />
                    <RANKING order="6" place="6" resultid="10789" />
                    <RANKING order="7" place="7" resultid="12335" />
                    <RANKING order="8" place="-1" resultid="10198" />
                    <RANKING order="9" place="-1" resultid="10929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12784" />
                    <RANKING order="2" place="2" resultid="10353" />
                    <RANKING order="3" place="3" resultid="10035" />
                    <RANKING order="4" place="4" resultid="12168" />
                    <RANKING order="5" place="5" resultid="10994" />
                    <RANKING order="6" place="6" resultid="10124" />
                    <RANKING order="7" place="7" resultid="12793" />
                    <RANKING order="8" place="8" resultid="10710" />
                    <RANKING order="9" place="-1" resultid="10217" />
                    <RANKING order="10" place="-1" resultid="12474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11995" />
                    <RANKING order="2" place="2" resultid="11336" />
                    <RANKING order="3" place="3" resultid="10958" />
                    <RANKING order="4" place="4" resultid="10283" />
                    <RANKING order="5" place="5" resultid="11079" />
                    <RANKING order="6" place="6" resultid="10965" />
                    <RANKING order="7" place="7" resultid="10979" />
                    <RANKING order="8" place="8" resultid="10974" />
                    <RANKING order="9" place="-1" resultid="10444" />
                    <RANKING order="10" place="-1" resultid="10746" />
                    <RANKING order="11" place="-1" resultid="10951" />
                    <RANKING order="12" place="-1" resultid="12374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11630" />
                    <RANKING order="2" place="2" resultid="11854" />
                    <RANKING order="3" place="3" resultid="11863" />
                    <RANKING order="4" place="4" resultid="11530" />
                    <RANKING order="5" place="5" resultid="11453" />
                    <RANKING order="6" place="6" resultid="10331" />
                    <RANKING order="7" place="7" resultid="10392" />
                    <RANKING order="8" place="8" resultid="11598" />
                    <RANKING order="9" place="9" resultid="10079" />
                    <RANKING order="10" place="10" resultid="12263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10901" />
                    <RANKING order="2" place="2" resultid="10432" />
                    <RANKING order="3" place="3" resultid="11060" />
                    <RANKING order="4" place="4" resultid="11903" />
                    <RANKING order="5" place="5" resultid="11898" />
                    <RANKING order="6" place="6" resultid="10075" />
                    <RANKING order="7" place="7" resultid="9762" />
                    <RANKING order="8" place="8" resultid="10532" />
                    <RANKING order="9" place="9" resultid="10757" />
                    <RANKING order="10" place="-1" resultid="11512" />
                    <RANKING order="11" place="-1" resultid="9743" />
                    <RANKING order="12" place="-1" resultid="11174" />
                    <RANKING order="13" place="-1" resultid="11873" />
                    <RANKING order="14" place="-1" resultid="12219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10233" />
                    <RANKING order="2" place="2" resultid="12159" />
                    <RANKING order="3" place="3" resultid="9719" />
                    <RANKING order="4" place="4" resultid="11405" />
                    <RANKING order="5" place="5" resultid="11327" />
                    <RANKING order="6" place="6" resultid="10399" />
                    <RANKING order="7" place="7" resultid="9684" />
                    <RANKING order="8" place="8" resultid="10268" />
                    <RANKING order="9" place="9" resultid="9903" />
                    <RANKING order="10" place="-1" resultid="9551" />
                    <RANKING order="11" place="-1" resultid="12117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11982" />
                    <RANKING order="2" place="2" resultid="12152" />
                    <RANKING order="3" place="3" resultid="9487" />
                    <RANKING order="4" place="4" resultid="11050" />
                    <RANKING order="5" place="5" resultid="11368" />
                    <RANKING order="6" place="-1" resultid="10738" />
                    <RANKING order="7" place="-1" resultid="12110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12196" />
                    <RANKING order="2" place="2" resultid="9948" />
                    <RANKING order="3" place="3" resultid="11032" />
                    <RANKING order="4" place="4" resultid="11575" />
                    <RANKING order="5" place="5" resultid="11821" />
                    <RANKING order="6" place="6" resultid="10054" />
                    <RANKING order="7" place="7" resultid="11544" />
                    <RANKING order="8" place="8" resultid="10813" />
                    <RANKING order="9" place="-1" resultid="9413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9483" />
                    <RANKING order="2" place="2" resultid="12422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9599" />
                    <RANKING order="2" place="2" resultid="12210" />
                    <RANKING order="3" place="3" resultid="10013" />
                    <RANKING order="4" place="4" resultid="9894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9980" />
                    <RANKING order="2" place="2" resultid="11386" />
                    <RANKING order="3" place="3" resultid="11977" />
                    <RANKING order="4" place="-1" resultid="9998" />
                    <RANKING order="5" place="-1" resultid="11022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10826" />
                    <RANKING order="2" place="-1" resultid="9957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10516" />
                    <RANKING order="2" place="2" resultid="12393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1697" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14088" daytime="10:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14089" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14090" daytime="10:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14091" daytime="10:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14092" daytime="10:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14093" daytime="10:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14094" daytime="10:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14095" daytime="10:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14096" daytime="10:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14097" daytime="10:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14098" daytime="10:45" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1664" daytime="10:20" gender="F" number="34" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1665" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9711" />
                    <RANKING order="2" place="2" resultid="10919" />
                    <RANKING order="3" place="3" resultid="10503" />
                    <RANKING order="4" place="4" resultid="10489" />
                    <RANKING order="5" place="5" resultid="10144" />
                    <RANKING order="6" place="6" resultid="10287" />
                    <RANKING order="7" place="7" resultid="9988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10096" />
                    <RANKING order="2" place="2" resultid="10131" />
                    <RANKING order="3" place="3" resultid="12771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12764" />
                    <RANKING order="2" place="2" resultid="12379" />
                    <RANKING order="3" place="3" resultid="10028" />
                    <RANKING order="4" place="4" resultid="10279" />
                    <RANKING order="5" place="5" resultid="11748" />
                    <RANKING order="6" place="6" resultid="10157" />
                    <RANKING order="7" place="-1" resultid="10314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11071" />
                    <RANKING order="2" place="2" resultid="12441" />
                    <RANKING order="3" place="3" resultid="11892" />
                    <RANKING order="4" place="4" resultid="9660" />
                    <RANKING order="5" place="-1" resultid="11739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10733" />
                    <RANKING order="2" place="2" resultid="11950" />
                    <RANKING order="3" place="3" resultid="12243" />
                    <RANKING order="4" place="4" resultid="10458" />
                    <RANKING order="5" place="5" resultid="10772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12236" />
                    <RANKING order="2" place="2" resultid="11589" />
                    <RANKING order="3" place="3" resultid="10778" />
                    <RANKING order="4" place="4" resultid="11942" />
                    <RANKING order="5" place="-1" resultid="9915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11398" />
                    <RANKING order="2" place="2" resultid="9517" />
                    <RANKING order="3" place="3" resultid="10246" />
                    <RANKING order="4" place="4" resultid="10910" />
                    <RANKING order="5" place="-1" resultid="11992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11289" />
                    <RANKING order="2" place="2" resultid="12251" />
                    <RANKING order="3" place="3" resultid="10766" />
                    <RANKING order="4" place="4" resultid="9668" />
                    <RANKING order="5" place="5" resultid="9677" />
                    <RANKING order="6" place="6" resultid="10473" />
                    <RANKING order="7" place="7" resultid="9972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12130" />
                    <RANKING order="2" place="2" resultid="9953" />
                    <RANKING order="3" place="3" resultid="12312" />
                    <RANKING order="4" place="4" resultid="11647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1676" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1677" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1678" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1679" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1680" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14083" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14084" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14085" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14086" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14087" daytime="10:25" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1721" daytime="11:00" gender="F" number="37" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1728" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11093" />
                    <RANKING order="2" place="2" resultid="10920" />
                    <RANKING order="3" place="3" resultid="9989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1729" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11681" />
                    <RANKING order="2" place="2" resultid="10888" />
                    <RANKING order="3" place="3" resultid="10097" />
                    <RANKING order="4" place="4" resultid="12258" />
                    <RANKING order="5" place="5" resultid="9838" />
                    <RANKING order="6" place="-1" resultid="12772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1730" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11662" />
                    <RANKING order="2" place="2" resultid="10525" />
                    <RANKING order="3" place="3" resultid="12779" />
                    <RANKING order="4" place="4" resultid="11672" />
                    <RANKING order="5" place="5" resultid="10309" />
                    <RANKING order="6" place="6" resultid="11749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1731" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10089" />
                    <RANKING order="2" place="2" resultid="11834" />
                    <RANKING order="3" place="3" resultid="12433" />
                    <RANKING order="4" place="-1" resultid="10465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1732" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10734" />
                    <RANKING order="2" place="2" resultid="11520" />
                    <RANKING order="3" place="3" resultid="10103" />
                    <RANKING order="4" place="4" resultid="11951" />
                    <RANKING order="5" place="-1" resultid="11825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1733" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11340" />
                    <RANKING order="2" place="2" resultid="11943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1734" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10247" />
                    <RANKING order="2" place="2" resultid="11296" />
                    <RANKING order="3" place="3" resultid="9847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1735" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11465" />
                    <RANKING order="2" place="2" resultid="11110" />
                    <RANKING order="3" place="3" resultid="10474" />
                    <RANKING order="4" place="-1" resultid="9973" />
                    <RANKING order="5" place="-1" resultid="12099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1737" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1740" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1741" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1742" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1743" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14102" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14103" daytime="11:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14104" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14105" daytime="11:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1698" daytime="10:45" gender="X" number="36" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1715" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10555" />
                    <RANKING order="2" place="2" resultid="10159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12822" />
                    <RANKING order="2" place="2" resultid="10365" />
                    <RANKING order="3" place="3" resultid="11907" />
                    <RANKING order="4" place="4" resultid="11541" />
                    <RANKING order="5" place="5" resultid="11751" />
                    <RANKING order="6" place="6" resultid="10830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1717" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9566" />
                    <RANKING order="2" place="2" resultid="11487" />
                    <RANKING order="3" place="3" resultid="11349" />
                    <RANKING order="4" place="4" resultid="12282" />
                    <RANKING order="5" place="5" resultid="11906" />
                    <RANKING order="6" place="6" resultid="11546" />
                    <RANKING order="7" place="7" resultid="12284" />
                    <RANKING order="8" place="8" resultid="10556" />
                    <RANKING order="9" place="-1" resultid="14186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1718" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9700" />
                    <RANKING order="2" place="2" resultid="11350" />
                    <RANKING order="3" place="3" resultid="11488" />
                    <RANKING order="4" place="4" resultid="10557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1719" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1720" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9981" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14099" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14100" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14101" daytime="10:55" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="12470" name="Aquasfera Masters Olsztyn">
          <CONTACT internet="annamariaaneczka@gmail.com" name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="12471">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="12472" heatid="13970" lane="9" entrytime="00:02:47.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="12473" heatid="14012" lane="8" entrytime="00:01:17.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="12474" heatid="14096" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11072" name="AquaStars Gdynia">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1978-11-20" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="11073">
              <RESULTS>
                <RESULT eventid="1113" points="335" reactiontime="+92" swimtime="00:02:44.04" resultid="11074" heatid="13925" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:02:05.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="367" reactiontime="+77" swimtime="00:00:33.56" resultid="11075" heatid="13951" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1239" points="275" reactiontime="+91" swimtime="00:03:15.25" resultid="11076" heatid="13967" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                    <SPLIT distance="150" swimtime="00:02:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="11077" heatid="14006" lane="8" entrytime="00:02:00.00" />
                <RESULT eventid="1440" points="461" reactiontime="+86" swimtime="00:00:29.02" resultid="11078" heatid="14022" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1681" points="424" reactiontime="+84" swimtime="00:00:35.16" resultid="11079" heatid="14089" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11080" heatid="14109" lane="5" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="12385" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1993-05-19" firstname="Łukasz" gender="M" lastname="Chmiel" nation="POL" license="100611700232" athleteid="12399">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="12400" heatid="13963" lane="5" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="12401" heatid="13977" lane="7" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="12402" heatid="14032" lane="3" />
                <RESULT eventid="1613" points="504" reactiontime="+75" swimtime="00:01:02.59" resultid="12403" heatid="14066" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="449" reactiontime="+41" swimtime="00:02:26.15" resultid="12404" heatid="14076" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:48.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-13" firstname="Tomasz" gender="M" lastname="Czermak" nation="POL" license="100611700216" athleteid="12405">
              <RESULTS>
                <RESULT eventid="1113" points="563" reactiontime="+79" swimtime="00:02:18.02" resultid="12406" heatid="13931" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                    <SPLIT distance="150" swimtime="00:01:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1165" points="519" reactiontime="+82" swimtime="00:18:03.80" resultid="12407" heatid="13943" lane="3" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                    <SPLIT distance="200" swimtime="00:02:16.10" />
                    <SPLIT distance="250" swimtime="00:02:51.74" />
                    <SPLIT distance="300" swimtime="00:03:27.68" />
                    <SPLIT distance="350" swimtime="00:04:03.90" />
                    <SPLIT distance="400" swimtime="00:04:40.28" />
                    <SPLIT distance="450" swimtime="00:05:16.26" />
                    <SPLIT distance="500" swimtime="00:05:52.45" />
                    <SPLIT distance="550" swimtime="00:06:28.90" />
                    <SPLIT distance="600" swimtime="00:07:05.58" />
                    <SPLIT distance="650" swimtime="00:07:42.10" />
                    <SPLIT distance="700" swimtime="00:08:18.70" />
                    <SPLIT distance="750" swimtime="00:08:55.19" />
                    <SPLIT distance="800" swimtime="00:09:31.81" />
                    <SPLIT distance="850" swimtime="00:10:08.51" />
                    <SPLIT distance="900" swimtime="00:10:45.13" />
                    <SPLIT distance="950" swimtime="00:11:21.80" />
                    <SPLIT distance="1000" swimtime="00:11:58.56" />
                    <SPLIT distance="1050" swimtime="00:12:35.64" />
                    <SPLIT distance="1100" swimtime="00:13:12.28" />
                    <SPLIT distance="1150" swimtime="00:13:48.77" />
                    <SPLIT distance="1200" swimtime="00:14:25.73" />
                    <SPLIT distance="1250" swimtime="00:15:02.47" />
                    <SPLIT distance="1300" swimtime="00:15:39.55" />
                    <SPLIT distance="1350" swimtime="00:16:16.08" />
                    <SPLIT distance="1400" swimtime="00:16:52.85" />
                    <SPLIT distance="1450" swimtime="00:17:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="545" reactiontime="+74" swimtime="00:02:35.48" resultid="12408" heatid="13970" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:54.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="432" reactiontime="+81" swimtime="00:02:27.40" resultid="12409" heatid="13995" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="572" reactiontime="+72" swimtime="00:01:09.76" resultid="12410" heatid="14013" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="486" reactiontime="+75" swimtime="00:02:09.66" resultid="12411" heatid="14053" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="551" reactiontime="+79" swimtime="00:00:32.21" resultid="12412" heatid="14098" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1744" points="505" swimtime="00:04:36.30" resultid="12413" heatid="14114" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                    <SPLIT distance="150" swimtime="00:01:39.14" />
                    <SPLIT distance="200" swimtime="00:02:14.39" />
                    <SPLIT distance="250" swimtime="00:02:50.10" />
                    <SPLIT distance="300" swimtime="00:03:26.30" />
                    <SPLIT distance="350" swimtime="00:04:02.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-29" firstname="Sławomir" gender="M" lastname="Smeja" nation="POL" license="100611700240" athleteid="12395">
              <RESULTS>
                <RESULT eventid="1165" points="654" reactiontime="+81" swimtime="00:16:43.38" resultid="12396" heatid="13943" lane="4" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.78" />
                    <SPLIT distance="150" swimtime="00:01:34.92" />
                    <SPLIT distance="200" swimtime="00:02:08.31" />
                    <SPLIT distance="250" swimtime="00:02:42.02" />
                    <SPLIT distance="300" swimtime="00:03:15.68" />
                    <SPLIT distance="350" swimtime="00:03:49.24" />
                    <SPLIT distance="400" swimtime="00:04:22.91" />
                    <SPLIT distance="450" swimtime="00:04:56.93" />
                    <SPLIT distance="500" swimtime="00:05:30.70" />
                    <SPLIT distance="550" swimtime="00:06:04.35" />
                    <SPLIT distance="600" swimtime="00:06:38.48" />
                    <SPLIT distance="650" swimtime="00:07:12.53" />
                    <SPLIT distance="700" swimtime="00:07:46.59" />
                    <SPLIT distance="750" swimtime="00:08:20.79" />
                    <SPLIT distance="800" swimtime="00:08:54.89" />
                    <SPLIT distance="850" swimtime="00:09:28.92" />
                    <SPLIT distance="900" swimtime="00:10:03.39" />
                    <SPLIT distance="950" swimtime="00:10:37.29" />
                    <SPLIT distance="1000" swimtime="00:11:11.24" />
                    <SPLIT distance="1050" swimtime="00:11:45.11" />
                    <SPLIT distance="1100" swimtime="00:12:18.91" />
                    <SPLIT distance="1150" swimtime="00:12:52.73" />
                    <SPLIT distance="1200" swimtime="00:13:26.52" />
                    <SPLIT distance="1250" swimtime="00:14:00.50" />
                    <SPLIT distance="1300" swimtime="00:14:34.07" />
                    <SPLIT distance="1350" swimtime="00:15:07.23" />
                    <SPLIT distance="1400" swimtime="00:15:40.47" />
                    <SPLIT distance="1450" swimtime="00:16:13.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="604" reactiontime="+81" swimtime="00:04:48.44" resultid="12397" heatid="14062" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="150" swimtime="00:01:42.46" />
                    <SPLIT distance="250" swimtime="00:03:01.97" />
                    <SPLIT distance="300" swimtime="00:03:43.87" />
                    <SPLIT distance="350" swimtime="00:04:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="641" reactiontime="+85" swimtime="00:04:15.19" resultid="12398" heatid="14114" lane="4" entrytime="00:04:07.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                    <SPLIT distance="100" swimtime="00:01:01.22" />
                    <SPLIT distance="150" swimtime="00:01:34.17" />
                    <SPLIT distance="200" swimtime="00:02:07.21" />
                    <SPLIT distance="250" swimtime="00:02:40.07" />
                    <SPLIT distance="300" swimtime="00:03:12.84" />
                    <SPLIT distance="350" swimtime="00:03:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="12386">
              <RESULTS>
                <RESULT eventid="1079" points="31" reactiontime="+107" swimtime="00:01:06.34" resultid="12387" heatid="13903" lane="3" />
                <RESULT comment="Rekord Polski" eventid="1165" points="27" reactiontime="+102" swimtime="00:47:50.02" resultid="12388" heatid="13939" lane="8" entrytime="00:47:39.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.62" />
                    <SPLIT distance="100" swimtime="00:02:49.12" />
                    <SPLIT distance="150" swimtime="00:04:25.30" />
                    <SPLIT distance="200" swimtime="00:05:58.29" />
                    <SPLIT distance="300" swimtime="00:09:05.30" />
                    <SPLIT distance="350" swimtime="00:10:39.51" />
                    <SPLIT distance="400" swimtime="00:12:13.59" />
                    <SPLIT distance="450" swimtime="00:13:51.32" />
                    <SPLIT distance="500" swimtime="00:15:23.95" />
                    <SPLIT distance="550" swimtime="00:17:04.16" />
                    <SPLIT distance="600" swimtime="00:18:37.18" />
                    <SPLIT distance="650" swimtime="00:20:13.42" />
                    <SPLIT distance="700" swimtime="00:21:48.60" />
                    <SPLIT distance="750" swimtime="00:23:28.01" />
                    <SPLIT distance="800" swimtime="00:25:04.56" />
                    <SPLIT distance="850" swimtime="00:26:42.33" />
                    <SPLIT distance="900" swimtime="00:28:20.14" />
                    <SPLIT distance="950" swimtime="00:30:00.45" />
                    <SPLIT distance="1000" swimtime="00:31:35.88" />
                    <SPLIT distance="1050" swimtime="00:33:15.98" />
                    <SPLIT distance="1100" swimtime="00:34:54.42" />
                    <SPLIT distance="1150" swimtime="00:39:54.69" />
                    <SPLIT distance="1200" swimtime="00:38:14.62" />
                    <SPLIT distance="1250" swimtime="00:43:14.08" />
                    <SPLIT distance="1300" swimtime="00:41:34.33" />
                    <SPLIT distance="1350" swimtime="00:46:25.50" />
                    <SPLIT distance="1400" swimtime="00:44:52.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="44" reactiontime="+98" swimtime="00:05:58.40" resultid="12389" heatid="13964" lane="8" entrytime="00:05:52.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.01" />
                    <SPLIT distance="100" swimtime="00:02:56.29" />
                    <SPLIT distance="150" swimtime="00:04:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="30" reactiontime="+80" swimtime="00:02:30.73" resultid="12390" heatid="13977" lane="3" entrytime="00:02:29.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="39" reactiontime="+56" swimtime="00:02:49.59" resultid="12391" heatid="14005" lane="3" entrytime="00:02:41.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="27" reactiontime="+130" swimtime="00:05:36.64" resultid="12392" heatid="14045" lane="7" entrytime="00:05:46.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.41" />
                    <SPLIT distance="100" swimtime="00:02:43.71" />
                    <SPLIT distance="150" swimtime="00:04:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="53" swimtime="00:01:10.23" resultid="12393" heatid="14089" lane="6" entrytime="00:01:08.08" />
                <RESULT eventid="1744" points="31" reactiontime="+101" swimtime="00:11:34.80" resultid="12394" heatid="14107" lane="8" entrytime="00:11:12.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.75" />
                    <SPLIT distance="100" swimtime="00:02:42.06" />
                    <SPLIT distance="150" swimtime="00:04:12.77" />
                    <SPLIT distance="200" swimtime="00:05:42.83" />
                    <SPLIT distance="250" swimtime="00:07:12.06" />
                    <SPLIT distance="300" swimtime="00:08:41.34" />
                    <SPLIT distance="350" swimtime="00:10:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CMUJKR" nation="POL" region="MAL" clubid="11169" name="Collegium Medicum UJ Masters Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="mariuszbaranik@gmail.com" name="Mariusz Baranik" phone="698128222" state="MAL" street="Białopradnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-08-22" firstname="Mirosław" gender="M" lastname="Woźniak" nation="POL" athleteid="11175">
              <RESULTS>
                <RESULT eventid="1113" points="339" reactiontime="+92" swimtime="00:02:43.43" resultid="11176" heatid="13928" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:02:06.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="389" reactiontime="+80" swimtime="00:01:04.24" resultid="11177" heatid="13984" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="305" reactiontime="+87" swimtime="00:01:26.04" resultid="11178" heatid="14009" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="355" reactiontime="+88" swimtime="00:00:31.65" resultid="11179" heatid="14024" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="11170">
              <RESULTS>
                <RESULT eventid="1079" points="426" reactiontime="+82" swimtime="00:00:27.77" resultid="11171" heatid="13914" lane="1" entrytime="00:00:27.20" />
                <RESULT eventid="1273" points="409" reactiontime="+86" swimtime="00:01:03.15" resultid="11172" heatid="13986" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="436" reactiontime="+77" swimtime="00:00:29.57" resultid="11173" heatid="14025" lane="5" entrytime="00:00:29.30" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="11174" heatid="14095" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LOD" clubid="10066" name="Delfin Masters Łódz">
          <CONTACT city="Łódz" email="cewa@poczta.fm" name="Cieplucha" phone="604627966" street="ul.Retkińska 74 m 18" zip="94-004" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-03" firstname="Piotr" gender="M" lastname="Gaede" nation="POL" athleteid="10076">
              <RESULTS>
                <RESULT eventid="1239" points="306" reactiontime="+87" swimtime="00:03:08.30" resultid="10077" heatid="13968" lane="0" entrytime="00:03:04.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="300" reactiontime="+83" swimtime="00:01:26.43" resultid="10078" heatid="14010" lane="0" entrytime="00:01:23.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="293" reactiontime="+81" swimtime="00:00:39.77" resultid="10079" heatid="14093" lane="4" entrytime="00:00:38.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="Cieplucha" nation="POL" athleteid="10080">
              <RESULTS>
                <RESULT eventid="1187" points="435" reactiontime="+66" swimtime="00:00:35.69" resultid="10081" heatid="13948" lane="0" entrytime="00:00:35.13" />
                <RESULT comment="Rekord Polski" eventid="1457" points="391" reactiontime="+64" swimtime="00:01:19.43" resultid="10082" heatid="14031" lane="1" entrytime="00:01:17.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="339" reactiontime="+70" swimtime="00:02:57.90" resultid="10083" heatid="14075" lane="1" entrytime="00:02:55.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:02:12.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-02-25" firstname="Jacek" gender="M" lastname="Kadłubiec" nation="POL" athleteid="10072">
              <RESULTS>
                <RESULT eventid="1239" points="318" reactiontime="+94" swimtime="00:03:06.06" resultid="10073" heatid="13969" lane="7" entrytime="00:02:51.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:26.09" />
                    <SPLIT distance="150" swimtime="00:02:14.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="318" reactiontime="+87" swimtime="00:01:24.82" resultid="10074" heatid="14010" lane="3" entrytime="00:01:20.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="325" swimtime="00:00:38.39" resultid="10075" heatid="14094" lane="6" entrytime="00:00:37.13" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="9415" name="Dynamo">
          <CONTACT city="Kharkiv" email="swimmer2003@ukr.net" name="Vadym Kutsenko" phone="038 057 7204282" street="Novgorodska" zip="61145" />
          <ATHLETES>
            <ATHLETE birthdate="1945-05-05" firstname="Vadym" gender="M" lastname="Kutsenko" nation="UKR" athleteid="9416">
              <RESULTS>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="9417" heatid="13941" lane="2" entrytime="00:22:40.49" entrycourse="LCM" />
                <RESULT eventid="1508" points="240" reactiontime="+110" swimtime="00:02:43.99" resultid="9418" heatid="14048" lane="7" entrytime="00:02:45.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:20.29" />
                    <SPLIT distance="150" swimtime="00:02:02.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="189" reactiontime="+127" swimtime="00:07:04.54" resultid="9419" heatid="14060" lane="6" entrytime="00:06:49.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:48.03" />
                    <SPLIT distance="150" swimtime="00:02:44.94" />
                    <SPLIT distance="200" swimtime="00:03:37.76" />
                    <SPLIT distance="250" swimtime="00:04:39.77" />
                    <SPLIT distance="300" swimtime="00:05:40.91" />
                    <SPLIT distance="350" swimtime="00:06:23.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="257" reactiontime="+128" swimtime="00:05:45.90" resultid="9420" heatid="14110" lane="6" entrytime="00:05:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:24.90" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                    <SPLIT distance="200" swimtime="00:02:53.49" />
                    <SPLIT distance="250" swimtime="00:03:37.60" />
                    <SPLIT distance="300" swimtime="00:04:21.08" />
                    <SPLIT distance="350" swimtime="00:05:04.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GBSPORT" nation="POL" region="PDK" clubid="10661" name="GB Sport Rzeszów">
          <CONTACT email="bartek@gbsport.pl" internet="www.gbsport.pl" name="Czarnota Bartłomiej" phone="603121020" state="PDK" />
          <ATHLETES>
            <ATHLETE birthdate="1977-02-01" firstname="Mariusz" gender="M" lastname="Wójcicki" nation="POL" athleteid="10677">
              <RESULTS>
                <RESULT eventid="1113" points="276" reactiontime="+86" swimtime="00:02:54.89" resultid="10678" heatid="13927" lane="0" entrytime="00:02:54.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:02:13.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="313" reactiontime="+67" swimtime="00:00:35.37" resultid="10679" heatid="13956" lane="7" entrytime="00:00:33.90" entrycourse="LCM" />
                <RESULT eventid="1341" points="250" reactiontime="+89" swimtime="00:02:56.81" resultid="10680" heatid="13992" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="252" reactiontime="+67" swimtime="00:01:22.13" resultid="10681" heatid="14036" lane="7" entrytime="00:01:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-05" firstname="Bartłomiej" gender="M" lastname="Czarnota" nation="POL" athleteid="10670">
              <RESULTS>
                <RESULT eventid="1079" points="495" reactiontime="+86" swimtime="00:00:26.42" resultid="10671" heatid="13912" lane="1" entrytime="00:00:28.90" entrycourse="LCM" />
                <RESULT eventid="1239" points="430" reactiontime="+90" swimtime="00:02:48.18" resultid="10672" heatid="13968" lane="6" entrytime="00:02:59.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:02:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="473" reactiontime="+85" swimtime="00:01:00.20" resultid="10673" heatid="13983" lane="3" entrytime="00:01:05.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="10674" heatid="14009" lane="9" entrytime="00:01:26.40" entrycourse="LCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="10675" heatid="14050" lane="7" entrytime="00:02:25.60" entrycourse="LCM" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="10676" heatid="14110" lane="7" entrytime="00:05:45.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-07-15" firstname="Grzegorz" gender="M" lastname="Wójcicki" nation="POL" athleteid="10682">
              <RESULTS>
                <RESULT eventid="1079" points="349" reactiontime="+75" swimtime="00:00:29.69" resultid="10683" heatid="13912" lane="8" entrytime="00:00:28.90" entrycourse="LCM" />
                <RESULT eventid="1205" points="241" reactiontime="+73" swimtime="00:00:38.58" resultid="10684" heatid="13954" lane="5" entrytime="00:00:36.20" entrycourse="LCM" />
                <RESULT eventid="1273" points="318" reactiontime="+74" swimtime="00:01:08.67" resultid="10685" heatid="13983" lane="2" entrytime="00:01:06.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="313" swimtime="00:00:33.01" resultid="10686" heatid="14022" lane="9" entrytime="00:00:33.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-17" firstname="Tomasz" gender="M" lastname="Pustelak" nation="POL" athleteid="10687">
              <RESULTS>
                <RESULT eventid="1079" points="374" reactiontime="+86" swimtime="00:00:29.02" resultid="10688" heatid="13913" lane="2" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="10689" heatid="13955" lane="1" entrytime="00:00:35.90" entrycourse="LCM" />
                <RESULT eventid="1273" points="361" swimtime="00:01:05.88" resultid="10690" heatid="13985" lane="9" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="10691" heatid="14023" lane="9" entrytime="00:00:32.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="10692" heatid="14056" lane="3" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10677" number="1" />
                    <RELAYPOSITION athleteid="10682" number="2" />
                    <RELAYPOSITION athleteid="10687" number="3" />
                    <RELAYPOSITION athleteid="10670" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="368" reactiontime="+69" swimtime="00:02:10.30" resultid="10693" heatid="13999" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:41.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10677" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="10670" number="2" />
                    <RELAYPOSITION athleteid="10682" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="10687" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9944" name="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Zuzanna" gender="F" lastname="Drążkiewicz" nation="POL" athleteid="9966">
              <RESULTS>
                <RESULT eventid="1062" points="48" reactiontime="+127" swimtime="00:01:05.13" resultid="9967" heatid="13896" lane="3" />
                <RESULT comment="(Time: 18:21), Przekroczony regulaminowy limit czasu." eventid="1147" reactiontime="+111" status="OTL" swimtime="00:00:00.00" resultid="9968" heatid="13935" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.63" />
                    <SPLIT distance="100" swimtime="00:02:33.97" />
                    <SPLIT distance="150" swimtime="00:03:59.87" />
                    <SPLIT distance="200" swimtime="00:05:25.48" />
                    <SPLIT distance="250" swimtime="00:06:53.43" />
                    <SPLIT distance="300" swimtime="00:08:22.40" />
                    <SPLIT distance="350" swimtime="00:09:49.17" />
                    <SPLIT distance="400" swimtime="00:11:16.89" />
                    <SPLIT distance="450" swimtime="00:12:43.11" />
                    <SPLIT distance="500" swimtime="00:14:08.95" />
                    <SPLIT distance="550" swimtime="00:15:34.10" />
                    <SPLIT distance="600" swimtime="00:17:01.91" />
                    <SPLIT distance="650" swimtime="00:18:28.87" />
                    <SPLIT distance="700" swimtime="00:19:52.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="58" reactiontime="+87" swimtime="00:01:09.79" resultid="9969" heatid="13944" lane="0" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="9970" heatid="13971" lane="9" />
                <RESULT eventid="1491" reactiontime="+108" status="DNF" swimtime="00:00:00.00" resultid="9971" heatid="14039" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="68" swimtime="00:01:12.07" resultid="9972" heatid="14083" lane="9" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="9973" heatid="14102" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="9949">
              <RESULTS>
                <RESULT eventid="1062" points="161" reactiontime="+102" swimtime="00:00:43.57" resultid="9950" heatid="13897" lane="8" entrytime="00:00:48.00" />
                <RESULT eventid="1187" points="114" reactiontime="+80" swimtime="00:00:55.67" resultid="9951" heatid="13945" lane="9" entrytime="00:00:56.00" />
                <RESULT eventid="1457" points="98" swimtime="00:02:05.68" resultid="9952" heatid="14028" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="123" swimtime="00:00:59.17" resultid="9953" heatid="14083" lane="6" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="9954">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="9955" heatid="13964" lane="4" entrytime="00:04:08.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="9956" heatid="14006" lane="2" entrytime="00:01:50.42" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="9957" heatid="14090" lane="3" entrytime="00:00:49.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="9945">
              <RESULTS>
                <RESULT eventid="1406" points="234" reactiontime="+98" swimtime="00:01:33.91" resultid="9946" heatid="14008" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="217" reactiontime="+124" swimtime="00:03:31.08" resultid="9947" heatid="13966" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:40.81" />
                    <SPLIT distance="150" swimtime="00:02:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="267" swimtime="00:00:41.00" resultid="9948" heatid="14092" lane="9" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="9974">
              <RESULTS>
                <RESULT eventid="1079" points="145" reactiontime="+110" swimtime="00:00:39.76" resultid="9975" heatid="13906" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1113" points="105" reactiontime="+119" swimtime="00:04:01.59" resultid="9976" heatid="13923" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.09" />
                    <SPLIT distance="100" swimtime="00:02:01.98" />
                    <SPLIT distance="150" swimtime="00:03:06.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="111" reactiontime="+101" swimtime="00:00:49.88" resultid="9977" heatid="13951" lane="5" entrytime="00:00:49.00" />
                <RESULT eventid="1273" points="112" reactiontime="+122" swimtime="00:01:37.21" resultid="9978" heatid="13979" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="128" swimtime="00:01:54.65" resultid="9979" heatid="14007" lane="9" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="178" reactiontime="+114" swimtime="00:00:46.93" resultid="9980" heatid="14091" lane="2" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="9958">
              <RESULTS>
                <RESULT eventid="1096" points="77" swimtime="00:04:55.55" resultid="9959" heatid="13919" lane="9" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.62" />
                    <SPLIT distance="100" swimtime="00:02:27.39" />
                    <SPLIT distance="150" swimtime="00:03:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="99" reactiontime="+71" swimtime="00:00:58.47" resultid="9960" heatid="13945" lane="8" entrytime="00:00:53.00" />
                <RESULT eventid="1324" points="44" reactiontime="+115" swimtime="00:05:42.50" resultid="9961" heatid="13990" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.02" />
                    <SPLIT distance="100" swimtime="00:02:43.53" />
                    <SPLIT distance="150" swimtime="00:04:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="43" reactiontime="+108" swimtime="00:01:09.34" resultid="9962" heatid="14014" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1457" points="92" reactiontime="+83" swimtime="00:02:08.59" resultid="9963" heatid="14029" lane="0" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="39" reactiontime="+107" swimtime="00:02:43.25" resultid="9964" heatid="14063" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="84" reactiontime="+78" swimtime="00:04:42.16" resultid="9965" heatid="14073" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:19.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="9981" heatid="14099" lane="4" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9958" number="1" />
                    <RELAYPOSITION athleteid="9954" number="2" />
                    <RELAYPOSITION athleteid="9974" number="3" />
                    <RELAYPOSITION athleteid="9949" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="9982" heatid="13933" lane="8" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9958" number="1" />
                    <RELAYPOSITION athleteid="9954" number="2" />
                    <RELAYPOSITION athleteid="9949" number="3" />
                    <RELAYPOSITION athleteid="9974" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10866" name="IKS Konstancin">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" license="103714700078" athleteid="10867">
              <RESULTS>
                <RESULT eventid="1079" points="430" swimtime="00:00:27.70" resultid="10868" heatid="13912" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="319" reactiontime="+79" swimtime="00:02:46.67" resultid="10869" heatid="13929" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:02:08.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="449" reactiontime="+73" swimtime="00:01:01.25" resultid="10870" heatid="13985" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="304" reactiontime="+83" swimtime="00:01:26.09" resultid="10871" heatid="14009" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="374" reactiontime="+79" swimtime="00:02:21.51" resultid="10872" heatid="14050" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:46.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="7000RUSE" nation="BUL" region="RUSE" clubid="10767" name="IRIS Ruse">
          <CONTACT city="Ruse" email="markomlight@abv.bg" name="Kamen Markov" phone="00359888806089" state="RUSE" street="Han Omurtaag 5" zip="7000" />
          <ATHLETES>
            <ATHLETE birthdate="1964-04-16" firstname="Kamen" gender="M" lastname="Markov" nation="BUL" license="BUL0346" athleteid="10796">
              <RESULTS>
                <RESULT eventid="1205" points="251" reactiontime="+82" swimtime="00:00:38.10" resultid="10797" heatid="13954" lane="6" entrytime="00:00:36.50" entrycourse="LCM" />
                <RESULT eventid="1273" points="260" reactiontime="+85" swimtime="00:01:13.43" resultid="10798" heatid="13982" lane="7" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="239" reactiontime="+75" swimtime="00:01:23.60" resultid="10799" heatid="14036" lane="9" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="173" reactiontime="+94" swimtime="00:03:03.03" resultid="10800" heatid="14048" lane="0" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="233" reactiontime="+84" swimtime="00:03:01.78" resultid="10801" heatid="14080" lane="1" entrytime="00:02:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:28.62" />
                    <SPLIT distance="150" swimtime="00:02:16.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-12-26" firstname="Krasimir" gender="M" lastname="Dinov" nation="BUL" license="BUL0350" athleteid="10810">
              <RESULTS>
                <RESULT eventid="1239" points="117" reactiontime="+106" swimtime="00:04:19.44" resultid="10811" heatid="13965" lane="0" entrytime="00:03:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.55" />
                    <SPLIT distance="100" swimtime="00:02:04.15" />
                    <SPLIT distance="150" swimtime="00:03:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="118" reactiontime="+96" swimtime="00:01:57.76" resultid="10812" heatid="14006" lane="5" entrytime="00:01:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="117" reactiontime="+98" swimtime="00:00:53.95" resultid="10813" heatid="14090" lane="1" entrytime="00:00:52.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-08-24" firstname="Nikola" gender="M" lastname="Gushterov" nation="BUL" license="BUL0359" athleteid="10784">
              <RESULTS>
                <RESULT eventid="1079" points="392" reactiontime="+82" swimtime="00:00:28.55" resultid="10785" heatid="13914" lane="6" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="350" reactiontime="+79" swimtime="00:01:06.56" resultid="10786" heatid="13985" lane="8" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="333" reactiontime="+78" swimtime="00:01:23.49" resultid="10787" heatid="14011" lane="5" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="362" reactiontime="+79" swimtime="00:00:31.47" resultid="10788" heatid="14024" lane="3" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1681" points="402" reactiontime="+79" swimtime="00:00:35.77" resultid="10789" heatid="14097" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-03-07" firstname="Konstantin" gender="M" lastname="Ivanov" nation="BUL" license="BUL0349" athleteid="10807">
              <RESULTS>
                <RESULT eventid="1341" points="79" reactiontime="+100" swimtime="00:04:19.66" resultid="10808" heatid="13993" lane="8" entrytime="00:03:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.47" />
                    <SPLIT distance="100" swimtime="00:02:03.30" />
                    <SPLIT distance="150" swimtime="00:03:12.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="123" reactiontime="+74" swimtime="00:03:44.90" resultid="10809" heatid="14078" lane="5" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.59" />
                    <SPLIT distance="100" swimtime="00:01:50.79" />
                    <SPLIT distance="150" swimtime="00:02:48.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Polina" gender="F" lastname="Davidova" nation="BUL" license="BUL0362" athleteid="10768">
              <RESULTS>
                <RESULT eventid="1062" points="197" reactiontime="+112" swimtime="00:00:40.78" resultid="10769" heatid="13898" lane="4" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="166" reactiontime="+56" swimtime="00:00:49.18" resultid="10770" heatid="13945" lane="4" entrytime="00:00:45.00" entrycourse="LCM" />
                <RESULT eventid="1423" points="117" reactiontime="+154" swimtime="00:00:49.91" resultid="10771" heatid="14015" lane="1" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1664" points="215" reactiontime="+96" swimtime="00:00:49.15" resultid="10772" heatid="14084" lane="4" entrytime="00:00:46.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-04-27" firstname="Nikolaj" gender="M" lastname="Handzhiev" nation="BUL" license="BUL0381" athleteid="10814">
              <RESULTS>
                <RESULT eventid="1113" points="122" reactiontime="+100" swimtime="00:03:49.26" resultid="10815" heatid="13923" lane="4" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:48.71" />
                    <SPLIT distance="150" swimtime="00:02:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="182" reactiontime="+105" swimtime="00:01:22.70" resultid="10816" heatid="13980" lane="0" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="167" reactiontime="+103" swimtime="00:03:05.14" resultid="10817" heatid="14046" lane="6" entrytime="00:03:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:26.78" />
                    <SPLIT distance="150" swimtime="00:02:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="155" reactiontime="+102" swimtime="00:06:49.30" resultid="10818" heatid="14108" lane="5" entrytime="00:06:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                    <SPLIT distance="200" swimtime="00:03:17.38" />
                    <SPLIT distance="250" swimtime="00:04:11.14" />
                    <SPLIT distance="300" swimtime="00:05:04.18" />
                    <SPLIT distance="350" swimtime="00:05:58.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-09-29" firstname="Evgenij" gender="M" lastname="Pejchev" nation="BUL" license="BUL0340" athleteid="10802">
              <RESULTS>
                <RESULT eventid="1079" points="217" reactiontime="+92" swimtime="00:00:34.78" resultid="10803" heatid="13907" lane="4" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="173" reactiontime="+94" swimtime="00:01:24.12" resultid="10804" heatid="13980" lane="8" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="151" swimtime="00:00:42.04" resultid="10805" heatid="14020" lane="9" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1613" reactiontime="+93" status="DNF" swimtime="00:00:00.00" resultid="10806" heatid="14067" lane="8" entrytime="00:01:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-07-25" firstname="Todor" gender="M" lastname="Todorov" nation="BUL" license="BUL0366" athleteid="10819">
              <RESULTS>
                <RESULT eventid="1079" points="69" reactiontime="+119" swimtime="00:00:50.88" resultid="10820" heatid="13904" lane="2" entrytime="00:00:47.00" entrycourse="LCM" />
                <RESULT eventid="1165" points="50" reactiontime="+119" swimtime="00:39:15.93" resultid="10821" heatid="13939" lane="1" entrytime="00:40:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.84" />
                    <SPLIT distance="100" swimtime="00:02:17.52" />
                    <SPLIT distance="150" swimtime="00:03:32.26" />
                    <SPLIT distance="200" swimtime="00:07:23.82" />
                    <SPLIT distance="250" swimtime="00:08:42.29" />
                    <SPLIT distance="300" swimtime="00:10:00.81" />
                    <SPLIT distance="350" swimtime="00:11:20.82" />
                    <SPLIT distance="400" swimtime="00:12:39.21" />
                    <SPLIT distance="450" swimtime="00:13:58.01" />
                    <SPLIT distance="500" swimtime="00:15:16.84" />
                    <SPLIT distance="550" swimtime="00:16:35.71" />
                    <SPLIT distance="600" swimtime="00:17:54.11" />
                    <SPLIT distance="650" swimtime="00:19:14.06" />
                    <SPLIT distance="700" swimtime="00:20:32.43" />
                    <SPLIT distance="750" swimtime="00:21:53.89" />
                    <SPLIT distance="800" swimtime="00:23:14.16" />
                    <SPLIT distance="850" swimtime="00:24:34.49" />
                    <SPLIT distance="900" swimtime="00:25:54.17" />
                    <SPLIT distance="950" swimtime="00:27:13.27" />
                    <SPLIT distance="1000" swimtime="00:28:30.02" />
                    <SPLIT distance="1050" swimtime="00:29:51.73" />
                    <SPLIT distance="1100" swimtime="00:31:11.55" />
                    <SPLIT distance="1150" swimtime="00:32:32.20" />
                    <SPLIT distance="1200" swimtime="00:33:53.36" />
                    <SPLIT distance="1450" swimtime="00:37:59.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="53" reactiontime="+92" swimtime="00:01:03.80" resultid="10822" heatid="13949" lane="5" entrytime="00:02:00.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="56" reactiontime="+106" swimtime="00:02:01.97" resultid="10823" heatid="13978" lane="8" entrytime="00:01:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="24" reactiontime="+119" swimtime="00:01:17.12" resultid="10824" heatid="14019" lane="0" entrytime="00:01:08.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="43" reactiontime="+67" swimtime="00:02:27.85" resultid="10825" heatid="14032" lane="5" entrytime="00:04:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K10 - Dłonie przeniesione poza linię bioder (z wyjątkiem pierwszego ruchu ramon po starcie i nawrotach (Time: 10:59), K-8, K-9" eventid="1681" reactiontime="+100" status="DSQ" swimtime="00:01:18.83" resultid="10826" heatid="14089" lane="8" entrytime="00:01:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-08" firstname="Veselina" gender="F" lastname="Borisova" nation="BUL" license="BUL0331" athleteid="10773">
              <RESULTS>
                <RESULT eventid="1062" points="233" reactiontime="+108" swimtime="00:00:38.54" resultid="10774" heatid="13899" lane="0" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1222" points="137" reactiontime="+101" swimtime="00:04:29.81" resultid="10775" heatid="13960" lane="3" entrytime="00:03:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.75" />
                    <SPLIT distance="100" swimtime="00:01:59.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="182" swimtime="00:01:31.79" resultid="10776" heatid="13973" lane="9" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="107" reactiontime="+104" swimtime="00:00:51.36" resultid="10777" heatid="14015" lane="8" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1664" points="194" reactiontime="+104" swimtime="00:00:50.91" resultid="10778" heatid="14084" lane="2" entrytime="00:00:48.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-05" firstname="Ivelin" gender="M" lastname="Ivanov" nation="BUL" license="BUL0344" athleteid="10790">
              <RESULTS>
                <RESULT eventid="1239" points="211" reactiontime="+100" swimtime="00:03:33.30" resultid="10791" heatid="13966" lane="5" entrytime="00:03:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:42.51" />
                    <SPLIT distance="150" swimtime="00:02:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="250" reactiontime="+103" swimtime="00:01:14.44" resultid="10792" heatid="13982" lane="4" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="227" reactiontime="+87" swimtime="00:01:34.81" resultid="10793" heatid="14008" lane="3" entrytime="00:01:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="195" swimtime="00:01:29.51" resultid="10794" heatid="14035" lane="4" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="201" swimtime="00:03:10.87" resultid="10795" heatid="14080" lane="8" entrytime="00:02:56.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-17" firstname="Jankov" gender="M" lastname="Javor" nation="BUL" license="BUL368" athleteid="10779">
              <RESULTS>
                <RESULT eventid="1079" points="341" reactiontime="+92" swimtime="00:00:29.91" resultid="10780" heatid="13914" lane="4" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1205" points="352" reactiontime="+75" swimtime="00:00:34.04" resultid="10781" heatid="13957" lane="3" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="314" reactiontime="+73" swimtime="00:01:16.38" resultid="10782" heatid="14038" lane="0" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="298" reactiontime="+76" swimtime="00:02:47.48" resultid="10783" heatid="14082" lane="7" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:02:02.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="165" reactiontime="+76" swimtime="00:02:34.59" resultid="10827" heatid="14055" lane="7" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                    <SPLIT distance="150" swimtime="00:01:59.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10790" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="10814" number="2" />
                    <RELAYPOSITION athleteid="10819" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="10796" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="148" reactiontime="+79" swimtime="00:02:56.59" resultid="10828" heatid="13997" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10796" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="10790" number="2" />
                    <RELAYPOSITION athleteid="10802" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="10819" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="238" reactiontime="+82" swimtime="00:02:16.86" resultid="10829" heatid="13933" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="150" swimtime="00:01:39.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10779" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="10768" number="2" />
                    <RELAYPOSITION athleteid="10773" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="10784" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="232" reactiontime="+65" swimtime="00:02:31.97" resultid="10830" heatid="14100" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10779" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="10768" number="2" />
                    <RELAYPOSITION athleteid="10784" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="10773" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="11805" name="K.S.niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="11806">
              <RESULTS>
                <RESULT eventid="1113" points="164" reactiontime="+123" swimtime="00:03:28.20" resultid="11807" heatid="13922" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                    <SPLIT distance="100" swimtime="00:01:40.57" />
                    <SPLIT distance="150" swimtime="00:02:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="177" swimtime="00:25:49.96" resultid="11808" heatid="13941" lane="9" entrytime="00:24:58.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:34.25" />
                    <SPLIT distance="150" swimtime="00:02:25.39" />
                    <SPLIT distance="200" swimtime="00:03:17.21" />
                    <SPLIT distance="250" swimtime="00:04:09.90" />
                    <SPLIT distance="300" swimtime="00:05:01.83" />
                    <SPLIT distance="350" swimtime="00:05:54.24" />
                    <SPLIT distance="400" swimtime="00:06:47.26" />
                    <SPLIT distance="450" swimtime="00:07:39.82" />
                    <SPLIT distance="500" swimtime="00:08:32.40" />
                    <SPLIT distance="550" swimtime="00:09:25.26" />
                    <SPLIT distance="600" swimtime="00:10:18.16" />
                    <SPLIT distance="650" swimtime="00:11:10.82" />
                    <SPLIT distance="700" swimtime="00:12:03.58" />
                    <SPLIT distance="750" swimtime="00:12:56.08" />
                    <SPLIT distance="800" swimtime="00:13:49.00" />
                    <SPLIT distance="850" swimtime="00:14:42.19" />
                    <SPLIT distance="900" swimtime="00:15:34.68" />
                    <SPLIT distance="950" swimtime="00:16:26.77" />
                    <SPLIT distance="1000" swimtime="00:17:19.53" />
                    <SPLIT distance="1050" swimtime="00:18:11.57" />
                    <SPLIT distance="1100" swimtime="00:19:03.80" />
                    <SPLIT distance="1150" swimtime="00:19:55.62" />
                    <SPLIT distance="1200" swimtime="00:20:47.86" />
                    <SPLIT distance="1250" swimtime="00:21:39.72" />
                    <SPLIT distance="1300" swimtime="00:22:31.05" />
                    <SPLIT distance="1350" swimtime="00:23:22.66" />
                    <SPLIT distance="1400" swimtime="00:24:13.75" />
                    <SPLIT distance="1450" swimtime="00:25:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="181" reactiontime="+70" swimtime="00:01:31.66" resultid="11809" heatid="14034" lane="6" entrytime="00:01:31.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="185" reactiontime="+67" swimtime="00:03:16.15" resultid="11810" heatid="14079" lane="7" entrytime="00:03:15.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:35.47" />
                    <SPLIT distance="150" swimtime="00:02:26.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-04" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="11815">
              <RESULTS>
                <RESULT eventid="1113" points="146" reactiontime="+98" swimtime="00:03:36.25" resultid="11816" heatid="13924" lane="0" entrytime="00:03:35.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="173" reactiontime="+82" swimtime="00:03:47.59" resultid="11817" heatid="13965" lane="2" entrytime="00:03:47.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:49.72" />
                    <SPLIT distance="150" swimtime="00:02:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="186" reactiontime="+89" swimtime="00:01:41.34" resultid="11818" heatid="14007" lane="2" entrytime="00:01:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="176" reactiontime="+107" swimtime="00:00:40.00" resultid="11819" heatid="14019" lane="3" entrytime="00:00:40.35" />
                <RESULT eventid="1613" points="116" reactiontime="+87" swimtime="00:01:41.97" resultid="11820" heatid="14067" lane="7" entrytime="00:01:39.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="203" reactiontime="+82" swimtime="00:00:44.91" resultid="11821" heatid="14091" lane="3" entrytime="00:00:43.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="11811">
              <RESULTS>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="11813" heatid="14059" lane="3" entrytime="00:08:20.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11814" heatid="14108" lane="9" entrytime="00:06:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="11822">
              <RESULTS>
                <RESULT eventid="1096" points="120" reactiontime="+107" swimtime="00:04:15.34" resultid="11823" heatid="13919" lane="7" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.52" />
                    <SPLIT distance="100" swimtime="00:02:09.96" />
                    <SPLIT distance="150" swimtime="00:03:16.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="11824" heatid="14039" lane="3" entrytime="00:03:35.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="11825" heatid="14102" lane="3" entrytime="00:07:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KR" nation="POL" region="KR" clubid="11351" name="Korona Kraków Masters">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="11431">
              <RESULTS>
                <RESULT eventid="1165" points="201" swimtime="00:24:45.29" resultid="11432" heatid="13940" lane="6" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:28.25" />
                    <SPLIT distance="150" swimtime="00:02:15.87" />
                    <SPLIT distance="200" swimtime="00:03:04.23" />
                    <SPLIT distance="250" swimtime="00:03:53.15" />
                    <SPLIT distance="300" swimtime="00:04:42.13" />
                    <SPLIT distance="350" swimtime="00:05:32.26" />
                    <SPLIT distance="400" swimtime="00:06:21.61" />
                    <SPLIT distance="450" swimtime="00:07:11.79" />
                    <SPLIT distance="500" swimtime="00:08:02.06" />
                    <SPLIT distance="550" swimtime="00:08:52.88" />
                    <SPLIT distance="600" swimtime="00:09:43.17" />
                    <SPLIT distance="650" swimtime="00:10:33.70" />
                    <SPLIT distance="700" swimtime="00:11:24.27" />
                    <SPLIT distance="750" swimtime="00:12:15.11" />
                    <SPLIT distance="800" swimtime="00:13:05.11" />
                    <SPLIT distance="850" swimtime="00:13:55.58" />
                    <SPLIT distance="900" swimtime="00:14:45.62" />
                    <SPLIT distance="950" swimtime="00:15:36.12" />
                    <SPLIT distance="1000" swimtime="00:16:26.64" />
                    <SPLIT distance="1050" swimtime="00:17:17.16" />
                    <SPLIT distance="1100" swimtime="00:18:07.06" />
                    <SPLIT distance="1150" swimtime="00:18:57.33" />
                    <SPLIT distance="1200" swimtime="00:19:47.46" />
                    <SPLIT distance="1250" swimtime="00:20:38.68" />
                    <SPLIT distance="1300" swimtime="00:21:29.26" />
                    <SPLIT distance="1350" swimtime="00:22:19.96" />
                    <SPLIT distance="1400" swimtime="00:23:09.92" />
                    <SPLIT distance="1450" swimtime="00:23:59.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="215" reactiontime="+92" swimtime="00:06:06.80" resultid="11433" heatid="14109" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:24.40" />
                    <SPLIT distance="150" swimtime="00:02:10.80" />
                    <SPLIT distance="200" swimtime="00:02:58.58" />
                    <SPLIT distance="250" swimtime="00:03:46.21" />
                    <SPLIT distance="300" swimtime="00:04:34.34" />
                    <SPLIT distance="350" swimtime="00:05:21.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="11441">
              <RESULTS>
                <RESULT eventid="1079" points="83" reactiontime="+100" swimtime="00:00:47.82" resultid="11442" heatid="13904" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1113" points="32" swimtime="00:05:57.78" resultid="11443" heatid="13923" lane="9" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.16" />
                    <SPLIT distance="100" swimtime="00:02:51.84" />
                    <SPLIT distance="150" swimtime="00:04:54.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="43" reactiontime="+82" swimtime="00:01:08.12" resultid="11444" heatid="13949" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1273" points="69" reactiontime="+123" swimtime="00:01:54.22" resultid="11445" heatid="13978" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="19" swimtime="00:01:22.67" resultid="11446" heatid="14019" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="1508" points="52" swimtime="00:04:31.68" resultid="11447" heatid="14045" lane="6" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.97" />
                    <SPLIT distance="100" swimtime="00:02:05.73" />
                    <SPLIT distance="150" swimtime="00:03:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11448" heatid="14077" lane="0" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz- Musiał" nation="POL" athleteid="11369">
              <RESULTS>
                <RESULT eventid="1062" points="137" reactiontime="+99" swimtime="00:00:45.98" resultid="11370" heatid="13897" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1147" points="121" reactiontime="+102" swimtime="00:16:24.57" resultid="11371" heatid="13935" lane="5" entrytime="00:15:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:51.21" />
                    <SPLIT distance="150" swimtime="00:02:52.05" />
                    <SPLIT distance="200" swimtime="00:03:54.18" />
                    <SPLIT distance="250" swimtime="00:04:56.41" />
                    <SPLIT distance="300" swimtime="00:06:04.50" />
                    <SPLIT distance="350" swimtime="00:07:07.96" />
                    <SPLIT distance="400" swimtime="00:08:11.08" />
                    <SPLIT distance="450" swimtime="00:09:14.52" />
                    <SPLIT distance="500" swimtime="00:10:15.99" />
                    <SPLIT distance="550" swimtime="00:11:18.74" />
                    <SPLIT distance="600" swimtime="00:12:21.75" />
                    <SPLIT distance="650" swimtime="00:13:24.12" />
                    <SPLIT distance="700" swimtime="00:14:25.32" />
                    <SPLIT distance="750" swimtime="00:15:26.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="74" reactiontime="+116" swimtime="00:04:49.79" resultid="11372" heatid="13990" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.87" />
                    <SPLIT distance="100" swimtime="00:02:17.35" />
                    <SPLIT distance="150" swimtime="00:03:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="93" reactiontime="+114" swimtime="00:09:51.21" resultid="11373" heatid="14057" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.62" />
                    <SPLIT distance="100" swimtime="00:02:22.58" />
                    <SPLIT distance="150" swimtime="00:03:42.08" />
                    <SPLIT distance="200" swimtime="00:05:00.36" />
                    <SPLIT distance="250" swimtime="00:06:25.53" />
                    <SPLIT distance="300" swimtime="00:07:49.12" />
                    <SPLIT distance="350" swimtime="00:08:52.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="72" reactiontime="+113" swimtime="00:02:13.19" resultid="11374" heatid="14063" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="83" reactiontime="+46" swimtime="00:04:44.34" resultid="11375" heatid="14073" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.56" />
                    <SPLIT distance="100" swimtime="00:02:15.92" />
                    <SPLIT distance="150" swimtime="00:03:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="11392">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="503" reactiontime="+76" swimtime="00:00:29.83" resultid="11393" heatid="13902" lane="0" entrytime="00:00:29.80" />
                <RESULT comment="Rekord Polski" eventid="1187" points="431" reactiontime="+60" swimtime="00:00:35.80" resultid="11394" heatid="13947" lane="5" entrytime="00:00:36.00" />
                <RESULT comment="Rekord Polski" eventid="1256" points="437" reactiontime="+71" swimtime="00:01:08.61" resultid="11395" heatid="13976" lane="8" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1388" points="420" reactiontime="+74" swimtime="00:01:25.89" resultid="11396" heatid="14001" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="423" reactiontime="+73" swimtime="00:00:32.53" resultid="11397" heatid="14017" lane="2" entrytime="00:00:32.50" />
                <RESULT comment="Rekord Polski" eventid="1664" points="506" reactiontime="+70" swimtime="00:00:36.99" resultid="11398" heatid="14087" lane="3" entrytime="00:00:36.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-04" firstname="Dawid" gender="M" lastname="Deszcz" nation="POL" athleteid="11471">
              <RESULTS>
                <RESULT eventid="1079" points="157" reactiontime="+98" swimtime="00:00:38.69" resultid="11472" heatid="13904" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Piotr" gender="M" lastname="Frankiewicz" nation="POL" athleteid="11473">
              <RESULTS>
                <RESULT eventid="1239" points="472" reactiontime="+76" swimtime="00:02:43.08" resultid="11474" heatid="13970" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:57.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="541" reactiontime="+75" swimtime="00:01:11.08" resultid="11475" heatid="14013" lane="4" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="556" reactiontime="+74" swimtime="00:00:32.12" resultid="11476" heatid="14098" lane="7" entrytime="00:00:31.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="11457">
              <RESULTS>
                <RESULT eventid="1062" points="342" reactiontime="+94" swimtime="00:00:33.92" resultid="11458" heatid="13900" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1147" points="277" reactiontime="+95" swimtime="00:12:27.35" resultid="11459" heatid="13937" lane="0" entrytime="00:12:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:23.04" />
                    <SPLIT distance="150" swimtime="00:02:09.63" />
                    <SPLIT distance="200" swimtime="00:02:57.13" />
                    <SPLIT distance="250" swimtime="00:03:45.11" />
                    <SPLIT distance="300" swimtime="00:04:32.59" />
                    <SPLIT distance="350" swimtime="00:05:20.86" />
                    <SPLIT distance="400" swimtime="00:06:08.71" />
                    <SPLIT distance="450" swimtime="00:06:56.96" />
                    <SPLIT distance="500" swimtime="00:07:44.96" />
                    <SPLIT distance="550" swimtime="00:08:33.17" />
                    <SPLIT distance="600" swimtime="00:09:20.86" />
                    <SPLIT distance="650" swimtime="00:10:08.56" />
                    <SPLIT distance="700" swimtime="00:10:56.10" />
                    <SPLIT distance="750" swimtime="00:11:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="312" reactiontime="+96" swimtime="00:01:16.71" resultid="11460" heatid="13974" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="11461" heatid="13991" lane="1" entrytime="00:03:20.00" />
                <RESULT eventid="1423" points="249" swimtime="00:00:38.80" resultid="11462" heatid="14016" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1491" points="279" reactiontime="+101" swimtime="00:02:52.85" resultid="11463" heatid="14042" lane="7" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1595" points="236" reactiontime="+103" swimtime="00:01:29.97" resultid="11464" heatid="14064" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="283" swimtime="00:06:02.92" resultid="11465" heatid="14104" lane="6" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:11.35" />
                    <SPLIT distance="200" swimtime="00:02:58.32" />
                    <SPLIT distance="250" swimtime="00:03:45.41" />
                    <SPLIT distance="300" swimtime="00:04:31.90" />
                    <SPLIT distance="350" swimtime="00:05:19.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="11434">
              <RESULTS>
                <RESULT eventid="1205" points="119" reactiontime="+101" swimtime="00:00:48.85" resultid="11435" heatid="13951" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1273" points="108" reactiontime="+86" swimtime="00:01:38.50" resultid="11436" heatid="13978" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="91" reactiontime="+78" swimtime="00:04:08.73" resultid="11437" heatid="14078" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.91" />
                    <SPLIT distance="100" swimtime="00:02:00.99" />
                    <SPLIT distance="150" swimtime="00:03:06.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="11466">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="11467" heatid="13899" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1222" points="344" reactiontime="+90" swimtime="00:03:18.45" resultid="11468" heatid="13961" lane="5" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:35.42" />
                    <SPLIT distance="150" swimtime="00:02:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="332" reactiontime="+95" swimtime="00:01:32.86" resultid="11469" heatid="14003" lane="0" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="204" reactiontime="+85" swimtime="00:01:38.57" resultid="11470" heatid="14029" lane="4" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="11376">
              <RESULTS>
                <RESULT eventid="1079" points="82" reactiontime="+152" swimtime="00:00:47.99" resultid="11377" heatid="13904" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1205" points="71" reactiontime="+99" swimtime="00:00:57.90" resultid="11378" heatid="13950" lane="9" entrytime="00:01:02.00" />
                <RESULT eventid="1474" points="72" reactiontime="+104" swimtime="00:02:04.76" resultid="11379" heatid="14033" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="72" reactiontime="+100" swimtime="00:04:28.55" resultid="11380" heatid="14078" lane="9" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.98" />
                    <SPLIT distance="100" swimtime="00:02:10.14" />
                    <SPLIT distance="150" swimtime="00:03:19.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="11399">
              <RESULTS>
                <RESULT eventid="1079" points="331" reactiontime="+92" swimtime="00:00:30.20" resultid="11400" heatid="13909" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1205" points="281" reactiontime="+81" swimtime="00:00:36.69" resultid="11401" heatid="13955" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1440" points="348" swimtime="00:00:31.88" resultid="11402" heatid="14024" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="264" reactiontime="+73" swimtime="00:01:20.96" resultid="11403" heatid="14035" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="274" reactiontime="+103" swimtime="00:01:16.67" resultid="11404" heatid="14069" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="317" reactiontime="+97" swimtime="00:00:38.72" resultid="11405" heatid="14093" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="11449">
              <RESULTS>
                <RESULT eventid="1239" points="338" reactiontime="+92" swimtime="00:03:02.33" resultid="11450" heatid="13964" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:15.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="336" reactiontime="+77" swimtime="00:01:23.27" resultid="11451" heatid="14010" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11452" heatid="14076" lane="4" />
                <RESULT eventid="1681" points="341" reactiontime="+78" swimtime="00:00:37.81" resultid="11453" heatid="14095" lane="7" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="11438">
              <RESULTS>
                <RESULT eventid="1062" points="280" reactiontime="+107" swimtime="00:00:36.27" resultid="11439" heatid="13899" lane="8" entrytime="00:00:36.50" />
                <RESULT eventid="1096" points="187" reactiontime="+110" swimtime="00:03:40.47" resultid="11440" heatid="13919" lane="6" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.32" />
                    <SPLIT distance="100" swimtime="00:01:46.69" />
                    <SPLIT distance="150" swimtime="00:02:50.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="11381">
              <RESULTS>
                <RESULT eventid="1079" points="93" swimtime="00:00:46.09" resultid="11382" heatid="13905" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1165" points="89" reactiontime="+120" swimtime="00:32:27.58" resultid="11383" heatid="13939" lane="2" entrytime="00:32:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                    <SPLIT distance="100" swimtime="00:02:05.62" />
                    <SPLIT distance="150" swimtime="00:03:13.96" />
                    <SPLIT distance="200" swimtime="00:04:20.98" />
                    <SPLIT distance="250" swimtime="00:05:27.93" />
                    <SPLIT distance="300" swimtime="00:06:34.70" />
                    <SPLIT distance="350" swimtime="00:07:42.38" />
                    <SPLIT distance="400" swimtime="00:08:47.23" />
                    <SPLIT distance="450" swimtime="00:09:52.96" />
                    <SPLIT distance="500" swimtime="00:10:58.62" />
                    <SPLIT distance="550" swimtime="00:12:05.50" />
                    <SPLIT distance="600" swimtime="00:13:11.43" />
                    <SPLIT distance="650" swimtime="00:14:16.82" />
                    <SPLIT distance="700" swimtime="00:15:20.73" />
                    <SPLIT distance="750" swimtime="00:16:25.84" />
                    <SPLIT distance="800" swimtime="00:17:30.76" />
                    <SPLIT distance="850" swimtime="00:18:35.43" />
                    <SPLIT distance="900" swimtime="00:19:40.53" />
                    <SPLIT distance="950" swimtime="00:20:44.11" />
                    <SPLIT distance="1000" swimtime="00:21:48.24" />
                    <SPLIT distance="1050" swimtime="00:22:52.34" />
                    <SPLIT distance="1100" swimtime="00:23:58.32" />
                    <SPLIT distance="1150" swimtime="00:25:03.14" />
                    <SPLIT distance="1200" swimtime="00:26:07.59" />
                    <SPLIT distance="1250" swimtime="00:27:13.84" />
                    <SPLIT distance="1300" swimtime="00:28:17.28" />
                    <SPLIT distance="1350" swimtime="00:29:22.73" />
                    <SPLIT distance="1400" swimtime="00:30:26.36" />
                    <SPLIT distance="1450" swimtime="00:31:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="93" reactiontime="+105" swimtime="00:01:43.42" resultid="11384" heatid="13978" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="71" reactiontime="+101" swimtime="00:04:05.91" resultid="11385" heatid="14045" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.33" />
                    <SPLIT distance="100" swimtime="00:01:56.24" />
                    <SPLIT distance="150" swimtime="00:03:02.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="77" reactiontime="+105" swimtime="00:01:02.02" resultid="11386" heatid="14089" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1744" points="77" swimtime="00:08:36.93" resultid="11387" heatid="14107" lane="6" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.42" />
                    <SPLIT distance="100" swimtime="00:02:03.72" />
                    <SPLIT distance="150" swimtime="00:03:13.51" />
                    <SPLIT distance="200" swimtime="00:04:19.21" />
                    <SPLIT distance="250" swimtime="00:05:28.22" />
                    <SPLIT distance="300" swimtime="00:06:32.69" />
                    <SPLIT distance="350" swimtime="00:07:39.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="11428">
              <RESULTS>
                <RESULT eventid="1079" points="504" reactiontime="+74" swimtime="00:00:26.26" resultid="11429" heatid="13916" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="492" reactiontime="+72" swimtime="00:00:59.41" resultid="11430" heatid="13986" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-03" firstname="Marcin" gender="M" lastname="Wyżga" nation="POL" athleteid="11424">
              <RESULTS>
                <RESULT eventid="1273" points="360" reactiontime="+83" swimtime="00:01:05.93" resultid="11425" heatid="13983" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="362" reactiontime="+81" swimtime="00:00:31.47" resultid="11426" heatid="14024" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11427" heatid="14076" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="11477">
              <RESULTS>
                <RESULT eventid="1062" points="234" reactiontime="+98" swimtime="00:00:38.48" resultid="11478" heatid="13898" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1096" points="159" reactiontime="+110" swimtime="00:03:52.38" resultid="11479" heatid="13918" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:53.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="11415">
              <RESULTS>
                <RESULT eventid="1062" points="52" swimtime="00:01:03.24" resultid="11416" heatid="13897" lane="9" entrytime="00:00:59.00" />
                <RESULT eventid="1096" points="42" reactiontime="+111" swimtime="00:06:02.19" resultid="11417" heatid="13918" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.69" />
                    <SPLIT distance="100" swimtime="00:03:05.51" />
                    <SPLIT distance="150" swimtime="00:04:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="65" reactiontime="+115" swimtime="00:05:45.75" resultid="11418" heatid="13959" lane="3" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.73" />
                    <SPLIT distance="100" swimtime="00:02:44.49" />
                    <SPLIT distance="150" swimtime="00:04:20.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="53" reactiontime="+112" swimtime="00:02:17.86" resultid="11419" heatid="13971" lane="8" entrytime="00:02:10.00" />
                <RESULT eventid="1423" points="28" reactiontime="+125" swimtime="00:01:20.00" resultid="11420" heatid="14014" lane="3" entrytime="00:01:15.00" />
                <RESULT comment="Rekord Polski" eventid="1555" points="42" reactiontime="+118" swimtime="00:12:50.42" resultid="11421" heatid="14057" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.32" />
                    <SPLIT distance="100" swimtime="00:03:10.74" />
                    <SPLIT distance="150" swimtime="00:04:59.88" />
                    <SPLIT distance="200" swimtime="00:06:53.20" />
                    <SPLIT distance="250" swimtime="00:08:31.35" />
                    <SPLIT distance="300" swimtime="00:12:47.52" />
                    <SPLIT distance="350" swimtime="00:11:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="26" reactiontime="+114" swimtime="00:03:07.67" resultid="11422" heatid="14063" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="54" reactiontime="+109" swimtime="00:10:27.85" resultid="11423" heatid="14102" lane="7" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.16" />
                    <SPLIT distance="100" swimtime="00:02:28.37" />
                    <SPLIT distance="200" swimtime="00:05:15.90" />
                    <SPLIT distance="250" swimtime="00:06:35.37" />
                    <SPLIT distance="300" swimtime="00:07:57.29" />
                    <SPLIT distance="350" swimtime="00:09:16.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-10-20" firstname="Janusz" gender="M" lastname="Toporski" nation="POL" athleteid="11360">
              <RESULTS>
                <RESULT eventid="1079" points="166" reactiontime="+86" swimtime="00:00:37.99" resultid="11361" heatid="13905" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1113" points="120" swimtime="00:03:50.87" resultid="11362" heatid="13924" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.16" />
                    <SPLIT distance="100" swimtime="00:02:03.08" />
                    <SPLIT distance="150" swimtime="00:03:02.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="148" reactiontime="+112" swimtime="00:04:00.08" resultid="11363" heatid="13965" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.38" />
                    <SPLIT distance="100" swimtime="00:01:59.57" />
                    <SPLIT distance="150" swimtime="00:03:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="94" swimtime="00:04:04.91" resultid="11364" heatid="13993" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                    <SPLIT distance="100" swimtime="00:01:58.42" />
                    <SPLIT distance="150" swimtime="00:03:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="131" reactiontime="+93" swimtime="00:01:53.88" resultid="11365" heatid="14006" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="126" reactiontime="+107" swimtime="00:08:05.75" resultid="11366" heatid="14059" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:56.24" />
                    <SPLIT distance="150" swimtime="00:03:04.44" />
                    <SPLIT distance="200" swimtime="00:04:10.57" />
                    <SPLIT distance="250" swimtime="00:05:12.59" />
                    <SPLIT distance="300" swimtime="00:06:15.19" />
                    <SPLIT distance="350" swimtime="00:07:11.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="87" reactiontime="+95" swimtime="00:01:52.23" resultid="11367" heatid="14066" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="133" reactiontime="+88" swimtime="00:00:51.64" resultid="11368" heatid="14090" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="11406">
              <RESULTS>
                <RESULT eventid="1079" points="202" reactiontime="+128" swimtime="00:00:35.58" resultid="11407" heatid="13908" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1113" points="128" reactiontime="+131" swimtime="00:03:45.92" resultid="11408" heatid="13924" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.31" />
                    <SPLIT distance="100" swimtime="00:01:53.21" />
                    <SPLIT distance="150" swimtime="00:03:01.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="217" reactiontime="+131" swimtime="00:01:18.00" resultid="11409" heatid="13981" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="58" reactiontime="+134" swimtime="00:04:47.47" resultid="11410" heatid="13992" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.81" />
                    <SPLIT distance="100" swimtime="00:02:12.33" />
                    <SPLIT distance="150" swimtime="00:03:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="162" reactiontime="+128" swimtime="00:03:06.92" resultid="11411" heatid="14047" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="150" swimtime="00:02:19.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="96" reactiontime="+139" swimtime="00:08:51.27" resultid="11412" heatid="14059" lane="5" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.81" />
                    <SPLIT distance="100" swimtime="00:02:06.33" />
                    <SPLIT distance="150" swimtime="00:03:16.89" />
                    <SPLIT distance="200" swimtime="00:04:30.56" />
                    <SPLIT distance="250" swimtime="00:05:41.47" />
                    <SPLIT distance="300" swimtime="00:06:54.19" />
                    <SPLIT distance="350" swimtime="00:07:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="80" swimtime="00:01:55.30" resultid="11413" heatid="14067" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="140" reactiontime="+134" swimtime="00:07:03.35" resultid="11414" heatid="14108" lane="4" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:40.74" />
                    <SPLIT distance="200" swimtime="00:03:26.53" />
                    <SPLIT distance="300" swimtime="00:05:15.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="11388">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="513" reactiontime="+79" swimtime="00:00:29.64" resultid="11389" heatid="13902" lane="8" entrytime="00:00:29.60" />
                <RESULT eventid="1256" points="488" reactiontime="+76" swimtime="00:01:06.10" resultid="11390" heatid="13976" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1423" points="408" reactiontime="+74" swimtime="00:00:32.93" resultid="11391" heatid="14017" lane="8" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="11454">
              <RESULTS>
                <RESULT eventid="1165" points="379" reactiontime="+92" swimtime="00:20:02.85" resultid="11455" heatid="13942" lane="7" entrytime="00:21:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:55.93" />
                    <SPLIT distance="200" swimtime="00:02:36.27" />
                    <SPLIT distance="250" swimtime="00:03:16.51" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                    <SPLIT distance="350" swimtime="00:04:36.66" />
                    <SPLIT distance="400" swimtime="00:05:16.52" />
                    <SPLIT distance="450" swimtime="00:05:56.45" />
                    <SPLIT distance="500" swimtime="00:06:36.21" />
                    <SPLIT distance="550" swimtime="00:07:15.99" />
                    <SPLIT distance="600" swimtime="00:07:55.63" />
                    <SPLIT distance="650" swimtime="00:08:35.46" />
                    <SPLIT distance="700" swimtime="00:09:15.19" />
                    <SPLIT distance="750" swimtime="00:09:54.90" />
                    <SPLIT distance="800" swimtime="00:10:35.19" />
                    <SPLIT distance="850" swimtime="00:11:15.15" />
                    <SPLIT distance="900" swimtime="00:11:55.56" />
                    <SPLIT distance="950" swimtime="00:12:35.32" />
                    <SPLIT distance="1000" swimtime="00:13:16.39" />
                    <SPLIT distance="1050" swimtime="00:13:57.46" />
                    <SPLIT distance="1100" swimtime="00:14:37.59" />
                    <SPLIT distance="1150" swimtime="00:15:17.94" />
                    <SPLIT distance="1200" swimtime="00:15:58.02" />
                    <SPLIT distance="1250" swimtime="00:16:41.98" />
                    <SPLIT distance="1300" swimtime="00:17:21.42" />
                    <SPLIT distance="1350" swimtime="00:18:05.29" />
                    <SPLIT distance="1400" swimtime="00:18:44.94" />
                    <SPLIT distance="1450" swimtime="00:19:24.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="377" reactiontime="+88" swimtime="00:02:34.23" resultid="11456" heatid="13995" lane="2" entrytime="00:02:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="337" reactiontime="+68" swimtime="00:02:14.19" resultid="11482" heatid="13999" lane="2" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11454" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="11449" number="2" />
                    <RELAYPOSITION athleteid="11424" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="11428" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Korona Kraków F" number="5">
              <RESULTS>
                <RESULT eventid="1381" points="83" reactiontime="+94" swimtime="00:03:33.59" resultid="11483" heatid="13997" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.33" />
                    <SPLIT distance="100" swimtime="00:02:03.88" />
                    <SPLIT distance="150" swimtime="00:02:45.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11376" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="11381" number="2" />
                    <RELAYPOSITION athleteid="11406" number="3" />
                    <RELAYPOSITION athleteid="11441" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="9">
              <RESULTS>
                <RESULT eventid="1548" points="231" reactiontime="+90" swimtime="00:02:18.15" resultid="11485" heatid="14055" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="150" swimtime="00:01:33.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11399" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="11406" number="2" />
                    <RELAYPOSITION athleteid="11449" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="11381" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1358" points="377" reactiontime="+60" swimtime="00:02:27.02" resultid="11481" heatid="13996" lane="6" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:01:52.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11392" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="11466" number="2" />
                    <RELAYPOSITION athleteid="11388" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="11457" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="6">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1525" points="394" reactiontime="+79" swimtime="00:02:11.74" resultid="11484" heatid="14054" lane="6" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11388" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="11466" number="2" />
                    <RELAYPOSITION athleteid="11457" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="11392" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków C" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1130" points="391" reactiontime="+72" swimtime="00:01:55.95" resultid="11480" heatid="13934" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:00.20" />
                    <SPLIT distance="150" swimtime="00:01:29.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11392" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="11454" number="2" />
                    <RELAYPOSITION athleteid="11388" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="11428" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D" number="2">
              <RESULTS>
                <RESULT eventid="1698" points="160" reactiontime="+50" swimtime="00:02:51.83" resultid="11488" heatid="14100" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.33" />
                    <SPLIT distance="100" swimtime="00:01:38.17" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11369" number="1" reactiontime="+50" />
                    <RELAYPOSITION athleteid="11399" number="2" />
                    <RELAYPOSITION athleteid="11457" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="11406" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków E" number="7">
              <RESULTS>
                <RESULT eventid="1130" points="205" reactiontime="+113" swimtime="00:02:23.72" resultid="11486" heatid="13933" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:46.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11438" number="1" reactiontime="+113" />
                    <RELAYPOSITION athleteid="11457" number="2" />
                    <RELAYPOSITION athleteid="11406" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="11360" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków C" number="8">
              <RESULTS>
                <RESULT eventid="1698" points="365" reactiontime="+67" swimtime="00:02:10.63" resultid="11487" heatid="14101" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:07.94" />
                    <SPLIT distance="150" swimtime="00:01:41.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11449" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="11473" number="2" />
                    <RELAYPOSITION athleteid="11392" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="11388" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="PŁYWAK" nation="POL" region="WAR" clubid="10911" name="KPiRS PŁYWAK">
          <CONTACT city="Płock" email="pawel.powichrowski@wp.pl" name="Powichrowski Paweł" phone="603694397" state="MAZ" street="Wiatraki 11 B" zip="09-402" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-30" firstname="Łukasz" gender="M" lastname="Szypryt" nation="POL" athleteid="10921">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="10922" heatid="13903" lane="4" />
                <RESULT eventid="1113" points="283" reactiontime="+85" swimtime="00:02:53.60" resultid="10923" heatid="13927" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="367" reactiontime="+64" swimtime="00:00:33.55" resultid="10924" heatid="13956" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1239" points="322" reactiontime="+86" swimtime="00:03:05.28" resultid="10925" heatid="13968" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                    <SPLIT distance="100" swimtime="00:01:32.05" />
                    <SPLIT distance="150" swimtime="00:02:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="326" reactiontime="+86" swimtime="00:01:24.14" resultid="10926" heatid="14011" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="313" reactiontime="+69" swimtime="00:01:16.43" resultid="10927" heatid="14036" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="235" reactiontime="+76" swimtime="00:03:01.15" resultid="10928" heatid="14080" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:31.12" />
                    <SPLIT distance="150" swimtime="00:02:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10929" heatid="14096" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-04-28" firstname="Karolina" gender="F" lastname="Kowalska" nation="POL" athleteid="10930">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="10931" heatid="13918" lane="1" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="10932" heatid="13937" lane="6" entrytime="00:10:58.63" />
                <RESULT eventid="1187" points="292" reactiontime="+109" swimtime="00:00:40.75" resultid="10933" heatid="13947" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1222" points="288" reactiontime="+97" swimtime="00:03:30.63" resultid="10934" heatid="13962" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                    <SPLIT distance="100" swimtime="00:01:40.42" />
                    <SPLIT distance="150" swimtime="00:02:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="300" reactiontime="+95" swimtime="00:00:36.48" resultid="10935" heatid="14016" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="1457" points="297" reactiontime="+108" swimtime="00:01:27.05" resultid="10936" heatid="14030" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="208" reactiontime="+96" swimtime="00:01:33.89" resultid="10937" heatid="14064" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="271" reactiontime="+101" swimtime="00:03:11.62" resultid="10938" heatid="14074" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.79" />
                    <SPLIT distance="100" swimtime="00:01:34.60" />
                    <SPLIT distance="150" swimtime="00:02:24.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-07-04" firstname="Agata" gender="F" lastname="Olejniczak" nation="POL" athleteid="10912">
              <RESULTS>
                <RESULT eventid="1062" points="519" reactiontime="+88" swimtime="00:00:29.52" resultid="10913" heatid="13902" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1096" points="317" reactiontime="+90" swimtime="00:03:04.93" resultid="10914" heatid="13920" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:19.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="363" reactiontime="+86" swimtime="00:00:37.92" resultid="10915" heatid="13947" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1222" points="336" reactiontime="+92" swimtime="00:03:19.95" resultid="10916" heatid="13962" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:36.17" />
                    <SPLIT distance="150" swimtime="00:02:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="387" reactiontime="+90" swimtime="00:01:28.29" resultid="10917" heatid="14003" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="365" reactiontime="+93" swimtime="00:02:38.05" resultid="10918" heatid="14043" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="407" reactiontime="+98" swimtime="00:00:39.77" resultid="10919" heatid="14087" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1721" points="260" reactiontime="+97" swimtime="00:06:13.40" resultid="10920" heatid="14105" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:22.74" />
                    <SPLIT distance="150" swimtime="00:02:09.09" />
                    <SPLIT distance="200" swimtime="00:02:57.37" />
                    <SPLIT distance="250" swimtime="00:03:46.15" />
                    <SPLIT distance="300" swimtime="00:04:35.09" />
                    <SPLIT distance="350" swimtime="00:05:24.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-23" firstname="Paweł" gender="M" lastname="Powichrowski" nation="POL" athleteid="10948">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="10949" heatid="13908" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="10950" heatid="13949" lane="2" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10951" heatid="14092" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-09" firstname="Piotr" gender="M" lastname="Mikuła" nation="POL" athleteid="10939">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="10940" heatid="13917" lane="7" entrytime="00:00:25.12" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="10941" heatid="13928" lane="7" entrytime="00:02:45.00" />
                <RESULT eventid="1205" points="389" reactiontime="+104" swimtime="00:00:32.91" resultid="10942" heatid="13949" lane="3" />
                <RESULT eventid="1273" points="571" reactiontime="+77" swimtime="00:00:56.54" resultid="10943" heatid="13989" lane="2" entrytime="00:00:56.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="415" reactiontime="+75" swimtime="00:01:17.62" resultid="10944" heatid="14010" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="388" reactiontime="+79" swimtime="00:02:19.83" resultid="10945" heatid="14044" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:03.75" />
                    <SPLIT distance="150" swimtime="00:01:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="526" reactiontime="+75" swimtime="00:00:32.71" resultid="10946" heatid="14097" lane="3" entrytime="00:00:33.39" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="10947" heatid="14113" lane="1" entrytime="00:04:55.83" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04211" nation="POL" region="11" clubid="11642" name="KS Delfin Gliwice">
          <CONTACT email="ksdelfin@op,pl" name="Cupiał Jarosław" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="11643">
              <RESULTS>
                <RESULT eventid="1187" points="44" reactiontime="+88" swimtime="00:01:16.53" resultid="11644" heatid="13944" lane="9" />
                <RESULT eventid="1222" points="102" reactiontime="+105" swimtime="00:04:57.63" resultid="11645" heatid="13959" lane="4" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.12" />
                    <SPLIT distance="100" swimtime="00:02:24.57" />
                    <SPLIT distance="150" swimtime="00:03:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="100" reactiontime="+119" swimtime="00:02:18.45" resultid="11646" heatid="14000" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="102" reactiontime="+103" swimtime="00:01:03.08" resultid="11647" heatid="14083" lane="1" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="9348" name="KS Extreme Team Oborniki">
          <CONTACT city="Oborniki" email="janwol@poczta.onet.pl" name="Wolniewicz Janusz" phone="791064667" street="Czarnkowska 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="9349">
              <RESULTS>
                <RESULT comment="(Time: 19:41), Przekroczony regulaminowy limit czasu." eventid="1165" reactiontime="+98" status="OTL" swimtime="00:31:10.63" resultid="9350" heatid="13939" lane="5" entrytime="00:29:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:43.43" />
                    <SPLIT distance="150" swimtime="00:02:42.67" />
                    <SPLIT distance="200" swimtime="00:03:42.91" />
                    <SPLIT distance="250" swimtime="00:04:42.99" />
                    <SPLIT distance="300" swimtime="00:05:43.55" />
                    <SPLIT distance="350" swimtime="00:06:45.34" />
                    <SPLIT distance="400" swimtime="00:07:46.38" />
                    <SPLIT distance="450" swimtime="00:08:47.91" />
                    <SPLIT distance="500" swimtime="00:09:48.85" />
                    <SPLIT distance="550" swimtime="00:10:51.47" />
                    <SPLIT distance="600" swimtime="00:11:54.01" />
                    <SPLIT distance="650" swimtime="00:12:57.48" />
                    <SPLIT distance="700" swimtime="00:14:00.15" />
                    <SPLIT distance="750" swimtime="00:15:04.36" />
                    <SPLIT distance="800" swimtime="00:16:08.10" />
                    <SPLIT distance="850" swimtime="00:17:11.52" />
                    <SPLIT distance="900" swimtime="00:18:14.83" />
                    <SPLIT distance="950" swimtime="00:19:18.65" />
                    <SPLIT distance="1000" swimtime="00:20:22.86" />
                    <SPLIT distance="1050" swimtime="00:21:27.90" />
                    <SPLIT distance="1100" swimtime="00:22:32.16" />
                    <SPLIT distance="1150" swimtime="00:23:36.84" />
                    <SPLIT distance="1200" swimtime="00:24:40.97" />
                    <SPLIT distance="1250" swimtime="00:25:49.05" />
                    <SPLIT distance="1300" swimtime="00:26:54.64" />
                    <SPLIT distance="1350" swimtime="00:28:00.60" />
                    <SPLIT distance="1400" swimtime="00:29:06.28" />
                    <SPLIT distance="1450" swimtime="00:30:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="162" reactiontime="+105" swimtime="00:01:26.03" resultid="9351" heatid="13979" lane="5" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="105" reactiontime="+94" swimtime="00:03:36.15" resultid="9352" heatid="14046" lane="8" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:43.96" />
                    <SPLIT distance="150" swimtime="00:02:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="118" reactiontime="+102" swimtime="00:07:28.45" resultid="9353" heatid="14107" lane="5" entrytime="00:07:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:41.62" />
                    <SPLIT distance="150" swimtime="00:02:38.94" />
                    <SPLIT distance="200" swimtime="00:03:37.43" />
                    <SPLIT distance="250" swimtime="00:04:36.65" />
                    <SPLIT distance="300" swimtime="00:05:35.04" />
                    <SPLIT distance="350" swimtime="00:06:34.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="9904" name="KS Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="9905">
              <RESULTS>
                <RESULT eventid="1113" points="302" swimtime="00:02:49.91" resultid="9906" heatid="13927" lane="9" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="327" reactiontime="+85" swimtime="00:00:34.86" resultid="9907" heatid="13949" lane="0" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="9908" heatid="13968" lane="1" entrytime="00:03:00.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="312" swimtime="00:01:16.58" resultid="9909" heatid="14036" lane="6" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="299" reactiontime="+79" swimtime="00:02:47.29" resultid="9910" heatid="14080" lane="4" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="12708" name="KS REKIN Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="12794">
              <RESULTS>
                <RESULT eventid="1079" points="536" reactiontime="+75" swimtime="00:00:25.73" resultid="12795" heatid="13915" lane="2" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1113" points="522" reactiontime="+76" swimtime="00:02:21.55" resultid="12796" heatid="13931" lane="7" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="100" swimtime="00:01:05.40" />
                    <SPLIT distance="150" swimtime="00:01:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="595" reactiontime="+59" swimtime="00:00:28.58" resultid="12797" heatid="13958" lane="3" entrytime="00:00:28.87" />
                <RESULT comment="Rekord Polski" eventid="1341" points="466" reactiontime="+80" swimtime="00:02:23.73" resultid="12798" heatid="13992" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                    <SPLIT distance="100" swimtime="00:01:02.78" />
                    <SPLIT distance="150" swimtime="00:01:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="572" reactiontime="+74" swimtime="00:00:27.02" resultid="12799" heatid="14018" lane="3" />
                <RESULT eventid="1474" points="557" reactiontime="+62" swimtime="00:01:03.10" resultid="12800" heatid="14038" lane="5" entrytime="00:01:02.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="534" reactiontime="+84" swimtime="00:01:01.37" resultid="12801" heatid="14066" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="481" reactiontime="+63" swimtime="00:02:22.76" resultid="12802" heatid="14082" lane="3" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="150" swimtime="00:01:45.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="12765">
              <RESULTS>
                <RESULT eventid="1062" points="367" reactiontime="+93" swimtime="00:00:33.13" resultid="12766" heatid="13901" lane="8" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="223" reactiontime="+105" swimtime="00:03:49.22" resultid="12767" heatid="13960" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                    <SPLIT distance="100" swimtime="00:01:49.36" />
                    <SPLIT distance="150" swimtime="00:02:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="313" swimtime="00:01:16.65" resultid="12768" heatid="13975" lane="9" entrytime="00:01:14.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="218" reactiontime="+101" swimtime="00:01:46.81" resultid="12769" heatid="14001" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="264" reactiontime="+105" swimtime="00:02:55.91" resultid="12770" heatid="14041" lane="0" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="243" reactiontime="+97" swimtime="00:00:47.21" resultid="12771" heatid="14084" lane="7" entrytime="00:00:49.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="12772" heatid="14104" lane="0" entrytime="00:06:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="StuczyńSki" nation="POL" athleteid="12780">
              <RESULTS>
                <RESULT eventid="1079" points="540" reactiontime="+78" swimtime="00:00:25.67" resultid="12781" heatid="13916" lane="7" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="513" reactiontime="+81" swimtime="00:00:58.59" resultid="12782" heatid="13989" lane="6" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="504" reactiontime="+80" swimtime="00:01:12.78" resultid="12783" heatid="14013" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="576" swimtime="00:00:31.75" resultid="12784" heatid="14098" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="12773">
              <RESULTS>
                <RESULT eventid="1147" points="260" reactiontime="+78" swimtime="00:12:42.94" resultid="12774" heatid="13936" lane="5" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:25.61" />
                    <SPLIT distance="150" swimtime="00:02:12.99" />
                    <SPLIT distance="200" swimtime="00:03:01.28" />
                    <SPLIT distance="250" swimtime="00:03:51.13" />
                    <SPLIT distance="300" swimtime="00:04:40.26" />
                    <SPLIT distance="350" swimtime="00:05:28.85" />
                    <SPLIT distance="400" swimtime="00:06:17.23" />
                    <SPLIT distance="450" swimtime="00:07:06.10" />
                    <SPLIT distance="500" swimtime="00:07:54.63" />
                    <SPLIT distance="550" swimtime="00:08:43.43" />
                    <SPLIT distance="600" swimtime="00:09:32.21" />
                    <SPLIT distance="650" swimtime="00:10:21.25" />
                    <SPLIT distance="700" swimtime="00:11:09.64" />
                    <SPLIT distance="750" swimtime="00:11:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="259" reactiontime="+84" swimtime="00:03:37.98" resultid="12775" heatid="13961" lane="0" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="100" swimtime="00:01:45.55" />
                    <SPLIT distance="150" swimtime="00:02:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="234" reactiontime="+79" swimtime="00:01:44.39" resultid="12776" heatid="14001" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="279" reactiontime="+78" swimtime="00:02:52.78" resultid="12777" heatid="14041" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="150" swimtime="00:02:08.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="251" reactiontime="+81" swimtime="00:03:16.61" resultid="12778" heatid="14074" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:36.15" />
                    <SPLIT distance="150" swimtime="00:02:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="276" reactiontime="+81" swimtime="00:06:06.02" resultid="12779" heatid="14103" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:25.91" />
                    <SPLIT distance="150" swimtime="00:02:12.43" />
                    <SPLIT distance="200" swimtime="00:02:59.99" />
                    <SPLIT distance="250" swimtime="00:03:47.22" />
                    <SPLIT distance="300" swimtime="00:04:34.89" />
                    <SPLIT distance="350" swimtime="00:05:21.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="12785">
              <RESULTS>
                <RESULT eventid="1079" points="514" reactiontime="+76" swimtime="00:00:26.09" resultid="12786" heatid="13915" lane="4" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1113" points="320" swimtime="00:02:46.65" resultid="12787" heatid="13931" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:16.48" />
                    <SPLIT distance="150" swimtime="00:02:05.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="449" reactiontime="+65" swimtime="00:00:31.39" resultid="12788" heatid="13958" lane="2" entrytime="00:00:29.90" />
                <RESULT eventid="1273" points="494" reactiontime="+78" swimtime="00:00:59.33" resultid="12789" heatid="13988" lane="8" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="506" reactiontime="+76" swimtime="00:00:28.13" resultid="12790" heatid="14026" lane="4" entrytime="00:00:27.90" />
                <RESULT eventid="1508" points="416" reactiontime="+74" swimtime="00:02:16.53" resultid="12791" heatid="14044" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="416" swimtime="00:01:06.70" resultid="12792" heatid="14071" lane="9" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="374" reactiontime="+82" swimtime="00:00:36.65" resultid="12793" heatid="14096" lane="1" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="12758">
              <RESULTS>
                <RESULT eventid="1062" points="547" reactiontime="+81" swimtime="00:00:29.01" resultid="12759" heatid="13902" lane="1" entrytime="00:00:29.47" entrycourse="SCM" />
                <RESULT eventid="1222" points="457" reactiontime="+80" swimtime="00:03:00.54" resultid="12760" heatid="13959" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="525" reactiontime="+78" swimtime="00:01:04.52" resultid="12761" heatid="13976" lane="6" entrytime="00:01:04.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="494" reactiontime="+76" swimtime="00:01:21.36" resultid="12762" heatid="14004" lane="5" entrytime="00:01:19.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="464" reactiontime="+80" swimtime="00:02:25.93" resultid="12763" heatid="14039" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="490" reactiontime="+76" swimtime="00:00:37.38" resultid="12764" heatid="14087" lane="5" entrytime="00:00:36.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Rekin Świebodzice B" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="390" reactiontime="+76" swimtime="00:01:56.10" resultid="12821" heatid="13932" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.79" />
                    <SPLIT distance="100" swimtime="00:00:54.18" />
                    <SPLIT distance="150" swimtime="00:01:29.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12780" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="12785" number="2" />
                    <RELAYPOSITION athleteid="12758" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="12773" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="382" reactiontime="+92" swimtime="00:02:08.68" resultid="12822" heatid="14099" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:40.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12765" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="12780" number="2" />
                    <RELAYPOSITION athleteid="12794" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="12758" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="10558" name="Ks Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502499565" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="11317">
              <RESULTS>
                <RESULT eventid="1079" points="439" reactiontime="+76" swimtime="00:00:27.50" resultid="11318" heatid="13913" lane="5" entrytime="00:00:27.90" />
                <RESULT eventid="1205" points="440" reactiontime="+67" swimtime="00:00:31.60" resultid="11319" heatid="13958" lane="9" entrytime="00:00:30.90" />
                <RESULT eventid="1474" points="461" reactiontime="+67" swimtime="00:01:07.22" resultid="11320" heatid="14037" lane="6" entrytime="00:01:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="11321" heatid="14049" lane="3" entrytime="00:02:32.00" />
                <RESULT eventid="1647" points="395" reactiontime="+68" swimtime="00:02:32.53" resultid="11322" heatid="14082" lane="0" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:13.32" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="11277">
              <RESULTS>
                <RESULT eventid="1079" points="356" reactiontime="+86" swimtime="00:00:29.48" resultid="11278" heatid="13911" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1165" points="315" reactiontime="+93" swimtime="00:21:19.98" resultid="11279" heatid="13942" lane="3" entrytime="00:21:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:17.86" />
                    <SPLIT distance="200" swimtime="00:02:41.64" />
                    <SPLIT distance="300" swimtime="00:04:05.94" />
                    <SPLIT distance="350" swimtime="00:04:47.97" />
                    <SPLIT distance="400" swimtime="00:06:55.47" />
                    <SPLIT distance="450" swimtime="00:06:12.66" />
                    <SPLIT distance="500" swimtime="00:08:21.33" />
                    <SPLIT distance="550" swimtime="00:07:37.88" />
                    <SPLIT distance="650" swimtime="00:09:03.98" />
                    <SPLIT distance="750" swimtime="00:10:30.50" />
                    <SPLIT distance="800" swimtime="00:09:47.58" />
                    <SPLIT distance="850" swimtime="00:11:57.01" />
                    <SPLIT distance="900" swimtime="00:11:14.04" />
                    <SPLIT distance="1000" swimtime="00:12:40.96" />
                    <SPLIT distance="1050" swimtime="00:14:51.12" />
                    <SPLIT distance="1100" swimtime="00:14:08.24" />
                    <SPLIT distance="1200" swimtime="00:15:34.62" />
                    <SPLIT distance="1250" swimtime="00:16:18.16" />
                    <SPLIT distance="1300" swimtime="00:17:02.56" />
                    <SPLIT distance="1350" swimtime="00:17:45.86" />
                    <SPLIT distance="1450" swimtime="00:19:12.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="401" reactiontime="+64" swimtime="00:00:32.60" resultid="11280" heatid="13955" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1474" points="355" reactiontime="+73" swimtime="00:01:13.30" resultid="11281" heatid="14036" lane="2" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="302" reactiontime="+79" swimtime="00:02:46.66" resultid="11282" heatid="14081" lane="0" entrytime="00:02:43.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:19.71" />
                    <SPLIT distance="150" swimtime="00:02:02.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="333" reactiontime="+91" swimtime="00:05:17.47" resultid="11283" heatid="14111" lane="2" entrytime="00:05:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:14.17" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                    <SPLIT distance="200" swimtime="00:02:34.70" />
                    <SPLIT distance="250" swimtime="00:03:15.93" />
                    <SPLIT distance="300" swimtime="00:03:57.57" />
                    <SPLIT distance="350" swimtime="00:04:38.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" athleteid="11284">
              <RESULTS>
                <RESULT eventid="1062" points="320" swimtime="00:00:34.66" resultid="11285" heatid="13900" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1222" points="322" reactiontime="+83" swimtime="00:03:22.82" resultid="11286" heatid="13961" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:36.77" />
                    <SPLIT distance="150" swimtime="00:02:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="317" reactiontime="+81" swimtime="00:01:34.32" resultid="11287" heatid="14003" lane="8" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="241" reactiontime="+84" swimtime="00:00:39.21" resultid="11288" heatid="14015" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1664" points="325" swimtime="00:00:42.84" resultid="11289" heatid="14085" lane="6" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-07" firstname="Elżbieta" gender="F" lastname="Krakowiak" nation="POL" license="100115600356" athleteid="11337">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1256" points="517" reactiontime="+94" swimtime="00:01:04.86" resultid="11338" heatid="13975" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="484" reactiontime="+98" swimtime="00:02:23.83" resultid="11339" heatid="14043" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="456" reactiontime="+74" swimtime="00:05:09.52" resultid="11340" heatid="14105" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:50.61" />
                    <SPLIT distance="200" swimtime="00:02:29.74" />
                    <SPLIT distance="250" swimtime="00:03:09.34" />
                    <SPLIT distance="300" swimtime="00:03:49.55" />
                    <SPLIT distance="350" swimtime="00:04:29.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="11290">
              <RESULTS>
                <RESULT eventid="1147" points="217" swimtime="00:13:30.67" resultid="11291" heatid="13936" lane="1" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:32.02" />
                    <SPLIT distance="150" swimtime="00:02:20.48" />
                    <SPLIT distance="200" swimtime="00:03:10.98" />
                    <SPLIT distance="250" swimtime="00:04:02.32" />
                    <SPLIT distance="300" swimtime="00:04:53.28" />
                    <SPLIT distance="350" swimtime="00:05:45.14" />
                    <SPLIT distance="400" swimtime="00:06:37.25" />
                    <SPLIT distance="450" swimtime="00:07:29.32" />
                    <SPLIT distance="500" swimtime="00:08:20.69" />
                    <SPLIT distance="550" swimtime="00:09:13.10" />
                    <SPLIT distance="600" swimtime="00:10:04.49" />
                    <SPLIT distance="650" swimtime="00:10:57.04" />
                    <SPLIT distance="700" swimtime="00:11:48.95" />
                    <SPLIT distance="750" swimtime="00:12:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="174" reactiontime="+129" swimtime="00:00:48.41" resultid="11292" heatid="13945" lane="2" entrytime="00:00:51.00" />
                <RESULT eventid="1256" points="212" swimtime="00:01:27.28" resultid="11293" heatid="13971" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="165" reactiontime="+127" swimtime="00:01:45.83" resultid="11294" heatid="14029" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="173" reactiontime="+113" swimtime="00:03:42.42" resultid="11295" heatid="14074" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.59" />
                    <SPLIT distance="100" swimtime="00:01:47.76" />
                    <SPLIT distance="150" swimtime="00:02:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="214" swimtime="00:06:38.17" resultid="11296" heatid="14103" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:22.34" />
                    <SPLIT distance="200" swimtime="00:03:13.12" />
                    <SPLIT distance="250" swimtime="00:04:04.94" />
                    <SPLIT distance="300" swimtime="00:04:56.99" />
                    <SPLIT distance="350" swimtime="00:05:48.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" athleteid="11306">
              <RESULTS>
                <RESULT eventid="1062" points="192" reactiontime="+88" swimtime="00:00:41.10" resultid="11307" heatid="13897" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1096" points="147" reactiontime="+101" swimtime="00:03:58.48" resultid="11308" heatid="13919" lane="2" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                    <SPLIT distance="100" swimtime="00:02:00.97" />
                    <SPLIT distance="150" swimtime="00:03:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="141" reactiontime="+78" swimtime="00:00:51.89" resultid="11309" heatid="13945" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1324" points="86" reactiontime="+92" swimtime="00:04:35.49" resultid="11310" heatid="13990" lane="3" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.92" />
                    <SPLIT distance="100" swimtime="00:02:08.96" />
                    <SPLIT distance="150" swimtime="00:03:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="141" reactiontime="+97" swimtime="00:08:35.53" resultid="11311" heatid="14057" lane="5" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.37" />
                    <SPLIT distance="100" swimtime="00:02:03.81" />
                    <SPLIT distance="150" swimtime="00:03:10.59" />
                    <SPLIT distance="200" swimtime="00:04:18.47" />
                    <SPLIT distance="250" swimtime="00:05:26.01" />
                    <SPLIT distance="300" swimtime="00:06:33.81" />
                    <SPLIT distance="350" swimtime="00:07:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="128" reactiontime="+74" swimtime="00:04:05.82" resultid="11312" heatid="14073" lane="5" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.74" />
                    <SPLIT distance="100" swimtime="00:04:05.93" />
                    <SPLIT distance="150" swimtime="00:03:05.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-31" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" athleteid="11328">
              <RESULTS>
                <RESULT eventid="1079" points="428" reactiontime="+81" swimtime="00:00:27.74" resultid="11329" heatid="13912" lane="3" entrytime="00:00:28.11" />
                <RESULT eventid="1113" points="317" reactiontime="+88" swimtime="00:02:47.06" resultid="11330" heatid="13928" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="391" swimtime="00:02:53.61" resultid="11331" heatid="13965" lane="9" entrytime="00:03:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                    <SPLIT distance="150" swimtime="00:02:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="421" reactiontime="+82" swimtime="00:01:02.56" resultid="11332" heatid="13984" lane="2" entrytime="00:01:04.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="436" reactiontime="+78" swimtime="00:01:16.33" resultid="11333" heatid="14011" lane="8" entrytime="00:01:19.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="344" swimtime="00:00:32.01" resultid="11334" heatid="14025" lane="9" entrytime="00:00:30.98" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="11335" heatid="14066" lane="5" entrytime="00:01:59.99" />
                <RESULT eventid="1681" points="462" reactiontime="+81" swimtime="00:00:34.16" resultid="11336" heatid="14096" lane="8" entrytime="00:00:35.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-03" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="11341">
              <RESULTS>
                <RESULT eventid="1273" points="421" swimtime="00:01:02.57" resultid="11342" heatid="13986" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="372" reactiontime="+77" swimtime="00:02:21.77" resultid="11343" heatid="14052" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="396" swimtime="00:04:59.68" resultid="11344" heatid="14113" lane="9" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:51.35" />
                    <SPLIT distance="200" swimtime="00:02:30.84" />
                    <SPLIT distance="250" swimtime="00:03:09.37" />
                    <SPLIT distance="300" swimtime="00:03:47.47" />
                    <SPLIT distance="350" swimtime="00:04:24.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="11270">
              <RESULTS>
                <RESULT eventid="1165" points="181" reactiontime="+105" swimtime="00:25:37.49" resultid="11271" heatid="13940" lane="4" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:21.64" />
                    <SPLIT distance="200" swimtime="00:03:12.32" />
                    <SPLIT distance="250" swimtime="00:04:04.01" />
                    <SPLIT distance="300" swimtime="00:04:55.05" />
                    <SPLIT distance="350" swimtime="00:05:47.05" />
                    <SPLIT distance="400" swimtime="00:06:38.41" />
                    <SPLIT distance="450" swimtime="00:07:29.90" />
                    <SPLIT distance="500" swimtime="00:08:22.32" />
                    <SPLIT distance="550" swimtime="00:09:13.73" />
                    <SPLIT distance="600" swimtime="00:10:05.84" />
                    <SPLIT distance="650" swimtime="00:10:57.74" />
                    <SPLIT distance="700" swimtime="00:11:49.61" />
                    <SPLIT distance="750" swimtime="00:12:41.89" />
                    <SPLIT distance="800" swimtime="00:13:34.03" />
                    <SPLIT distance="850" swimtime="00:14:26.06" />
                    <SPLIT distance="900" swimtime="00:15:18.25" />
                    <SPLIT distance="950" swimtime="00:16:10.02" />
                    <SPLIT distance="1000" swimtime="00:17:02.22" />
                    <SPLIT distance="1050" swimtime="00:17:54.26" />
                    <SPLIT distance="1100" swimtime="00:18:46.21" />
                    <SPLIT distance="1150" swimtime="00:19:38.22" />
                    <SPLIT distance="1200" swimtime="00:20:29.92" />
                    <SPLIT distance="1250" swimtime="00:21:21.45" />
                    <SPLIT distance="1300" swimtime="00:22:13.90" />
                    <SPLIT distance="1350" swimtime="00:23:05.57" />
                    <SPLIT distance="1400" swimtime="00:23:57.77" />
                    <SPLIT distance="1450" swimtime="00:24:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="188" reactiontime="+101" swimtime="00:03:14.61" resultid="11272" heatid="13994" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:33.50" />
                    <SPLIT distance="150" swimtime="00:02:23.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="187" reactiontime="+104" swimtime="00:00:39.21" resultid="11273" heatid="14020" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1508" points="198" reactiontime="+104" swimtime="00:02:54.82" resultid="11274" heatid="14047" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="150" swimtime="00:02:11.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="197" reactiontime="+111" swimtime="00:01:25.55" resultid="11275" heatid="14068" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="132" reactiontime="+85" swimtime="00:03:39.38" resultid="11276" heatid="14078" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                    <SPLIT distance="100" swimtime="00:01:51.49" />
                    <SPLIT distance="150" swimtime="00:02:49.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="11323">
              <RESULTS>
                <RESULT eventid="1113" points="254" reactiontime="+87" swimtime="00:02:59.86" resultid="11324" heatid="13925" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:19.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="307" reactiontime="+89" swimtime="00:03:08.19" resultid="11325" heatid="13967" lane="7" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                    <SPLIT distance="150" swimtime="00:02:18.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="296" reactiontime="+83" swimtime="00:01:26.83" resultid="11326" heatid="14008" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="313" reactiontime="+90" swimtime="00:00:38.88" resultid="11327" heatid="14091" lane="1" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="11297">
              <RESULTS>
                <RESULT eventid="1113" points="526" reactiontime="+79" swimtime="00:02:21.19" resultid="11298" heatid="13931" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1165" points="526" reactiontime="+79" swimtime="00:17:58.35" resultid="11299" heatid="13943" lane="5" entrytime="00:18:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.36" />
                    <SPLIT distance="200" swimtime="00:02:18.12" />
                    <SPLIT distance="250" swimtime="00:02:53.76" />
                    <SPLIT distance="300" swimtime="00:03:29.56" />
                    <SPLIT distance="350" swimtime="00:04:05.50" />
                    <SPLIT distance="400" swimtime="00:04:41.64" />
                    <SPLIT distance="450" swimtime="00:05:17.88" />
                    <SPLIT distance="500" swimtime="00:05:54.34" />
                    <SPLIT distance="550" swimtime="00:06:30.65" />
                    <SPLIT distance="600" swimtime="00:07:07.03" />
                    <SPLIT distance="650" swimtime="00:07:43.56" />
                    <SPLIT distance="700" swimtime="00:08:19.97" />
                    <SPLIT distance="750" swimtime="00:08:56.28" />
                    <SPLIT distance="800" swimtime="00:09:32.32" />
                    <SPLIT distance="850" swimtime="00:10:09.08" />
                    <SPLIT distance="900" swimtime="00:10:45.86" />
                    <SPLIT distance="950" swimtime="00:11:22.41" />
                    <SPLIT distance="1000" swimtime="00:11:59.41" />
                    <SPLIT distance="1050" swimtime="00:12:35.92" />
                    <SPLIT distance="1100" swimtime="00:13:11.89" />
                    <SPLIT distance="1150" swimtime="00:13:47.82" />
                    <SPLIT distance="1200" swimtime="00:14:23.78" />
                    <SPLIT distance="1250" swimtime="00:15:00.03" />
                    <SPLIT distance="1300" swimtime="00:15:36.13" />
                    <SPLIT distance="1350" swimtime="00:16:12.25" />
                    <SPLIT distance="1400" swimtime="00:16:48.28" />
                    <SPLIT distance="1450" swimtime="00:17:24.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="462" reactiontime="+76" swimtime="00:02:44.26" resultid="11300" heatid="13970" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="504" reactiontime="+76" swimtime="00:02:20.07" resultid="11301" heatid="13995" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="534" reactiontime="+73" swimtime="00:02:05.70" resultid="11302" heatid="14053" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="100" swimtime="00:01:01.00" />
                    <SPLIT distance="150" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="473" reactiontime="+80" swimtime="00:05:12.74" resultid="11303" heatid="14062" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:50.18" />
                    <SPLIT distance="200" swimtime="00:02:32.10" />
                    <SPLIT distance="250" swimtime="00:03:16.29" />
                    <SPLIT distance="300" swimtime="00:04:01.57" />
                    <SPLIT distance="350" swimtime="00:04:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="511" reactiontime="+76" swimtime="00:01:02.31" resultid="11304" heatid="14071" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="532" reactiontime="+79" swimtime="00:04:31.50" resultid="11305" heatid="14114" lane="3" entrytime="00:04:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="150" swimtime="00:01:39.16" />
                    <SPLIT distance="200" swimtime="00:02:13.65" />
                    <SPLIT distance="250" swimtime="00:02:48.12" />
                    <SPLIT distance="300" swimtime="00:03:22.80" />
                    <SPLIT distance="350" swimtime="00:03:57.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-28" firstname="Łukasz" gender="M" lastname="Stolarczyk" nation="POL" athleteid="11313">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="11314" heatid="13989" lane="9" entrytime="00:00:57.30" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="11315" heatid="14027" lane="9" entrytime="00:00:27.90" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="11316" heatid="14071" lane="8" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="KS WARTA POZNAŃ ZMIENNA MĘSKA" number="2">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="11346" heatid="13999" lane="6" entrytime="00:02:02.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11317" number="1" />
                    <RELAYPOSITION athleteid="11328" number="2" />
                    <RELAYPOSITION athleteid="11313" number="3" />
                    <RELAYPOSITION athleteid="11297" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="KS WARTA POZNAŃ ZMIENNA MĘSKA" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="275" reactiontime="+83" swimtime="00:02:23.63" resultid="11347" heatid="13998" lane="0" entrytime="00:02:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:54.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11277" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="11323" number="2" />
                    <RELAYPOSITION athleteid="11270" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="11341" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="KS WARTA POZNAŃ ZMIENNA PAŃ" number="4">
              <RESULTS>
                <RESULT eventid="1358" points="228" reactiontime="+121" swimtime="00:02:53.78" resultid="11348" heatid="13996" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.32" />
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                    <SPLIT distance="150" swimtime="00:02:24.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11290" number="1" reactiontime="+121" />
                    <RELAYPOSITION athleteid="11284" number="2" />
                    <RELAYPOSITION athleteid="11306" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="11337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="KS WARTA POZNAŃ DOWOLNA MIXED" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="227" swimtime="00:02:18.91" resultid="11345" heatid="13933" lane="1" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:49.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11290" number="1" />
                    <RELAYPOSITION athleteid="11323" number="2" />
                    <RELAYPOSITION athleteid="11284" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="11277" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="KS WARTA POZNAŃ ZMIENNA MIXED" number="5">
              <RESULTS>
                <RESULT eventid="1698" points="355" reactiontime="+74" swimtime="00:02:11.83" resultid="11349" heatid="14101" lane="0" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:42.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11317" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="11284" number="2" />
                    <RELAYPOSITION athleteid="11297" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="11337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="KS WARTA POZNAŃ ZMIENNA MIXED" number="6">
              <RESULTS>
                <RESULT eventid="1698" points="168" reactiontime="+89" swimtime="00:02:49.28" resultid="11350" heatid="14100" lane="9" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:29.10" />
                    <SPLIT distance="150" swimtime="00:02:18.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11290" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="11323" number="2" />
                    <RELAYPOSITION athleteid="11306" number="3" />
                    <RELAYPOSITION athleteid="11277" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="WAR" clubid="11648" name="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="11649">
              <RESULTS>
                <RESULT eventid="1079" points="524" reactiontime="+86" swimtime="00:00:25.92" resultid="11650" heatid="13917" lane="1" entrytime="00:00:25.50" />
                <RESULT comment="Rekord Polski" eventid="1205" points="630" reactiontime="+64" swimtime="00:00:28.03" resultid="11651" heatid="13958" lane="4" entrytime="00:00:28.25" />
                <RESULT eventid="1440" points="627" reactiontime="+77" swimtime="00:00:26.20" resultid="11652" heatid="14018" lane="4" />
                <RESULT comment="Rekord Polski" eventid="1474" points="601" reactiontime="+62" swimtime="00:01:01.52" resultid="11653" heatid="14038" lane="4" entrytime="00:01:01.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="534" reactiontime="+63" swimtime="00:02:17.92" resultid="11654" heatid="14082" lane="4" entrytime="00:02:17.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="150" swimtime="00:01:41.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="11655">
              <RESULTS>
                <RESULT eventid="1062" points="503" reactiontime="+80" swimtime="00:00:29.82" resultid="11656" heatid="13902" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1096" points="447" reactiontime="+88" swimtime="00:02:44.89" resultid="11657" heatid="13921" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:02:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1187" points="526" reactiontime="+73" swimtime="00:00:33.52" resultid="11658" heatid="13948" lane="4" entrytime="00:00:32.50" />
                <RESULT comment="Rekord Polski" eventid="1457" points="493" reactiontime="+76" swimtime="00:01:13.56" resultid="11659" heatid="14031" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="390" swimtime="00:02:34.53" resultid="11660" heatid="14043" lane="6" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1630" points="465" reactiontime="+77" swimtime="00:02:40.04" resultid="11661" heatid="14075" lane="4" entrytime="00:02:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:01:59.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="383" reactiontime="+93" swimtime="00:05:28.19" resultid="11662" heatid="14105" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="200" swimtime="00:02:36.64" />
                    <SPLIT distance="300" swimtime="00:04:03.57" />
                    <SPLIT distance="350" swimtime="00:04:47.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="12483" name="MAREA klub Košice">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1991-03-13" firstname="Peter" gender="M" lastname="Hrinda" nation="SVK" athleteid="12484">
              <RESULTS>
                <RESULT eventid="1681" points="651" reactiontime="+72" swimtime="00:00:30.48" resultid="12485" heatid="14098" lane="5" entrytime="00:00:29.92" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10084" name="Masters Białystok">
          <CONTACT city="Białystok" email="epiwo@wp.pl" name="Piwowarczyk" phone="600330566" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="10085">
              <RESULTS>
                <RESULT eventid="1147" points="408" reactiontime="+87" swimtime="00:10:56.85" resultid="10086" heatid="13937" lane="4" entrytime="00:10:24.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:55.01" />
                    <SPLIT distance="200" swimtime="00:02:35.53" />
                    <SPLIT distance="250" swimtime="00:03:16.03" />
                    <SPLIT distance="300" swimtime="00:03:56.53" />
                    <SPLIT distance="350" swimtime="00:04:37.50" />
                    <SPLIT distance="400" swimtime="00:05:18.40" />
                    <SPLIT distance="450" swimtime="00:05:59.69" />
                    <SPLIT distance="500" swimtime="00:06:40.83" />
                    <SPLIT distance="550" swimtime="00:07:21.69" />
                    <SPLIT distance="600" swimtime="00:08:04.76" />
                    <SPLIT distance="650" swimtime="00:08:47.98" />
                    <SPLIT distance="700" swimtime="00:09:31.71" />
                    <SPLIT distance="750" swimtime="00:10:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="458" reactiontime="+85" swimtime="00:01:07.53" resultid="10087" heatid="13976" lane="2" entrytime="00:01:05.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="467" reactiontime="+86" swimtime="00:02:25.56" resultid="10088" heatid="14043" lane="7" entrytime="00:02:22.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="443" reactiontime="+84" swimtime="00:05:12.52" resultid="10089" heatid="14105" lane="4" entrytime="00:05:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:51.07" />
                    <SPLIT distance="200" swimtime="00:02:31.18" />
                    <SPLIT distance="250" swimtime="00:03:11.31" />
                    <SPLIT distance="300" swimtime="00:03:52.16" />
                    <SPLIT distance="350" swimtime="00:04:33.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12424" name="Masters Team Biała Podlaska">
          <CONTACT city="Biała Podlaska" email="wilhelmg@poczta.onet.pl" name="Gromisz" zip="21-500" />
          <ATHLETES>
            <ATHLETE birthdate="1990-09-04" firstname="Krzysztof" gender="M" lastname="Rola" nation="POL" athleteid="12449">
              <RESULTS>
                <RESULT eventid="1079" points="484" swimtime="00:00:26.62" resultid="12450" heatid="13917" lane="9" entrytime="00:00:25.78" />
                <RESULT eventid="1205" points="442" reactiontime="+68" swimtime="00:00:31.55" resultid="12451" heatid="13957" lane="6" entrytime="00:00:31.20" />
                <RESULT eventid="1273" points="458" reactiontime="+72" swimtime="00:01:00.85" resultid="12452" heatid="13987" lane="1" entrytime="00:00:59.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="494" swimtime="00:00:28.37" resultid="12453" heatid="14026" lane="9" entrytime="00:00:29.12" />
                <RESULT eventid="1474" points="403" swimtime="00:01:10.28" resultid="12454" heatid="14037" lane="7" entrytime="00:01:10.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-11-29" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="12425">
              <RESULTS>
                <RESULT eventid="1062" points="498" reactiontime="+84" swimtime="00:00:29.92" resultid="12426" heatid="13901" lane="4" entrytime="00:00:31.05" />
                <RESULT eventid="1096" points="410" reactiontime="+87" swimtime="00:02:49.67" resultid="12427" heatid="13921" lane="1" entrytime="00:02:49.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:02:08.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="467" reactiontime="+100" swimtime="00:01:07.07" resultid="12428" heatid="13975" lane="6" entrytime="00:01:09.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="273" reactiontime="+95" swimtime="00:03:07.63" resultid="12429" heatid="13991" lane="6" entrytime="00:03:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:18.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="462" swimtime="00:00:31.60" resultid="12430" heatid="14017" lane="6" entrytime="00:00:32.20" />
                <RESULT eventid="1555" points="343" reactiontime="+105" swimtime="00:06:23.37" resultid="12431" heatid="14058" lane="3" entrytime="00:06:04.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="150" swimtime="00:02:14.97" />
                    <SPLIT distance="200" swimtime="00:03:05.72" />
                    <SPLIT distance="250" swimtime="00:03:57.86" />
                    <SPLIT distance="300" swimtime="00:04:52.91" />
                    <SPLIT distance="350" swimtime="00:05:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="417" reactiontime="+87" swimtime="00:01:14.44" resultid="12432" heatid="14065" lane="2" entrytime="00:01:16.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="340" reactiontime="+91" swimtime="00:05:41.22" resultid="12433" heatid="14105" lane="7" entrytime="00:05:12.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                    <SPLIT distance="200" swimtime="00:02:45.34" />
                    <SPLIT distance="250" swimtime="00:03:29.89" />
                    <SPLIT distance="300" swimtime="00:04:14.49" />
                    <SPLIT distance="350" swimtime="00:04:58.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Michał" gender="M" lastname="Jagiełło" nation="POL" athleteid="12442">
              <RESULTS>
                <RESULT eventid="1079" points="584" reactiontime="+79" swimtime="00:00:25.01" resultid="12443" heatid="13917" lane="2" entrytime="00:00:25.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="560" reactiontime="+81" swimtime="00:00:56.88" resultid="12444" heatid="13987" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="516" reactiontime="+77" swimtime="00:00:27.96" resultid="12445" heatid="14026" lane="3" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-07" firstname="Robert" gender="M" lastname="Jagiełło" nation="POL" athleteid="12446">
              <RESULTS>
                <RESULT eventid="1079" points="201" reactiontime="+101" swimtime="00:00:35.69" resultid="12447" heatid="13907" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1273" points="137" reactiontime="+95" swimtime="00:01:30.90" resultid="12448" heatid="13980" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-27" firstname="Renata" gender="F" lastname="Kasprowicz" nation="POL" athleteid="12434">
              <RESULTS>
                <RESULT eventid="1062" points="445" reactiontime="+87" swimtime="00:00:31.06" resultid="12435" heatid="13901" lane="2" entrytime="00:00:31.85" />
                <RESULT eventid="1096" points="288" reactiontime="+84" swimtime="00:03:10.97" resultid="12436" heatid="13920" lane="8" entrytime="00:03:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:25.39" />
                    <SPLIT distance="150" swimtime="00:02:20.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="325" reactiontime="+81" swimtime="00:03:22.19" resultid="12437" heatid="13962" lane="7" entrytime="00:03:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:34.82" />
                    <SPLIT distance="150" swimtime="00:02:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="350" reactiontime="+93" swimtime="00:01:13.87" resultid="12438" heatid="13975" lane="0" entrytime="00:01:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="346" reactiontime="+87" swimtime="00:01:31.66" resultid="12439" heatid="14003" lane="6" entrytime="00:01:31.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="356" reactiontime="+80" swimtime="00:00:34.46" resultid="12440" heatid="14017" lane="7" entrytime="00:00:32.78" />
                <RESULT eventid="1664" points="374" swimtime="00:00:40.90" resultid="12441" heatid="14086" lane="6" entrytime="00:00:40.26" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="10892" name="Masters Unia Oświęcim">
          <ATHLETES>
            <ATHLETE birthdate="1969-11-05" firstname="Sławomir" gender="M" lastname="Formas" nation="POL" athleteid="10897">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1239" points="499" reactiontime="+82" swimtime="00:02:40.08" resultid="10898" heatid="13969" lane="4" entrytime="00:02:47.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1406" points="530" reactiontime="+76" swimtime="00:01:11.55" resultid="10899" heatid="14013" lane="8" entrytime="00:01:13.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="368" reactiontime="+80" swimtime="00:02:22.28" resultid="10900" heatid="14052" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1681" points="549" swimtime="00:00:32.26" resultid="10901" heatid="14098" lane="9" entrytime="00:00:32.52" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" nation="POL" athleteid="10906">
              <RESULTS>
                <RESULT eventid="1256" points="330" reactiontime="+89" swimtime="00:01:15.29" resultid="10907" heatid="13974" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="292" reactiontime="+98" swimtime="00:01:36.91" resultid="10908" heatid="14002" lane="2" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="287" reactiontime="+92" swimtime="00:02:51.14" resultid="10909" heatid="14041" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:21.52" />
                    <SPLIT distance="150" swimtime="00:02:06.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="289" reactiontime="+84" swimtime="00:00:44.57" resultid="10910" heatid="14086" lane="8" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="10893">
              <RESULTS>
                <RESULT eventid="1205" points="263" reactiontime="+68" swimtime="00:00:37.49" resultid="10894" heatid="13953" lane="4" entrytime="00:00:38.05" />
                <RESULT eventid="1474" points="242" reactiontime="+83" swimtime="00:01:23.33" resultid="10895" heatid="14035" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="220" reactiontime="+70" swimtime="00:03:05.14" resultid="10896" heatid="14079" lane="4" entrytime="00:03:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:16.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" athleteid="10902">
              <RESULTS>
                <RESULT eventid="1187" points="352" reactiontime="+80" swimtime="00:00:38.31" resultid="10903" heatid="13947" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1457" points="325" reactiontime="+76" swimtime="00:01:24.53" resultid="10904" heatid="14030" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="292" reactiontime="+82" swimtime="00:03:06.93" resultid="10905" heatid="14074" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:22.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" points="264" reactiontime="+77" swimtime="00:02:25.61" resultid="11546" heatid="14101" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:22.45" />
                    <SPLIT distance="150" swimtime="00:01:51.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10893" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="10897" number="2" />
                    <RELAYPOSITION athleteid="10902" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="10906" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="10367" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="10425">
              <RESULTS>
                <RESULT eventid="1079" points="441" reactiontime="+71" swimtime="00:00:27.46" resultid="10426" heatid="13914" lane="8" entrytime="00:00:27.30" entrycourse="LCM" />
                <RESULT eventid="1113" points="379" reactiontime="+88" swimtime="00:02:37.40" resultid="10427" heatid="13929" lane="7" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:15.67" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="10428" heatid="13968" lane="4" entrytime="00:02:55.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="450" reactiontime="+79" swimtime="00:01:01.21" resultid="10429" heatid="13986" lane="5" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="405" reactiontime="+78" swimtime="00:01:18.28" resultid="10430" heatid="14012" lane="9" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="311" reactiontime="+109" swimtime="00:05:59.90" resultid="10431" heatid="14061" lane="2" entrytime="00:05:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:24.73" />
                    <SPLIT distance="150" swimtime="00:02:12.12" />
                    <SPLIT distance="200" swimtime="00:02:58.57" />
                    <SPLIT distance="250" swimtime="00:03:51.20" />
                    <SPLIT distance="300" swimtime="00:04:42.79" />
                    <SPLIT distance="350" swimtime="00:05:22.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="470" reactiontime="+81" swimtime="00:00:33.96" resultid="10432" heatid="14096" lane="7" entrytime="00:00:35.50" entrycourse="LCM" />
                <RESULT eventid="1744" points="342" reactiontime="+65" swimtime="00:05:14.55" resultid="10433" heatid="14112" lane="6" entrytime="00:05:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:52.06" />
                    <SPLIT distance="200" swimtime="00:02:32.98" />
                    <SPLIT distance="250" swimtime="00:03:13.68" />
                    <SPLIT distance="300" swimtime="00:03:55.38" />
                    <SPLIT distance="350" swimtime="00:04:36.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" athleteid="10388">
              <RESULTS>
                <RESULT eventid="1113" points="135" swimtime="00:03:41.95" resultid="10389" heatid="13924" lane="9" entrytime="00:03:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:57.05" />
                    <SPLIT distance="150" swimtime="00:02:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="225" reactiontime="+112" swimtime="00:03:28.60" resultid="10390" heatid="13966" lane="0" entrytime="00:03:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.09" />
                    <SPLIT distance="100" swimtime="00:01:43.09" />
                    <SPLIT distance="150" swimtime="00:02:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="253" reactiontime="+100" swimtime="00:01:31.51" resultid="10391" heatid="14008" lane="7" entrytime="00:01:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="333" reactiontime="+93" swimtime="00:00:38.08" resultid="10392" heatid="14093" lane="8" entrytime="00:00:39.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-27" firstname="Michał" gender="M" lastname="Klupa" nation="POL" athleteid="10475">
              <RESULTS>
                <RESULT eventid="1205" points="542" reactiontime="+57" swimtime="00:00:29.47" resultid="10476" heatid="13958" lane="5" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1474" points="471" reactiontime="+62" swimtime="00:01:06.72" resultid="10477" heatid="14038" lane="3" entrytime="00:01:02.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="397" reactiontime="+79" swimtime="00:05:31.74" resultid="10478" heatid="14061" lane="3" entrytime="00:05:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:13.75" />
                    <SPLIT distance="200" swimtime="00:02:36.70" />
                    <SPLIT distance="250" swimtime="00:03:26.04" />
                    <SPLIT distance="300" swimtime="00:04:15.98" />
                    <SPLIT distance="350" swimtime="00:04:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="457" reactiontime="+61" swimtime="00:02:25.26" resultid="10479" heatid="14082" lane="5" entrytime="00:02:18.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:48.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="412" reactiontime="+70" swimtime="00:04:55.53" resultid="10480" heatid="14112" lane="5" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:06.19" />
                    <SPLIT distance="150" swimtime="00:01:43.49" />
                    <SPLIT distance="200" swimtime="00:02:21.18" />
                    <SPLIT distance="250" swimtime="00:02:59.74" />
                    <SPLIT distance="300" swimtime="00:03:38.54" />
                    <SPLIT distance="350" swimtime="00:04:18.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="10517">
              <RESULTS>
                <RESULT eventid="1062" points="456" reactiontime="+77" swimtime="00:00:30.81" resultid="10518" heatid="13901" lane="3" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1147" points="353" reactiontime="+83" swimtime="00:11:29.38" resultid="10519" heatid="13937" lane="1" entrytime="00:11:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:16.98" />
                    <SPLIT distance="150" swimtime="00:01:59.99" />
                    <SPLIT distance="200" swimtime="00:02:43.97" />
                    <SPLIT distance="250" swimtime="00:03:28.14" />
                    <SPLIT distance="300" swimtime="00:04:12.33" />
                    <SPLIT distance="350" swimtime="00:04:56.83" />
                    <SPLIT distance="400" swimtime="00:05:41.39" />
                    <SPLIT distance="450" swimtime="00:06:25.84" />
                    <SPLIT distance="500" swimtime="00:07:09.34" />
                    <SPLIT distance="550" swimtime="00:07:54.27" />
                    <SPLIT distance="600" swimtime="00:08:37.93" />
                    <SPLIT distance="650" swimtime="00:09:22.27" />
                    <SPLIT distance="700" swimtime="00:10:05.78" />
                    <SPLIT distance="750" swimtime="00:10:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="460" reactiontime="+64" swimtime="00:00:35.04" resultid="10520" heatid="13948" lane="2" entrytime="00:00:34.50" entrycourse="LCM" />
                <RESULT eventid="1324" points="273" reactiontime="+80" swimtime="00:03:07.75" resultid="10521" heatid="13990" lane="4" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:17.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="449" reactiontime="+73" swimtime="00:01:15.88" resultid="10522" heatid="14031" lane="2" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="366" swimtime="00:02:37.93" resultid="10523" heatid="14043" lane="9" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:57.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="409" reactiontime="+64" swimtime="00:02:47.09" resultid="10524" heatid="14075" lane="2" entrytime="00:02:44.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="378" swimtime="00:05:29.44" resultid="10525" heatid="14105" lane="9" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:00.06" />
                    <SPLIT distance="200" swimtime="00:02:43.47" />
                    <SPLIT distance="250" swimtime="00:03:25.57" />
                    <SPLIT distance="300" swimtime="00:04:08.07" />
                    <SPLIT distance="350" swimtime="00:04:50.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-12" firstname="Janusz" gender="M" lastname="Mrozik" nation="POL" athleteid="10540">
              <RESULTS>
                <RESULT eventid="1239" points="63" swimtime="00:05:19.19" resultid="10541" heatid="13964" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.15" />
                    <SPLIT distance="100" swimtime="00:02:37.30" />
                    <SPLIT distance="150" swimtime="00:03:59.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="41" reactiontime="+115" swimtime="00:02:15.42" resultid="10542" heatid="13977" lane="5" entrytime="00:02:06.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Karolina" gender="F" lastname="Górka" nation="POL" athleteid="10496">
              <RESULTS>
                <RESULT eventid="1062" points="442" reactiontime="+69" swimtime="00:00:31.13" resultid="10497" heatid="13901" lane="6" entrytime="00:00:31.74" entrycourse="LCM" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="10498" heatid="13921" lane="8" entrytime="00:02:50.00" entrycourse="LCM" />
                <RESULT eventid="1222" points="349" reactiontime="+74" swimtime="00:03:17.41" resultid="10499" heatid="13961" lane="8" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:33.76" />
                    <SPLIT distance="150" swimtime="00:02:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="391" reactiontime="+73" swimtime="00:01:11.20" resultid="10500" heatid="13975" lane="7" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="348" reactiontime="+72" swimtime="00:01:31.41" resultid="10501" heatid="14004" lane="9" entrytime="00:01:28.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="282" reactiontime="+78" swimtime="00:02:52.14" resultid="10502" heatid="14042" lane="2" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="362" reactiontime="+70" swimtime="00:00:41.36" resultid="10503" heatid="14086" lane="7" entrytime="00:00:41.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="10414">
              <RESULTS>
                <RESULT eventid="1062" points="117" reactiontime="+129" swimtime="00:00:48.43" resultid="10415" heatid="13896" lane="4" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="108" reactiontime="+80" swimtime="00:00:56.66" resultid="10416" heatid="13944" lane="5" entrytime="00:00:57.00" entrycourse="LCM" />
                <RESULT eventid="1222" points="123" reactiontime="+122" swimtime="00:04:38.97" resultid="10417" heatid="13960" lane="0" entrytime="00:04:30.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.26" />
                    <SPLIT distance="100" swimtime="00:02:15.31" />
                    <SPLIT distance="150" swimtime="00:03:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="113" reactiontime="+75" swimtime="00:02:00.13" resultid="10418" heatid="14029" lane="9" entrytime="00:02:05.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="113" reactiontime="+93" swimtime="00:04:16.25" resultid="10419" heatid="14073" lane="7" entrytime="00:04:26.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.56" />
                    <SPLIT distance="100" swimtime="00:02:07.08" />
                    <SPLIT distance="150" swimtime="00:03:13.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="10490">
              <RESULTS>
                <RESULT eventid="1079" points="487" reactiontime="+73" swimtime="00:00:26.56" resultid="10491" heatid="13915" lane="3" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1273" points="460" reactiontime="+75" swimtime="00:01:00.75" resultid="10492" heatid="13987" lane="8" entrytime="00:00:59.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="10493" heatid="14025" lane="3" entrytime="00:00:29.69" entrycourse="LCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="10494" heatid="14051" lane="0" entrytime="00:02:20.69" entrycourse="LCM" />
                <RESULT eventid="1681" points="441" reactiontime="+76" swimtime="00:00:34.70" resultid="10495" heatid="14093" lane="7" entrytime="00:00:38.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="10420">
              <RESULTS>
                <RESULT eventid="1222" points="534" reactiontime="+81" swimtime="00:02:51.46" resultid="10421" heatid="13962" lane="4" entrytime="00:02:48.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:05.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="596" reactiontime="+81" swimtime="00:01:01.85" resultid="10422" heatid="13976" lane="4" entrytime="00:01:01.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="526" reactiontime="+82" swimtime="00:01:19.67" resultid="10423" heatid="14004" lane="4" entrytime="00:01:18.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="577" reactiontime="+83" swimtime="00:02:15.70" resultid="10424" heatid="14043" lane="4" entrytime="00:02:13.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="150" swimtime="00:01:40.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="10510">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1079" points="124" reactiontime="+116" swimtime="00:00:41.87" resultid="10511" heatid="13905" lane="5" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="76" reactiontime="+126" swimtime="00:04:28.79" resultid="10512" heatid="13923" lane="1" entrytime="00:04:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.17" />
                    <SPLIT distance="100" swimtime="00:02:19.01" />
                    <SPLIT distance="150" swimtime="00:03:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1205" points="69" reactiontime="+88" swimtime="00:00:58.36" resultid="10513" heatid="13950" lane="8" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="97" reactiontime="+127" swimtime="00:01:41.88" resultid="10514" heatid="13978" lane="5" entrytime="00:01:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="86" reactiontime="+122" swimtime="00:03:50.89" resultid="10515" heatid="14045" lane="4" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.88" />
                    <SPLIT distance="150" swimtime="00:02:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="88" swimtime="00:00:59.39" resultid="10516" heatid="14089" lane="9" entrytime="00:00:58.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="10393">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="10394" heatid="13926" lane="8" entrytime="00:03:00.00" entrycourse="LCM" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="10395" heatid="13965" lane="7" entrytime="00:03:50.00" entrycourse="LCM" />
                <RESULT eventid="1341" points="142" reactiontime="+93" swimtime="00:03:33.29" resultid="10396" heatid="13994" lane="2" entrytime="00:03:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:30.96" />
                    <SPLIT distance="150" swimtime="00:02:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="257" reactiontime="+95" swimtime="00:01:31.03" resultid="10397" heatid="14009" lane="0" entrytime="00:01:25.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="10398" heatid="14068" lane="5" entrytime="00:01:24.80" entrycourse="LCM" />
                <RESULT eventid="1681" points="287" reactiontime="+88" swimtime="00:00:40.02" resultid="10399" heatid="14093" lane="3" entrytime="00:00:38.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="10504">
              <RESULTS>
                <RESULT eventid="1079" points="67" reactiontime="+120" swimtime="00:00:51.44" resultid="10505" heatid="13904" lane="1" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1205" points="67" reactiontime="+65" swimtime="00:00:58.96" resultid="10506" heatid="13950" lane="1" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="62" reactiontime="+98" swimtime="00:01:58.38" resultid="10507" heatid="13977" lane="4" entrytime="00:01:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="61" reactiontime="+73" swimtime="00:02:11.72" resultid="10508" heatid="14033" lane="0" entrytime="00:02:06.00" entrycourse="LCM" />
                <RESULT eventid="1647" points="39" reactiontime="+62" swimtime="00:05:28.25" resultid="10509" heatid="14077" lane="2" entrytime="00:04:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.43" />
                    <SPLIT distance="100" swimtime="00:04:47.45" />
                    <SPLIT distance="150" swimtime="00:03:34.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-22" firstname="Mateusz" gender="M" lastname="Dybek" nation="POL" athleteid="10534">
              <RESULTS>
                <RESULT eventid="1079" points="470" swimtime="00:00:26.88" resultid="10535" heatid="13916" lane="9" entrytime="00:00:26.30" entrycourse="LCM" />
                <RESULT comment="(Time: 21:07), Przekroczony regulaminowy limit czasu." eventid="1165" status="OTL" swimtime="00:21:38.60" resultid="10536" heatid="13942" lane="6" entrytime="00:21:11.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="150" swimtime="00:01:57.04" />
                    <SPLIT distance="200" swimtime="00:02:39.30" />
                    <SPLIT distance="250" swimtime="00:03:21.56" />
                    <SPLIT distance="300" swimtime="00:04:04.85" />
                    <SPLIT distance="350" swimtime="00:04:47.91" />
                    <SPLIT distance="400" swimtime="00:05:31.61" />
                    <SPLIT distance="450" swimtime="00:06:14.82" />
                    <SPLIT distance="500" swimtime="00:06:58.85" />
                    <SPLIT distance="550" swimtime="00:07:41.93" />
                    <SPLIT distance="600" swimtime="00:08:26.22" />
                    <SPLIT distance="650" swimtime="00:09:10.19" />
                    <SPLIT distance="700" swimtime="00:09:54.92" />
                    <SPLIT distance="750" swimtime="00:10:38.94" />
                    <SPLIT distance="800" swimtime="00:11:23.74" />
                    <SPLIT distance="850" swimtime="00:12:06.54" />
                    <SPLIT distance="900" swimtime="00:12:50.42" />
                    <SPLIT distance="950" swimtime="00:13:33.83" />
                    <SPLIT distance="1000" swimtime="00:14:17.60" />
                    <SPLIT distance="1050" swimtime="00:15:01.18" />
                    <SPLIT distance="1100" swimtime="00:15:45.17" />
                    <SPLIT distance="1150" swimtime="00:16:29.17" />
                    <SPLIT distance="1200" swimtime="00:17:13.88" />
                    <SPLIT distance="1250" swimtime="00:17:58.09" />
                    <SPLIT distance="1300" swimtime="00:18:42.50" />
                    <SPLIT distance="1350" swimtime="00:19:27.04" />
                    <SPLIT distance="1400" swimtime="00:20:11.52" />
                    <SPLIT distance="1450" swimtime="00:20:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="473" reactiontime="+82" swimtime="00:01:00.18" resultid="10537" heatid="13988" lane="1" entrytime="00:00:58.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="357" reactiontime="+75" swimtime="00:02:23.73" resultid="10538" heatid="14051" lane="5" entrytime="00:02:15.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:47.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="327" swimtime="00:05:19.16" resultid="10539" heatid="14112" lane="9" entrytime="00:05:15.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:52.71" />
                    <SPLIT distance="200" swimtime="00:02:33.89" />
                    <SPLIT distance="250" swimtime="00:03:14.43" />
                    <SPLIT distance="300" swimtime="00:03:56.00" />
                    <SPLIT distance="350" swimtime="00:04:38.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzta" gender="F" lastname="Wach" nation="POL" athleteid="10453">
              <RESULTS>
                <RESULT eventid="1062" points="244" reactiontime="+84" swimtime="00:00:37.93" resultid="10454" heatid="13899" lane="7" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="275" reactiontime="+66" swimtime="00:00:41.57" resultid="10455" heatid="13946" lane="6" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="232" reactiontime="+91" swimtime="00:01:24.68" resultid="10456" heatid="13973" lane="6" entrytime="00:01:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="255" reactiontime="+67" swimtime="00:01:31.62" resultid="10457" heatid="14030" lane="1" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="239" reactiontime="+84" swimtime="00:00:47.49" resultid="10458" heatid="14084" lane="3" entrytime="00:00:47.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-08-12" firstname="Konrad" gender="M" lastname="Plutecki" nation="POL" athleteid="10445">
              <RESULTS>
                <RESULT eventid="1079" points="461" reactiontime="+80" swimtime="00:00:27.05" resultid="10446" heatid="13916" lane="0" entrytime="00:00:26.06" entrycourse="LCM" />
                <RESULT eventid="1205" points="358" reactiontime="+72" swimtime="00:00:33.84" resultid="10447" heatid="13956" lane="6" entrytime="00:00:33.33" entrycourse="LCM" />
                <RESULT eventid="1273" points="483" reactiontime="+77" swimtime="00:00:59.75" resultid="10448" heatid="13988" lane="2" entrytime="00:00:58.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="378" reactiontime="+73" swimtime="00:01:20.07" resultid="10449" heatid="14011" lane="3" entrytime="00:01:18.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="378" reactiontime="+78" swimtime="00:02:20.96" resultid="10450" heatid="14051" lane="4" entrytime="00:02:15.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="363" reactiontime="+74" swimtime="00:02:36.80" resultid="10451" heatid="14081" lane="6" entrytime="00:02:35.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="150" swimtime="00:01:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="384" reactiontime="+75" swimtime="00:05:02.71" resultid="10452" heatid="14112" lane="4" entrytime="00:04:59.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:11.09" />
                    <SPLIT distance="150" swimtime="00:01:50.68" />
                    <SPLIT distance="200" swimtime="00:02:29.70" />
                    <SPLIT distance="250" swimtime="00:03:08.66" />
                    <SPLIT distance="300" swimtime="00:03:47.74" />
                    <SPLIT distance="350" swimtime="00:04:26.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-04-02" firstname="Jacek" gender="M" lastname="Tyczyński" nation="POL" athleteid="10543">
              <RESULTS>
                <RESULT eventid="1165" points="373" reactiontime="+90" swimtime="00:20:09.59" resultid="10544" heatid="13943" lane="2" entrytime="00:19:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:50.31" />
                    <SPLIT distance="200" swimtime="00:02:29.94" />
                    <SPLIT distance="250" swimtime="00:03:10.16" />
                    <SPLIT distance="300" swimtime="00:03:50.98" />
                    <SPLIT distance="350" swimtime="00:04:31.35" />
                    <SPLIT distance="400" swimtime="00:05:11.85" />
                    <SPLIT distance="450" swimtime="00:05:52.55" />
                    <SPLIT distance="500" swimtime="00:06:33.39" />
                    <SPLIT distance="550" swimtime="00:07:14.26" />
                    <SPLIT distance="600" swimtime="00:07:54.85" />
                    <SPLIT distance="650" swimtime="00:08:35.84" />
                    <SPLIT distance="700" swimtime="00:09:17.62" />
                    <SPLIT distance="750" swimtime="00:09:58.61" />
                    <SPLIT distance="800" swimtime="00:10:40.01" />
                    <SPLIT distance="850" swimtime="00:11:20.05" />
                    <SPLIT distance="900" swimtime="00:12:00.37" />
                    <SPLIT distance="950" swimtime="00:12:40.87" />
                    <SPLIT distance="1000" swimtime="00:13:22.88" />
                    <SPLIT distance="1050" swimtime="00:14:03.70" />
                    <SPLIT distance="1100" swimtime="00:14:44.92" />
                    <SPLIT distance="1150" swimtime="00:15:26.35" />
                    <SPLIT distance="1200" swimtime="00:16:07.53" />
                    <SPLIT distance="1250" swimtime="00:16:48.05" />
                    <SPLIT distance="1300" swimtime="00:17:28.37" />
                    <SPLIT distance="1350" swimtime="00:18:08.36" />
                    <SPLIT distance="1400" swimtime="00:18:49.21" />
                    <SPLIT distance="1450" swimtime="00:19:29.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="10400">
              <RESULTS>
                <RESULT eventid="1187" points="445" reactiontime="+54" swimtime="00:00:35.42" resultid="10401" heatid="13947" lane="7" entrytime="00:00:37.80" entrycourse="LCM" />
                <RESULT eventid="1457" points="421" reactiontime="+59" swimtime="00:01:17.49" resultid="10402" heatid="14031" lane="8" entrytime="00:01:19.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="324" reactiontime="+87" swimtime="00:06:30.44" resultid="10403" heatid="14057" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:36.51" />
                    <SPLIT distance="150" swimtime="00:02:24.79" />
                    <SPLIT distance="200" swimtime="00:03:12.46" />
                    <SPLIT distance="250" swimtime="00:04:09.50" />
                    <SPLIT distance="300" swimtime="00:05:05.55" />
                    <SPLIT distance="350" swimtime="00:05:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="384" reactiontime="+62" swimtime="00:02:50.59" resultid="10404" heatid="14075" lane="0" entrytime="00:02:58.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:08.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" athleteid="10466">
              <RESULTS>
                <RESULT eventid="1062" points="113" reactiontime="+116" swimtime="00:00:49.05" resultid="10467" heatid="13897" lane="1" entrytime="00:00:47.00" entrycourse="LCM" />
                <RESULT eventid="1096" points="83" reactiontime="+132" swimtime="00:04:48.29" resultid="10468" heatid="13918" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.50" />
                    <SPLIT distance="100" swimtime="00:02:23.71" />
                    <SPLIT distance="150" swimtime="00:03:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="93" reactiontime="+96" swimtime="00:00:59.69" resultid="10469" heatid="13944" lane="2" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="92" reactiontime="+119" swimtime="00:01:55.13" resultid="10470" heatid="13971" lane="7" entrytime="00:01:51.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="115" reactiontime="+129" swimtime="00:02:12.10" resultid="10471" heatid="14001" lane="0" entrytime="00:02:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="74" swimtime="00:02:17.88" resultid="10472" heatid="14028" lane="4" entrytime="00:02:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="114" reactiontime="+128" swimtime="00:01:00.78" resultid="10473" heatid="14083" lane="2" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1721" points="88" reactiontime="+143" swimtime="00:08:54.81" resultid="10474" heatid="14102" lane="2" entrytime="00:09:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                    <SPLIT distance="100" swimtime="00:01:57.35" />
                    <SPLIT distance="150" swimtime="00:03:05.18" />
                    <SPLIT distance="200" swimtime="00:04:14.30" />
                    <SPLIT distance="250" swimtime="00:05:24.07" />
                    <SPLIT distance="300" swimtime="00:06:35.13" />
                    <SPLIT distance="350" swimtime="00:07:47.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-30" firstname="Szymon" gender="M" lastname="Łenyk" nation="POL" athleteid="10438">
              <RESULTS>
                <RESULT eventid="1079" points="194" reactiontime="+114" swimtime="00:00:36.09" resultid="10439" heatid="13903" lane="2" />
                <RESULT comment="(Time: 19:41), Przekroczony regulaminowy limit czasu." eventid="1165" reactiontime="+128" status="OTL" swimtime="00:00:00.00" resultid="10440" heatid="13939" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:39.22" />
                    <SPLIT distance="150" swimtime="00:02:36.33" />
                    <SPLIT distance="200" swimtime="00:03:37.45" />
                    <SPLIT distance="250" swimtime="00:04:37.62" />
                    <SPLIT distance="300" swimtime="00:05:39.75" />
                    <SPLIT distance="350" swimtime="00:06:42.31" />
                    <SPLIT distance="400" swimtime="00:07:44.04" />
                    <SPLIT distance="450" swimtime="00:08:45.77" />
                    <SPLIT distance="500" swimtime="00:09:47.88" />
                    <SPLIT distance="550" swimtime="00:10:50.87" />
                    <SPLIT distance="600" swimtime="00:11:53.91" />
                    <SPLIT distance="650" swimtime="00:12:56.40" />
                    <SPLIT distance="700" swimtime="00:13:59.24" />
                    <SPLIT distance="750" swimtime="00:15:02.19" />
                    <SPLIT distance="800" swimtime="00:16:05.11" />
                    <SPLIT distance="850" swimtime="00:17:08.17" />
                    <SPLIT distance="900" swimtime="00:18:10.68" />
                    <SPLIT distance="950" swimtime="00:19:12.51" />
                    <SPLIT distance="1000" swimtime="00:20:14.89" />
                    <SPLIT distance="1050" swimtime="00:21:17.49" />
                    <SPLIT distance="1100" swimtime="00:22:19.75" />
                    <SPLIT distance="1150" swimtime="00:23:23.56" />
                    <SPLIT distance="1200" swimtime="00:24:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="110" reactiontime="+99" swimtime="00:00:50.12" resultid="10441" heatid="13949" lane="8" />
                <RESULT eventid="1273" points="151" reactiontime="+105" swimtime="00:01:27.94" resultid="10442" heatid="13977" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="10443" heatid="14032" lane="6" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 10:55)" eventid="1681" reactiontime="+94" status="DSQ" swimtime="00:00:49.75" resultid="10444" heatid="14088" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="10405">
              <RESULTS>
                <RESULT eventid="1062" points="129" reactiontime="+118" swimtime="00:00:46.94" resultid="10406" heatid="13897" lane="0" entrytime="00:00:49.00" entrycourse="LCM" />
                <RESULT eventid="1096" points="89" reactiontime="+114" swimtime="00:04:41.87" resultid="10407" heatid="13918" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.29" />
                    <SPLIT distance="100" swimtime="00:02:15.70" />
                    <SPLIT distance="150" swimtime="00:03:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="109" reactiontime="+73" swimtime="00:00:56.51" resultid="10408" heatid="13944" lane="4" entrytime="00:00:57.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="99" reactiontime="+110" swimtime="00:01:52.22" resultid="10409" heatid="13971" lane="0" entrytime="00:02:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:59)" eventid="1423" reactiontime="+70" status="DSQ" swimtime="00:01:01.41" resultid="10410" heatid="14014" lane="4" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1457" points="89" reactiontime="+83" swimtime="00:02:09.79" resultid="10411" heatid="14028" lane="5" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="56" reactiontime="+128" swimtime="00:02:24.92" resultid="10412" heatid="14063" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="91" reactiontime="+87" swimtime="00:04:35.19" resultid="10413" heatid="14073" lane="8" entrytime="00:04:39.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.39" />
                    <SPLIT distance="100" swimtime="00:02:14.17" />
                    <SPLIT distance="150" swimtime="00:03:26.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-10" firstname="Witold" gender="M" lastname="Śmiałek" nation="POL" athleteid="10434">
              <RESULTS>
                <RESULT eventid="1079" points="158" reactiontime="+93" swimtime="00:00:38.62" resultid="10435" heatid="13905" lane="3" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1205" points="118" reactiontime="+85" swimtime="00:00:49.01" resultid="10436" heatid="13949" lane="7" />
                <RESULT eventid="1474" points="85" reactiontime="+114" swimtime="00:01:58.04" resultid="10437" heatid="14032" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzta" gender="F" lastname="Skalska" nation="POL" athleteid="10459">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="10460" heatid="13918" lane="8" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="10461" heatid="13961" lane="9" entrytime="00:03:34.31" entrycourse="LCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="10462" heatid="13973" lane="8" entrytime="00:01:29.74" entrycourse="LCM" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="10463" heatid="14015" lane="2" entrytime="00:00:45.26" entrycourse="LCM" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="10464" heatid="14040" lane="6" entrytime="00:03:17.32" entrycourse="LCM" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="10465" heatid="14103" lane="9" entrytime="00:07:10.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="10526">
              <RESULTS>
                <RESULT eventid="1079" points="361" reactiontime="+81" swimtime="00:00:29.34" resultid="10527" heatid="13911" lane="6" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT eventid="1113" points="218" reactiontime="+90" swimtime="00:03:09.35" resultid="10528" heatid="13926" lane="7" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:02:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="364" reactiontime="+81" swimtime="00:01:05.66" resultid="10529" heatid="13983" lane="8" entrytime="00:01:07.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="256" reactiontime="+89" swimtime="00:00:35.32" resultid="10530" heatid="14020" lane="4" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1508" points="264" swimtime="00:02:38.96" resultid="10531" heatid="14049" lane="9" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="236" reactiontime="+85" swimtime="00:00:42.73" resultid="10532" heatid="14092" lane="2" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1744" points="238" reactiontime="+92" swimtime="00:05:55.03" resultid="10533" heatid="14110" lane="0" entrytime="00:05:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:19.07" />
                    <SPLIT distance="150" swimtime="00:02:05.22" />
                    <SPLIT distance="200" swimtime="00:02:52.95" />
                    <SPLIT distance="250" swimtime="00:03:40.52" />
                    <SPLIT distance="300" swimtime="00:04:27.55" />
                    <SPLIT distance="350" swimtime="00:05:14.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-03-22" firstname="Sandra" gender="F" lastname="Wolska" nation="POL" athleteid="10481">
              <RESULTS>
                <RESULT eventid="1062" points="352" reactiontime="+89" swimtime="00:00:33.58" resultid="10482" heatid="13901" lane="1" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1096" points="286" reactiontime="+92" swimtime="00:03:11.40" resultid="10483" heatid="13920" lane="2" entrytime="00:03:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:01:34.46" />
                    <SPLIT distance="150" swimtime="00:02:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="337" reactiontime="+90" swimtime="00:03:19.77" resultid="10484" heatid="13961" lane="3" entrytime="00:03:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:02:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="166" swimtime="00:03:41.28" resultid="10485" heatid="13991" lane="9" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:41.78" />
                    <SPLIT distance="150" swimtime="00:02:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="267" reactiontime="+91" swimtime="00:02:55.37" resultid="10486" heatid="14039" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:20.79" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="272" reactiontime="+94" swimtime="00:06:53.80" resultid="10487" heatid="14058" lane="2" entrytime="00:06:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:38.81" />
                    <SPLIT distance="150" swimtime="00:02:32.98" />
                    <SPLIT distance="200" swimtime="00:03:25.98" />
                    <SPLIT distance="250" swimtime="00:04:20.57" />
                    <SPLIT distance="300" swimtime="00:05:16.19" />
                    <SPLIT distance="350" swimtime="00:06:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="216" reactiontime="+80" swimtime="00:03:26.72" resultid="10488" heatid="14072" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.69" />
                    <SPLIT distance="100" swimtime="00:01:41.85" />
                    <SPLIT distance="150" swimtime="00:02:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="346" reactiontime="+87" swimtime="00:00:41.96" resultid="10489" heatid="14087" lane="8" entrytime="00:00:38.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Wisła 4" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="476" reactiontime="+59" swimtime="00:01:59.59" resultid="10548" heatid="13999" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                    <SPLIT distance="150" swimtime="00:01:33.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10475" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="10425" number="2" />
                    <RELAYPOSITION athleteid="10534" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="10490" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="10549" heatid="14056" lane="4" entrytime="00:01:44.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10425" number="1" />
                    <RELAYPOSITION athleteid="10475" number="2" />
                    <RELAYPOSITION athleteid="10534" number="3" />
                    <RELAYPOSITION athleteid="10490" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Wisła 5" number="5">
              <RESULTS>
                <RESULT eventid="1381" points="210" reactiontime="+92" swimtime="00:02:37.05" resultid="10550" heatid="13998" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.24" />
                    <SPLIT distance="100" swimtime="00:01:30.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10438" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="10388" number="2" />
                    <RELAYPOSITION athleteid="10393" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="10526" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="251" reactiontime="+87" swimtime="00:02:14.46" resultid="10551" heatid="14055" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="150" swimtime="00:01:44.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10438" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="10388" number="2" />
                    <RELAYPOSITION athleteid="10393" number="3" />
                    <RELAYPOSITION athleteid="10526" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Wisła 6" number="6">
              <RESULTS>
                <RESULT eventid="1381" points="65" swimtime="00:03:51.65" resultid="10552" heatid="13997" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.77" />
                    <SPLIT distance="100" swimtime="00:02:01.04" />
                    <SPLIT distance="150" swimtime="00:03:27.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10504" number="1" />
                    <RELAYPOSITION athleteid="10510" number="2" />
                    <RELAYPOSITION athleteid="10540" number="3" reactiontime="+96" />
                    <RELAYPOSITION athleteid="10434" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Wisła 7" number="7">
              <RESULTS>
                <RESULT eventid="1358" points="254" reactiontime="+65" swimtime="00:02:47.60" resultid="10553" heatid="13996" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:36.01" />
                    <SPLIT distance="150" swimtime="00:02:10.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10517" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="10414" number="2" />
                    <RELAYPOSITION athleteid="10400" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="10453" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="263" reactiontime="+78" swimtime="00:02:30.67" resultid="10554" heatid="14054" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:08.89" />
                    <SPLIT distance="150" swimtime="00:01:56.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10517" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="10453" number="2" />
                    <RELAYPOSITION athleteid="10414" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="10400" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Wisła 1" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="83" reactiontime="+113" swimtime="00:03:13.84" resultid="10545" heatid="13932" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                    <SPLIT distance="100" swimtime="00:01:41.09" />
                    <SPLIT distance="150" swimtime="00:02:34.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10405" number="1" reactiontime="+113" />
                    <RELAYPOSITION athleteid="10504" number="2" />
                    <RELAYPOSITION athleteid="10466" number="3" reactiontime="+108" />
                    <RELAYPOSITION athleteid="10434" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Wisła 2" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="330" reactiontime="+78" swimtime="00:02:02.70" resultid="10546" heatid="13932" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:00:58.40" />
                    <SPLIT distance="150" swimtime="00:01:36.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10517" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="10534" number="2" />
                    <RELAYPOSITION athleteid="10453" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="10490" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" name="Wisła 3" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="342" reactiontime="+83" swimtime="00:02:01.22" resultid="10547" heatid="13933" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="150" swimtime="00:01:34.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10481" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="10445" number="2" />
                    <RELAYPOSITION athleteid="10496" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10543" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="Wisła 8" number="8">
              <RESULTS>
                <RESULT eventid="1698" points="362" swimtime="00:02:11.04" resultid="10555" heatid="14101" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="150" swimtime="00:01:45.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10517" number="1" />
                    <RELAYPOSITION athleteid="10490" number="2" />
                    <RELAYPOSITION athleteid="10400" number="3" />
                    <RELAYPOSITION athleteid="10475" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Wisła 9" number="9">
              <RESULTS>
                <RESULT eventid="1698" points="141" reactiontime="+81" swimtime="00:02:59.39" resultid="10556" heatid="14100" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                    <SPLIT distance="100" swimtime="00:01:33.86" />
                    <SPLIT distance="150" swimtime="00:02:09.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10414" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="10388" number="2" />
                    <RELAYPOSITION athleteid="10393" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="10466" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Wisła 10" number="10">
              <RESULTS>
                <RESULT eventid="1698" points="138" reactiontime="+69" swimtime="00:03:00.77" resultid="10557" heatid="14099" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:01:39.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10453" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="10405" number="2" />
                    <RELAYPOSITION athleteid="10534" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="10504" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11707" name="MASTERS Zdzieszowice">
          <CONTACT city="Zdzieszowice" email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" state="OPO" zip="47-330" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-13" firstname="Magda" gender="F" lastname="Gorostiza" nation="POL" athleteid="11743">
              <RESULTS>
                <RESULT eventid="1222" points="257" reactiontime="+97" swimtime="00:03:38.74" resultid="11744" heatid="13962" lane="0" entrytime="00:03:15.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:43.33" />
                    <SPLIT distance="150" swimtime="00:02:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="263" reactiontime="+97" swimtime="00:01:21.23" resultid="11745" heatid="13972" lane="3" entrytime="00:01:30.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="288" reactiontime="+93" swimtime="00:01:37.35" resultid="11746" heatid="14002" lane="4" entrytime="00:01:35.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="237" reactiontime="+92" swimtime="00:03:02.49" resultid="11747" heatid="14041" lane="7" entrytime="00:02:52.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:27.07" />
                    <SPLIT distance="150" swimtime="00:02:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="325" reactiontime="+91" swimtime="00:00:42.84" resultid="11748" heatid="14086" lane="3" entrytime="00:00:40.01" />
                <RESULT eventid="1721" points="210" reactiontime="+99" swimtime="00:06:40.60" resultid="11749" heatid="14104" lane="7" entrytime="00:05:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                    <SPLIT distance="150" swimtime="00:02:20.01" />
                    <SPLIT distance="200" swimtime="00:03:11.13" />
                    <SPLIT distance="250" swimtime="00:04:03.16" />
                    <SPLIT distance="300" swimtime="00:04:56.20" />
                    <SPLIT distance="350" swimtime="00:05:48.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="11708">
              <RESULTS>
                <RESULT eventid="1113" points="470" reactiontime="+77" swimtime="00:02:26.54" resultid="11709" heatid="13931" lane="3" entrytime="00:02:19.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="349" swimtime="00:20:36.30" resultid="11710" heatid="13939" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:16.32" />
                    <SPLIT distance="150" swimtime="00:01:57.46" />
                    <SPLIT distance="200" swimtime="00:02:38.93" />
                    <SPLIT distance="250" swimtime="00:03:20.21" />
                    <SPLIT distance="300" swimtime="00:04:01.33" />
                    <SPLIT distance="350" swimtime="00:04:42.15" />
                    <SPLIT distance="400" swimtime="00:05:23.62" />
                    <SPLIT distance="450" swimtime="00:06:04.96" />
                    <SPLIT distance="500" swimtime="00:06:45.98" />
                    <SPLIT distance="550" swimtime="00:07:26.66" />
                    <SPLIT distance="600" swimtime="00:08:08.04" />
                    <SPLIT distance="650" swimtime="00:08:49.35" />
                    <SPLIT distance="700" swimtime="00:09:30.65" />
                    <SPLIT distance="750" swimtime="00:10:11.90" />
                    <SPLIT distance="800" swimtime="00:10:53.59" />
                    <SPLIT distance="850" swimtime="00:11:35.41" />
                    <SPLIT distance="900" swimtime="00:12:17.34" />
                    <SPLIT distance="950" swimtime="00:12:59.10" />
                    <SPLIT distance="1000" swimtime="00:13:40.95" />
                    <SPLIT distance="1050" swimtime="00:14:22.38" />
                    <SPLIT distance="1100" swimtime="00:15:04.12" />
                    <SPLIT distance="1150" swimtime="00:15:46.11" />
                    <SPLIT distance="1200" swimtime="00:16:27.86" />
                    <SPLIT distance="1250" swimtime="00:17:09.73" />
                    <SPLIT distance="1300" swimtime="00:17:51.55" />
                    <SPLIT distance="1350" swimtime="00:18:32.95" />
                    <SPLIT distance="1400" swimtime="00:19:14.69" />
                    <SPLIT distance="1450" swimtime="00:19:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="11711" heatid="13977" lane="6" />
                <RESULT eventid="1341" points="402" reactiontime="+77" swimtime="00:02:31.05" resultid="11712" heatid="13995" lane="5" entrytime="00:02:29.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="459" reactiontime="+82" swimtime="00:02:12.20" resultid="11713" heatid="14045" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="440" reactiontime="+75" swimtime="00:05:20.39" resultid="11714" heatid="14062" lane="5" entrytime="00:05:08.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:56.44" />
                    <SPLIT distance="200" swimtime="00:02:39.18" />
                    <SPLIT distance="250" swimtime="00:03:23.52" />
                    <SPLIT distance="300" swimtime="00:04:08.90" />
                    <SPLIT distance="350" swimtime="00:04:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="481" reactiontime="+78" swimtime="00:01:03.55" resultid="11715" heatid="14071" lane="7" entrytime="00:01:01.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="434" reactiontime="+80" swimtime="00:04:50.65" resultid="11716" heatid="14113" lane="5" entrytime="00:04:45.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                    <SPLIT distance="200" swimtime="00:02:25.60" />
                    <SPLIT distance="250" swimtime="00:03:02.48" />
                    <SPLIT distance="300" swimtime="00:03:39.57" />
                    <SPLIT distance="350" swimtime="00:04:16.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="11717">
              <RESULTS>
                <RESULT eventid="1079" points="405" reactiontime="+80" swimtime="00:00:28.25" resultid="11718" heatid="13910" lane="4" entrytime="00:00:30.01" />
                <RESULT eventid="1113" points="345" swimtime="00:02:42.48" resultid="11719" heatid="13930" lane="9" entrytime="00:02:36.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="11720" heatid="13984" lane="3" entrytime="00:01:03.21" />
                <RESULT eventid="1341" points="329" reactiontime="+94" swimtime="00:02:41.52" resultid="11721" heatid="13995" lane="6" entrytime="00:02:36.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="335" swimtime="00:01:23.35" resultid="11722" heatid="14010" lane="6" entrytime="00:01:20.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="308" swimtime="00:06:00.69" resultid="11723" heatid="14062" lane="9" entrytime="00:05:41.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                    <SPLIT distance="200" swimtime="00:02:57.11" />
                    <SPLIT distance="250" swimtime="00:03:50.55" />
                    <SPLIT distance="300" swimtime="00:04:43.02" />
                    <SPLIT distance="350" swimtime="00:05:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="346" reactiontime="+89" swimtime="00:01:10.96" resultid="11724" heatid="14070" lane="3" entrytime="00:01:08.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11725" heatid="14112" lane="2" entrytime="00:05:05.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Grzegorz" gender="M" lastname="Sierka" nation="POL" athleteid="11740">
              <RESULTS>
                <RESULT eventid="1440" points="495" reactiontime="+83" swimtime="00:00:28.34" resultid="11741" heatid="14027" lane="1" entrytime="00:00:27.65" />
                <RESULT eventid="1474" points="436" reactiontime="+67" swimtime="00:01:08.45" resultid="11742" heatid="14038" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-18" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="11726">
              <RESULTS>
                <RESULT eventid="1096" points="298" reactiontime="+102" swimtime="00:03:08.74" resultid="11727" heatid="13920" lane="0" entrytime="00:03:10.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="283" reactiontime="+77" swimtime="00:00:41.17" resultid="11728" heatid="13947" lane="1" entrytime="00:00:37.86" />
                <RESULT eventid="1256" points="292" reactiontime="+93" swimtime="00:01:18.43" resultid="11729" heatid="13974" lane="7" entrytime="00:01:17.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="267" reactiontime="+99" swimtime="00:00:37.93" resultid="11730" heatid="14016" lane="2" entrytime="00:00:36.61" />
                <RESULT eventid="1457" points="286" reactiontime="+77" swimtime="00:01:28.19" resultid="11731" heatid="14030" lane="7" entrytime="00:01:28.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="285" reactiontime="+83" swimtime="00:03:08.31" resultid="11732" heatid="14074" lane="2" entrytime="00:03:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:32.55" />
                    <SPLIT distance="150" swimtime="00:02:21.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-23" firstname="Katarzyna" gender="F" lastname="Gniot" nation="POL" athleteid="11733">
              <RESULTS>
                <RESULT eventid="1062" points="223" reactiontime="+107" swimtime="00:00:39.13" resultid="11734" heatid="13897" lane="3" entrytime="00:00:43.22" />
                <RESULT eventid="1187" points="118" reactiontime="+72" swimtime="00:00:55.09" resultid="11735" heatid="13946" lane="8" entrytime="00:00:42.34" />
                <RESULT eventid="1256" points="178" reactiontime="+117" swimtime="00:01:32.46" resultid="11736" heatid="13972" lane="0" entrytime="00:01:35.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="170" reactiontime="+95" swimtime="00:01:56.08" resultid="11737" heatid="14002" lane="8" entrytime="00:01:45.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="104" reactiontime="+93" swimtime="00:02:03.20" resultid="11738" heatid="14029" lane="7" entrytime="00:01:50.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="11739" heatid="14085" lane="0" entrytime="00:00:45.55" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="249" reactiontime="+103" swimtime="00:02:14.84" resultid="11750" heatid="13933" lane="6" entrytime="00:02:15.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11726" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="11733" number="2" />
                    <RELAYPOSITION athleteid="11717" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="11708" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="280" reactiontime="+76" swimtime="00:02:22.68" resultid="11751" heatid="14100" lane="3" entrytime="00:02:20.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11726" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="11743" number="2" />
                    <RELAYPOSITION athleteid="11717" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="11708" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10952" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos" phone="604184311" street="Rafał" />
          <ATHLETES>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="10975">
              <RESULTS>
                <RESULT eventid="1079" points="429" reactiontime="+83" swimtime="00:00:27.71" resultid="10976" heatid="13916" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="359" reactiontime="+100" swimtime="00:01:05.97" resultid="10977" heatid="13985" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="334" reactiontime="+103" swimtime="00:00:32.32" resultid="10978" heatid="14022" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1681" points="360" swimtime="00:00:37.13" resultid="10979" heatid="14096" lane="9" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="10980">
              <RESULTS>
                <RESULT eventid="1113" points="240" reactiontime="+90" swimtime="00:03:03.20" resultid="10981" heatid="13930" lane="8" entrytime="00:02:34.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="150" swimtime="00:02:18.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="10983" heatid="13983" lane="9" entrytime="00:01:07.89" />
                <RESULT eventid="1474" points="257" reactiontime="+85" swimtime="00:01:21.67" resultid="10984" heatid="14035" lane="3" entrytime="00:01:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="10985" heatid="14068" lane="4" entrytime="00:01:22.01" />
                <RESULT eventid="1744" points="270" swimtime="00:05:40.11" resultid="10986" heatid="14110" lane="9" entrytime="00:05:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                    <SPLIT distance="200" swimtime="00:02:46.47" />
                    <SPLIT distance="250" swimtime="00:03:30.82" />
                    <SPLIT distance="300" swimtime="00:04:16.25" />
                    <SPLIT distance="350" swimtime="00:04:59.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="10959">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:32)" eventid="1079" reactiontime="+68" status="DSQ" swimtime="00:00:27.11" resultid="10960" heatid="13912" lane="4" entrytime="00:00:28.04" />
                <RESULT eventid="1113" points="409" reactiontime="+91" swimtime="00:02:33.50" resultid="10961" heatid="13929" lane="4" entrytime="00:02:38.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="456" reactiontime="+82" swimtime="00:01:00.93" resultid="10962" heatid="13985" lane="5" entrytime="00:01:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="448" reactiontime="+91" swimtime="00:00:29.30" resultid="10963" heatid="14025" lane="1" entrytime="00:00:30.32" />
                <RESULT eventid="1508" points="389" swimtime="00:02:19.67" resultid="10964" heatid="14051" lane="9" entrytime="00:02:22.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                    <SPLIT distance="150" swimtime="00:01:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="398" reactiontime="+105" swimtime="00:00:35.89" resultid="10965" heatid="14094" lane="1" entrytime="00:00:37.69" />
                <RESULT eventid="1744" points="351" reactiontime="+90" swimtime="00:05:11.81" resultid="10966" heatid="14111" lane="5" entrytime="00:05:18.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:46.77" />
                    <SPLIT distance="200" swimtime="00:02:25.98" />
                    <SPLIT distance="250" swimtime="00:03:07.10" />
                    <SPLIT distance="300" swimtime="00:03:48.76" />
                    <SPLIT distance="350" swimtime="00:04:31.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="10967">
              <RESULTS>
                <RESULT eventid="1079" points="279" reactiontime="+103" swimtime="00:00:31.99" resultid="10968" heatid="13907" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1113" points="169" reactiontime="+114" swimtime="00:03:25.83" resultid="10969" heatid="13925" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:41.41" />
                    <SPLIT distance="150" swimtime="00:02:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="10970" heatid="13953" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="10971" heatid="13967" lane="9" entrytime="00:03:20.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="10972" heatid="14008" lane="1" entrytime="00:01:31.00" />
                <RESULT eventid="1647" points="158" reactiontime="+88" swimtime="00:03:26.99" resultid="10973" heatid="14079" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="1681" points="249" reactiontime="+92" swimtime="00:00:41.97" resultid="10974" heatid="14092" lane="7" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="10953">
              <RESULTS>
                <RESULT eventid="1113" points="361" reactiontime="+81" swimtime="00:02:39.99" resultid="10954" heatid="13929" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="388" reactiontime="+84" swimtime="00:02:54.08" resultid="10955" heatid="13969" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="415" reactiontime="+79" swimtime="00:01:17.61" resultid="10956" heatid="14012" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="394" swimtime="00:00:30.58" resultid="10957" heatid="14025" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1681" points="460" reactiontime="+77" swimtime="00:00:34.22" resultid="10958" heatid="14097" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="10987">
              <RESULTS>
                <RESULT eventid="1113" points="412" reactiontime="+88" swimtime="00:02:33.10" resultid="10988" heatid="13927" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="467" reactiontime="+60" swimtime="00:00:30.98" resultid="10989" heatid="13955" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1341" points="259" reactiontime="+92" swimtime="00:02:54.74" resultid="10990" heatid="13994" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="10991" heatid="14011" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1474" points="433" reactiontime="+61" swimtime="00:01:08.61" resultid="10992" heatid="14037" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="10993" heatid="14047" lane="3" entrytime="00:02:50.00" />
                <RESULT eventid="1681" points="462" reactiontime="+83" swimtime="00:00:34.17" resultid="10994" heatid="14095" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="423" reactiontime="+63" swimtime="00:02:04.42" resultid="10995" heatid="13999" lane="9" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:06.70" />
                    <SPLIT distance="150" swimtime="00:01:36.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10987" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="10953" number="2" />
                    <RELAYPOSITION athleteid="10959" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="10975" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="438" reactiontime="+85" swimtime="00:01:51.65" resultid="10996" heatid="14056" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="100" swimtime="00:00:56.22" />
                    <SPLIT distance="150" swimtime="00:01:23.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10967" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="10987" number="2" />
                    <RELAYPOSITION athleteid="10959" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="10975" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASTKRAS" nation="POL" region="LU" clubid="9745" name="Masterskrasnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="9750">
              <RESULTS>
                <RESULT eventid="1079" points="284" reactiontime="+63" swimtime="00:00:31.78" resultid="9751" heatid="13910" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1165" points="150" reactiontime="+97" swimtime="00:27:17.51" resultid="9752" heatid="13940" lane="2" entrytime="00:25:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:31.18" />
                    <SPLIT distance="200" swimtime="00:03:26.36" />
                    <SPLIT distance="250" swimtime="00:04:21.91" />
                    <SPLIT distance="300" swimtime="00:05:18.52" />
                    <SPLIT distance="350" swimtime="00:06:14.04" />
                    <SPLIT distance="400" swimtime="00:07:11.48" />
                    <SPLIT distance="450" swimtime="00:08:05.81" />
                    <SPLIT distance="500" swimtime="00:09:01.89" />
                    <SPLIT distance="550" swimtime="00:09:58.31" />
                    <SPLIT distance="600" swimtime="00:10:55.25" />
                    <SPLIT distance="650" swimtime="00:11:51.11" />
                    <SPLIT distance="700" swimtime="00:12:47.98" />
                    <SPLIT distance="750" swimtime="00:13:43.02" />
                    <SPLIT distance="800" swimtime="00:14:39.67" />
                    <SPLIT distance="850" swimtime="00:15:34.87" />
                    <SPLIT distance="900" swimtime="00:16:31.64" />
                    <SPLIT distance="950" swimtime="00:17:26.24" />
                    <SPLIT distance="1000" swimtime="00:18:23.98" />
                    <SPLIT distance="1050" swimtime="00:19:18.03" />
                    <SPLIT distance="1100" swimtime="00:20:14.33" />
                    <SPLIT distance="1150" swimtime="00:21:10.22" />
                    <SPLIT distance="1200" swimtime="00:22:04.08" />
                    <SPLIT distance="1250" swimtime="00:22:58.44" />
                    <SPLIT distance="1300" swimtime="00:23:53.69" />
                    <SPLIT distance="1350" swimtime="00:24:47.78" />
                    <SPLIT distance="1400" swimtime="00:25:41.22" />
                    <SPLIT distance="1450" swimtime="00:26:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="227" reactiontime="+60" swimtime="00:00:39.39" resultid="9753" heatid="13953" lane="3" entrytime="00:00:38.20" />
                <RESULT eventid="1341" points="82" reactiontime="+90" swimtime="00:04:16.22" resultid="9754" heatid="13992" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                    <SPLIT distance="100" swimtime="00:02:01.93" />
                    <SPLIT distance="150" swimtime="00:03:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="9755" heatid="14034" lane="5" entrytime="00:01:29.30" />
                <RESULT eventid="1578" points="146" reactiontime="+95" swimtime="00:07:43.02" resultid="9756" heatid="14060" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.25" />
                    <SPLIT distance="100" swimtime="00:01:56.29" />
                    <SPLIT distance="150" swimtime="00:02:55.02" />
                    <SPLIT distance="200" swimtime="00:03:53.37" />
                    <SPLIT distance="250" swimtime="00:05:00.19" />
                    <SPLIT distance="300" swimtime="00:06:05.62" />
                    <SPLIT distance="350" swimtime="00:06:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="132" reactiontime="+81" swimtime="00:01:37.67" resultid="9757" heatid="14068" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="9758" heatid="14079" lane="1" entrytime="00:03:18.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-02-09" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="9746">
              <RESULTS>
                <RESULT eventid="1273" points="189" swimtime="00:01:21.70" resultid="9747" heatid="13981" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="164" reactiontime="+94" swimtime="00:03:06.34" resultid="9748" heatid="14047" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                    <SPLIT distance="150" swimtime="00:02:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="168" reactiontime="+98" swimtime="00:06:38.58" resultid="9749" heatid="14114" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:02:15.35" />
                    <SPLIT distance="200" swimtime="00:03:07.33" />
                    <SPLIT distance="250" swimtime="00:03:59.18" />
                    <SPLIT distance="300" swimtime="00:04:52.62" />
                    <SPLIT distance="350" swimtime="00:05:46.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="9759">
              <RESULTS>
                <RESULT eventid="1239" points="308" reactiontime="+92" swimtime="00:03:07.87" resultid="9760" heatid="13967" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                    <SPLIT distance="150" swimtime="00:02:19.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="319" reactiontime="+94" swimtime="00:01:24.71" resultid="9761" heatid="14009" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="301" reactiontime="+101" swimtime="00:00:39.39" resultid="9762" heatid="14094" lane="0" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="9763">
              <RESULTS>
                <RESULT eventid="1205" points="96" reactiontime="+82" swimtime="00:00:52.48" resultid="9764" heatid="13950" lane="2" entrytime="00:00:56.29" />
                <RESULT eventid="1239" points="91" reactiontime="+96" swimtime="00:04:41.48" resultid="9765" heatid="13964" lane="5" entrytime="00:04:15.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.43" />
                    <SPLIT distance="100" swimtime="00:02:13.42" />
                    <SPLIT distance="150" swimtime="00:03:29.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="94" reactiontime="+97" swimtime="00:02:07.06" resultid="9766" heatid="14006" lane="7" entrytime="00:01:59.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="96" reactiontime="+99" swimtime="00:00:48.84" resultid="9767" heatid="14019" lane="7" entrytime="00:00:55.27" />
                <RESULT eventid="1613" points="57" reactiontime="+102" swimtime="00:02:09.13" resultid="9768" heatid="14066" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" nation="POL" region="PDK" clubid="9433" name="Mkp Bobry Dębica">
          <CONTACT name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1991-10-29" firstname="Marcin" gender="M" lastname="Potoczny" nation="POL" athleteid="9615">
              <RESULTS>
                <RESULT eventid="1079" points="145" reactiontime="+84" swimtime="00:00:39.78" resultid="9616" heatid="13905" lane="0" entrytime="00:00:43.29" />
                <RESULT eventid="1205" points="104" reactiontime="+76" swimtime="00:00:50.98" resultid="9617" heatid="13951" lane="6" entrytime="00:00:49.71" />
                <RESULT eventid="1273" points="135" reactiontime="+90" swimtime="00:01:31.43" resultid="9618" heatid="13978" lane="6" entrytime="00:01:44.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="109" reactiontime="+80" swimtime="00:03:32.98" resultid="12461" heatid="14044" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:37.72" />
                    <SPLIT distance="150" swimtime="00:02:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="118" swimtime="00:07:28.25" resultid="12462" heatid="14107" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:01:38.81" />
                    <SPLIT distance="150" swimtime="00:02:36.66" />
                    <SPLIT distance="200" swimtime="00:03:34.58" />
                    <SPLIT distance="250" swimtime="00:04:34.24" />
                    <SPLIT distance="300" swimtime="00:05:33.44" />
                    <SPLIT distance="350" swimtime="00:06:33.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-11" firstname="Przemysław" gender="M" lastname="Jurek" nation="POL" athleteid="9605">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1079" points="563" reactiontime="+82" swimtime="00:00:25.32" resultid="9606" heatid="13917" lane="3" entrytime="00:00:24.80" />
                <RESULT eventid="1113" points="449" reactiontime="+86" swimtime="00:02:28.82" resultid="9607" heatid="13931" lane="8" entrytime="00:02:25.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:07.73" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="567" reactiontime="+86" swimtime="00:00:56.65" resultid="9608" heatid="13989" lane="5" entrytime="00:00:55.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="494" reactiontime="+88" swimtime="00:00:28.37" resultid="9609" heatid="14027" lane="0" entrytime="00:00:27.78" />
                <RESULT eventid="1613" points="510" reactiontime="+88" swimtime="00:01:02.33" resultid="9610" heatid="14071" lane="2" entrytime="00:01:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-25" firstname="Adam" gender="M" lastname="Wytrwał" nation="POL" athleteid="9625">
              <RESULTS>
                <RESULT eventid="1165" points="274" reactiontime="+104" swimtime="00:22:20.18" resultid="9626" heatid="13942" lane="1" entrytime="00:21:25.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                    <SPLIT distance="200" swimtime="00:02:46.00" />
                    <SPLIT distance="250" swimtime="00:03:30.74" />
                    <SPLIT distance="300" swimtime="00:04:14.94" />
                    <SPLIT distance="350" swimtime="00:05:00.40" />
                    <SPLIT distance="400" swimtime="00:05:45.70" />
                    <SPLIT distance="450" swimtime="00:06:31.13" />
                    <SPLIT distance="500" swimtime="00:07:16.16" />
                    <SPLIT distance="550" swimtime="00:08:01.58" />
                    <SPLIT distance="600" swimtime="00:08:47.07" />
                    <SPLIT distance="650" swimtime="00:09:32.46" />
                    <SPLIT distance="700" swimtime="00:10:17.21" />
                    <SPLIT distance="750" swimtime="00:11:02.84" />
                    <SPLIT distance="800" swimtime="00:11:48.03" />
                    <SPLIT distance="850" swimtime="00:12:33.36" />
                    <SPLIT distance="900" swimtime="00:13:18.83" />
                    <SPLIT distance="950" swimtime="00:14:04.17" />
                    <SPLIT distance="1000" swimtime="00:14:50.94" />
                    <SPLIT distance="1050" swimtime="00:15:36.64" />
                    <SPLIT distance="1100" swimtime="00:16:21.43" />
                    <SPLIT distance="1150" swimtime="00:18:36.88" />
                    <SPLIT distance="1200" swimtime="00:17:51.56" />
                    <SPLIT distance="1250" swimtime="00:20:07.57" />
                    <SPLIT distance="1300" swimtime="00:19:22.02" />
                    <SPLIT distance="1400" swimtime="00:20:52.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" athleteid="9611">
              <RESULTS>
                <RESULT eventid="1165" points="355" reactiontime="+104" swimtime="00:20:29.72" resultid="9612" heatid="13942" lane="2" entrytime="00:21:19.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:15.83" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                    <SPLIT distance="200" swimtime="00:02:36.97" />
                    <SPLIT distance="250" swimtime="00:03:17.51" />
                    <SPLIT distance="300" swimtime="00:03:58.67" />
                    <SPLIT distance="350" swimtime="00:04:39.36" />
                    <SPLIT distance="400" swimtime="00:05:20.49" />
                    <SPLIT distance="450" swimtime="00:06:01.06" />
                    <SPLIT distance="500" swimtime="00:06:42.48" />
                    <SPLIT distance="550" swimtime="00:07:22.50" />
                    <SPLIT distance="600" swimtime="00:08:03.29" />
                    <SPLIT distance="650" swimtime="00:08:44.01" />
                    <SPLIT distance="700" swimtime="00:09:25.49" />
                    <SPLIT distance="750" swimtime="00:10:06.63" />
                    <SPLIT distance="800" swimtime="00:10:47.92" />
                    <SPLIT distance="850" swimtime="00:11:29.25" />
                    <SPLIT distance="900" swimtime="00:12:10.93" />
                    <SPLIT distance="950" swimtime="00:12:51.77" />
                    <SPLIT distance="1000" swimtime="00:13:33.47" />
                    <SPLIT distance="1050" swimtime="00:14:15.19" />
                    <SPLIT distance="1100" swimtime="00:14:57.19" />
                    <SPLIT distance="1150" swimtime="00:15:39.47" />
                    <SPLIT distance="1200" swimtime="00:16:21.01" />
                    <SPLIT distance="1250" swimtime="00:17:02.42" />
                    <SPLIT distance="1300" swimtime="00:17:44.39" />
                    <SPLIT distance="1350" swimtime="00:18:25.85" />
                    <SPLIT distance="1400" swimtime="00:19:08.35" />
                    <SPLIT distance="1450" swimtime="00:19:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="309" reactiontime="+96" swimtime="00:02:44.91" resultid="9613" heatid="13992" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="285" reactiontime="+98" swimtime="00:06:10.21" resultid="9614" heatid="14059" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:02:08.80" />
                    <SPLIT distance="200" swimtime="00:03:00.33" />
                    <SPLIT distance="250" swimtime="00:03:53.85" />
                    <SPLIT distance="300" swimtime="00:04:48.86" />
                    <SPLIT distance="350" swimtime="00:05:30.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-14" firstname="Jan" gender="M" lastname="Wałaszek" nation="POL" athleteid="9627">
              <RESULTS>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="9628" heatid="13940" lane="0" entrytime="00:26:41.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-23" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="500308600142" athleteid="9629">
              <RESULTS>
                <RESULT eventid="1187" points="395" reactiontime="+75" swimtime="00:00:36.88" resultid="9630" heatid="13948" lane="7" entrytime="00:00:34.90" />
                <RESULT eventid="1457" points="392" reactiontime="+76" swimtime="00:01:19.36" resultid="9631" heatid="14031" lane="6" entrytime="00:01:14.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="403" reactiontime="+73" swimtime="00:02:47.91" resultid="9632" heatid="14075" lane="6" entrytime="00:02:41.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:05.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-08" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="9619">
              <RESULTS>
                <RESULT eventid="1113" points="127" reactiontime="+118" swimtime="00:03:46.35" resultid="9620" heatid="13923" lane="3" entrytime="00:03:46.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:48.44" />
                    <SPLIT distance="150" swimtime="00:02:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="176" reactiontime="+122" swimtime="00:25:53.04" resultid="9621" heatid="13940" lane="7" entrytime="00:25:12.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                    <SPLIT distance="150" swimtime="00:02:14.95" />
                    <SPLIT distance="200" swimtime="00:03:07.36" />
                    <SPLIT distance="250" swimtime="00:03:59.31" />
                    <SPLIT distance="300" swimtime="00:04:52.56" />
                    <SPLIT distance="350" swimtime="00:05:46.15" />
                    <SPLIT distance="400" swimtime="00:06:38.53" />
                    <SPLIT distance="450" swimtime="00:07:31.05" />
                    <SPLIT distance="500" swimtime="00:08:25.14" />
                    <SPLIT distance="550" swimtime="00:09:18.77" />
                    <SPLIT distance="600" swimtime="00:10:13.20" />
                    <SPLIT distance="650" swimtime="00:11:07.43" />
                    <SPLIT distance="700" swimtime="00:12:02.04" />
                    <SPLIT distance="750" swimtime="00:12:55.77" />
                    <SPLIT distance="800" swimtime="00:13:50.18" />
                    <SPLIT distance="850" swimtime="00:14:43.81" />
                    <SPLIT distance="900" swimtime="00:15:38.16" />
                    <SPLIT distance="950" swimtime="00:16:31.84" />
                    <SPLIT distance="1000" swimtime="00:17:26.28" />
                    <SPLIT distance="1050" swimtime="00:18:21.06" />
                    <SPLIT distance="1100" swimtime="00:19:15.10" />
                    <SPLIT distance="1150" swimtime="00:20:08.81" />
                    <SPLIT distance="1200" swimtime="00:21:03.29" />
                    <SPLIT distance="1250" swimtime="00:21:57.29" />
                    <SPLIT distance="1300" swimtime="00:22:52.16" />
                    <SPLIT distance="1350" swimtime="00:23:46.54" />
                    <SPLIT distance="1400" swimtime="00:24:40.96" />
                    <SPLIT distance="1450" swimtime="00:25:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="207" reactiontime="+116" swimtime="00:01:19.22" resultid="9622" heatid="13979" lane="4" entrytime="00:01:21.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="193" reactiontime="+118" swimtime="00:02:56.36" resultid="9623" heatid="14046" lane="3" entrytime="00:03:03.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:21.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="196" swimtime="00:06:18.43" resultid="9624" heatid="14108" lane="6" entrytime="00:06:30.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:11.77" />
                    <SPLIT distance="200" swimtime="00:03:01.13" />
                    <SPLIT distance="250" swimtime="00:03:51.35" />
                    <SPLIT distance="300" swimtime="00:04:41.22" />
                    <SPLIT distance="350" swimtime="00:05:31.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="ZAC" clubid="9360" name="MKP Szczecin">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" internet="numer kodowy 001/16" name="Kowalczyk Piotr" phone="509758055" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="11565">
              <RESULTS>
                <RESULT eventid="1222" points="93" swimtime="00:05:06.13" resultid="11566" heatid="13960" lane="9" entrytime="00:04:57.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.94" />
                    <SPLIT distance="100" swimtime="00:02:30.56" />
                    <SPLIT distance="150" swimtime="00:03:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="78" swimtime="00:02:30.26" resultid="11567" heatid="14001" lane="9" entrytime="00:02:20.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="78" swimtime="00:01:08.85" resultid="11568" heatid="14083" lane="8" entrytime="00:01:09.73" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="11553">
              <RESULTS>
                <RESULT eventid="1079" points="309" reactiontime="+99" swimtime="00:00:30.91" resultid="11554" heatid="13909" lane="3" entrytime="00:00:31.20" />
                <RESULT eventid="1165" points="254" reactiontime="+119" swimtime="00:22:54.79" resultid="11555" heatid="13941" lane="1" entrytime="00:22:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:08.28" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:05:12.83" />
                    <SPLIT distance="200" swimtime="00:02:53.59" />
                    <SPLIT distance="250" swimtime="00:06:44.50" />
                    <SPLIT distance="300" swimtime="00:04:26.42" />
                    <SPLIT distance="350" swimtime="00:08:15.54" />
                    <SPLIT distance="400" swimtime="00:05:59.07" />
                    <SPLIT distance="450" swimtime="00:09:48.33" />
                    <SPLIT distance="500" swimtime="00:07:30.26" />
                    <SPLIT distance="550" swimtime="00:11:21.83" />
                    <SPLIT distance="600" swimtime="00:09:02.01" />
                    <SPLIT distance="650" swimtime="00:12:54.24" />
                    <SPLIT distance="700" swimtime="00:10:35.36" />
                    <SPLIT distance="750" swimtime="00:14:27.26" />
                    <SPLIT distance="800" swimtime="00:12:08.86" />
                    <SPLIT distance="850" swimtime="00:16:00.59" />
                    <SPLIT distance="900" swimtime="00:13:40.26" />
                    <SPLIT distance="950" swimtime="00:17:33.65" />
                    <SPLIT distance="1000" swimtime="00:15:13.70" />
                    <SPLIT distance="1050" swimtime="00:19:07.74" />
                    <SPLIT distance="1100" swimtime="00:16:46.65" />
                    <SPLIT distance="1150" swimtime="00:20:40.43" />
                    <SPLIT distance="1200" swimtime="00:18:20.95" />
                    <SPLIT distance="1250" swimtime="00:22:12.13" />
                    <SPLIT distance="1300" swimtime="00:19:54.00" />
                    <SPLIT distance="1400" swimtime="00:21:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="296" reactiontime="+104" swimtime="00:01:10.32" resultid="11556" heatid="13982" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="251" swimtime="00:02:41.50" resultid="11557" heatid="14048" lane="9" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:02:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11558" heatid="14110" lane="1" entrytime="00:05:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="11547">
              <RESULTS>
                <RESULT eventid="1165" points="331" swimtime="00:20:58.47" resultid="11548" heatid="13943" lane="9" entrytime="00:20:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                    <SPLIT distance="200" swimtime="00:02:33.86" />
                    <SPLIT distance="250" swimtime="00:04:39.06" />
                    <SPLIT distance="300" swimtime="00:03:57.00" />
                    <SPLIT distance="350" swimtime="00:06:03.72" />
                    <SPLIT distance="400" swimtime="00:05:21.33" />
                    <SPLIT distance="450" swimtime="00:07:29.31" />
                    <SPLIT distance="500" swimtime="00:06:46.24" />
                    <SPLIT distance="550" swimtime="00:08:54.38" />
                    <SPLIT distance="600" swimtime="00:08:11.59" />
                    <SPLIT distance="650" swimtime="00:10:19.70" />
                    <SPLIT distance="700" swimtime="00:09:37.11" />
                    <SPLIT distance="750" swimtime="00:11:45.90" />
                    <SPLIT distance="800" swimtime="00:11:02.14" />
                    <SPLIT distance="850" swimtime="00:13:10.96" />
                    <SPLIT distance="900" swimtime="00:12:28.79" />
                    <SPLIT distance="950" swimtime="00:14:37.37" />
                    <SPLIT distance="1000" swimtime="00:13:53.90" />
                    <SPLIT distance="1050" swimtime="00:16:04.44" />
                    <SPLIT distance="1100" swimtime="00:15:20.92" />
                    <SPLIT distance="1150" swimtime="00:17:30.71" />
                    <SPLIT distance="1200" swimtime="00:16:47.58" />
                    <SPLIT distance="1250" swimtime="00:18:56.29" />
                    <SPLIT distance="1300" swimtime="00:18:14.03" />
                    <SPLIT distance="1400" swimtime="00:19:39.28" />
                    <SPLIT distance="1450" swimtime="00:20:21.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="391" reactiontime="+84" swimtime="00:01:04.13" resultid="11549" heatid="13985" lane="6" entrytime="00:01:02.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="350" reactiontime="+87" swimtime="00:02:24.60" resultid="11550" heatid="14051" lane="7" entrytime="00:02:19.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11551" heatid="14080" lane="3" entrytime="00:02:48.00" />
                <RESULT eventid="1744" points="372" reactiontime="+91" swimtime="00:05:05.73" resultid="11552" heatid="14112" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:51.76" />
                    <SPLIT distance="200" swimtime="00:02:31.40" />
                    <SPLIT distance="250" swimtime="00:03:10.63" />
                    <SPLIT distance="300" swimtime="00:03:50.64" />
                    <SPLIT distance="350" swimtime="00:04:29.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="11559">
              <RESULTS>
                <RESULT eventid="1113" points="358" reactiontime="+98" swimtime="00:02:40.41" resultid="11560" heatid="13930" lane="2" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:02:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="425" reactiontime="+109" swimtime="00:19:18.43" resultid="11561" heatid="13943" lane="0" entrytime="00:19:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                    <SPLIT distance="200" swimtime="00:02:23.55" />
                    <SPLIT distance="250" swimtime="00:03:00.75" />
                    <SPLIT distance="300" swimtime="00:03:38.30" />
                    <SPLIT distance="350" swimtime="00:04:16.16" />
                    <SPLIT distance="400" swimtime="00:04:54.28" />
                    <SPLIT distance="450" swimtime="00:05:32.21" />
                    <SPLIT distance="500" swimtime="00:06:10.55" />
                    <SPLIT distance="550" swimtime="00:06:49.27" />
                    <SPLIT distance="600" swimtime="00:07:28.16" />
                    <SPLIT distance="650" swimtime="00:08:07.04" />
                    <SPLIT distance="700" swimtime="00:08:46.64" />
                    <SPLIT distance="750" swimtime="00:09:26.57" />
                    <SPLIT distance="800" swimtime="00:10:06.81" />
                    <SPLIT distance="850" swimtime="00:10:46.29" />
                    <SPLIT distance="900" swimtime="00:11:25.83" />
                    <SPLIT distance="950" swimtime="00:12:05.12" />
                    <SPLIT distance="1000" swimtime="00:12:44.60" />
                    <SPLIT distance="1050" swimtime="00:13:23.89" />
                    <SPLIT distance="1100" swimtime="00:14:03.45" />
                    <SPLIT distance="1150" swimtime="00:14:42.18" />
                    <SPLIT distance="1200" swimtime="00:15:21.52" />
                    <SPLIT distance="1250" swimtime="00:16:00.97" />
                    <SPLIT distance="1300" swimtime="00:16:40.31" />
                    <SPLIT distance="1350" swimtime="00:17:20.18" />
                    <SPLIT distance="1400" swimtime="00:18:00.02" />
                    <SPLIT distance="1450" swimtime="00:18:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="330" reactiontime="+100" swimtime="00:02:41.33" resultid="11562" heatid="13995" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:02:00.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="416" reactiontime="+102" swimtime="00:05:26.39" resultid="11563" heatid="14062" lane="2" entrytime="00:05:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:13.33" />
                    <SPLIT distance="150" swimtime="00:01:56.52" />
                    <SPLIT distance="200" swimtime="00:02:37.83" />
                    <SPLIT distance="250" swimtime="00:03:26.05" />
                    <SPLIT distance="300" swimtime="00:04:15.22" />
                    <SPLIT distance="350" swimtime="00:04:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="444" reactiontime="+96" swimtime="00:04:48.34" resultid="11564" heatid="14114" lane="0" entrytime="00:04:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:42.85" />
                    <SPLIT distance="200" swimtime="00:02:19.73" />
                    <SPLIT distance="250" swimtime="00:02:56.34" />
                    <SPLIT distance="300" swimtime="00:03:33.72" />
                    <SPLIT distance="350" swimtime="00:04:11.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-31" firstname="Konrad" gender="M" lastname="Tekiel" nation="POL" athleteid="11576">
              <RESULTS>
                <RESULT eventid="1508" points="139" reactiontime="+110" swimtime="00:03:16.79" resultid="11577" heatid="14047" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:33.05" />
                    <SPLIT distance="150" swimtime="00:02:24.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="139" reactiontime="+102" swimtime="00:07:04.07" resultid="11578" heatid="14108" lane="1" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="100" swimtime="00:01:43.37" />
                    <SPLIT distance="150" swimtime="00:02:38.76" />
                    <SPLIT distance="200" swimtime="00:03:33.80" />
                    <SPLIT distance="250" swimtime="00:04:29.05" />
                    <SPLIT distance="300" swimtime="00:05:22.75" />
                    <SPLIT distance="350" swimtime="00:06:15.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="11571">
              <RESULTS>
                <RESULT eventid="1113" points="160" reactiontime="+103" swimtime="00:03:29.80" resultid="11572" heatid="13924" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="11573" heatid="13965" lane="4" entrytime="00:03:40.00" />
                <RESULT eventid="1406" points="201" reactiontime="+90" swimtime="00:01:38.84" resultid="11574" heatid="14007" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="240" reactiontime="+88" swimtime="00:00:42.48" resultid="11575" heatid="14090" lane="7" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="11569">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="11570" heatid="13906" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-09" firstname="Piotr" gender="M" lastname="Nowicki" nation="POL" athleteid="11579">
              <RESULTS>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="11580" heatid="14047" lane="8" entrytime="00:02:55.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11581" heatid="14108" lane="0" entrytime="00:06:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="9DDZ" nation="POL" region="DOL" clubid="12070" name="Mks Dziewiątka Dzierżoniów">
          <CONTACT name="Piotr Kuszka" phone="604226649" />
          <ATHLETES>
            <ATHLETE birthdate="1989-01-17" firstname="Piotr" gender="M" lastname="Gołębiowski" nation="POL" athleteid="12075">
              <RESULTS>
                <RESULT eventid="1205" points="379" reactiontime="+72" swimtime="00:00:33.20" resultid="12076" heatid="13958" lane="0" entrytime="00:00:30.50" />
                <RESULT eventid="1273" points="447" reactiontime="+94" swimtime="00:01:01.33" resultid="12077" heatid="13986" lane="8" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="487" reactiontime="+89" swimtime="00:00:28.50" resultid="12078" heatid="14027" lane="8" entrytime="00:00:27.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-03" firstname="Krzysztof" gender="M" lastname="Pawlaczek" nation="POL" athleteid="12071">
              <RESULTS>
                <RESULT eventid="1239" points="363" reactiontime="+83" swimtime="00:02:57.93" resultid="12072" heatid="13969" lane="0" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="380" reactiontime="+82" swimtime="00:01:19.94" resultid="12073" heatid="14011" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="409" reactiontime="+84" swimtime="00:00:30.20" resultid="12074" heatid="14024" lane="5" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-14" firstname="Piotr" gender="M" lastname="Kuszka" nation="POL" athleteid="12083">
              <RESULTS>
                <RESULT eventid="1239" points="215" reactiontime="+95" swimtime="00:03:32.00" resultid="12084" heatid="13966" lane="3" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:42.29" />
                    <SPLIT distance="150" swimtime="00:02:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="210" swimtime="00:01:18.81" resultid="12085" heatid="13980" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="215" reactiontime="+96" swimtime="00:01:36.66" resultid="12086" heatid="14007" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="189" reactiontime="+94" swimtime="00:00:39.04" resultid="12087" heatid="14019" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-09-02" firstname="Małgorzata" gender="F" lastname="Morańda" nation="POL" athleteid="12079">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="12080" heatid="13944" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="12081" heatid="13971" lane="2" entrytime="00:01:50.00" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="12082" heatid="14001" lane="8" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01111" nation="POL" region="SLA" clubid="11094" name="Mks Mos Katowice">
          <CONTACT city="KATOWICE" email="zanuli@wp.pl" name="ORPEL ANNA" phone="502348487" state="ŚLĄSK" street="PADEREWSKIEGO 46A" zip="40-282" />
          <ATHLETES>
            <ATHLETE birthdate="1994-12-04" firstname="Paweł" gender="M" lastname="Ulfik" nation="POL" license="101111200016" athleteid="11095">
              <RESULTS>
                <RESULT eventid="1205" points="414" reactiontime="+68" swimtime="00:00:32.23" resultid="11096" heatid="13954" lane="1" entrytime="00:00:36.54" />
                <RESULT eventid="1239" points="348" reactiontime="+87" swimtime="00:03:00.42" resultid="11097" heatid="13969" lane="1" entrytime="00:02:52.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:13.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="368" reactiontime="+79" swimtime="00:01:20.80" resultid="11098" heatid="14011" lane="1" entrytime="00:01:19.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="380" reactiontime="+69" swimtime="00:01:11.65" resultid="11099" heatid="14037" lane="2" entrytime="00:01:10.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="382" reactiontime="+61" swimtime="00:02:34.15" resultid="11100" heatid="14081" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="392" swimtime="00:00:36.08" resultid="11101" heatid="14097" lane="9" entrytime="00:00:34.81" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01011" nation="POL" region="SLA" clubid="12179" name="MKS Park Wodny Tarnowskie Góry">
          <CONTACT city="Tarnowskie Góry" name="Macner Dagmara" phone="509691784" state="SLA" street="Obwodnica 8" zip="42-600" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-15" firstname="Mateusz" gender="M" lastname="Kotkowski" nameprefix="MK" nation="POL" license="1" athleteid="12180">
              <RESULTS>
                <RESULT eventid="1079" points="492" reactiontime="+73" swimtime="00:00:26.48" resultid="12181" heatid="13916" lane="8" entrytime="00:00:26.03" />
                <RESULT eventid="1113" points="438" reactiontime="+75" swimtime="00:02:30.06" resultid="12182" heatid="13929" lane="8" entrytime="00:02:40.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="511" reactiontime="+77" swimtime="00:00:58.64" resultid="12183" heatid="13988" lane="7" entrytime="00:00:58.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="485" reactiontime="+82" swimtime="00:00:28.54" resultid="12184" heatid="14026" lane="2" entrytime="00:00:28.27" />
                <RESULT eventid="1508" points="459" swimtime="00:02:12.19" resultid="12185" heatid="14052" lane="9" entrytime="00:02:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:04.11" />
                    <SPLIT distance="150" swimtime="00:01:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="444" swimtime="00:04:48.36" resultid="12186" heatid="14114" lane="9" entrytime="00:04:41.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="150" swimtime="00:01:40.15" />
                    <SPLIT distance="200" swimtime="00:02:17.18" />
                    <SPLIT distance="250" swimtime="00:02:54.89" />
                    <SPLIT distance="300" swimtime="00:03:33.82" />
                    <SPLIT distance="350" swimtime="00:04:12.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-30" firstname="Kajetan" gender="M" lastname="Smoliński" nameprefix="SK" nation="POL" license="2" athleteid="12187">
              <RESULTS>
                <RESULT eventid="1079" points="500" reactiontime="+78" swimtime="00:00:26.33" resultid="12188" heatid="13916" lane="3" entrytime="00:00:25.97" />
                <RESULT eventid="1273" points="483" reactiontime="+74" swimtime="00:00:59.78" resultid="12189" heatid="13989" lane="8" entrytime="00:00:57.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="12190" heatid="14026" lane="7" entrytime="00:00:28.33" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00811" nation="POL" region="SLA" clubid="9916" name="MKS Pałac Młodzieży Katowice">
          <CONTACT city="Katowice" email="r.puchalski@duosport.pl" name="Puchalski Robert" state="ŚLĄSK" street="Mikołowska 26" zip="40-066" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-01" firstname="Błażej" gender="M" lastname="Kornaga" nation="POL" athleteid="9917">
              <RESULTS>
                <RESULT eventid="1079" points="371" swimtime="00:00:29.09" resultid="9918" heatid="13904" lane="9" />
                <RESULT eventid="1273" points="365" reactiontime="+84" swimtime="00:01:05.60" resultid="9919" heatid="13984" lane="8" entrytime="00:01:04.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="298" reactiontime="+79" swimtime="00:02:32.62" resultid="9920" heatid="14050" lane="1" entrytime="00:02:27.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="274" reactiontime="+92" swimtime="00:05:38.46" resultid="9921" heatid="14111" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:00.55" />
                    <SPLIT distance="200" swimtime="00:02:44.46" />
                    <SPLIT distance="250" swimtime="00:03:29.44" />
                    <SPLIT distance="300" swimtime="00:04:14.22" />
                    <SPLIT distance="350" swimtime="00:04:58.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-08-16" firstname="Jacek" gender="M" lastname="Syska" nation="POL" athleteid="9922">
              <RESULTS>
                <RESULT eventid="1079" points="236" reactiontime="+91" swimtime="00:00:33.79" resultid="9923" heatid="13903" lane="5" />
                <RESULT eventid="1440" points="237" reactiontime="+87" swimtime="00:00:36.24" resultid="9924" heatid="14020" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" region="DOL" clubid="10090" name="Mks Swim Academy Termy Jakuba Oława" shortname="Mks Swim Academy Termy Jakuba ">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOL" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE birthdate="1991-07-06" firstname="Agnieszka" gender="F" lastname="Burdelak" nation="POL" license="5045016000019" athleteid="10091">
              <RESULTS>
                <RESULT eventid="1062" points="512" reactiontime="+70" swimtime="00:00:29.66" resultid="10092" heatid="13902" lane="6" entrytime="00:00:28.90" />
                <RESULT eventid="1222" points="444" reactiontime="+72" swimtime="00:03:02.21" resultid="10093" heatid="13962" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="456" swimtime="00:01:23.56" resultid="10094" heatid="14004" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="419" reactiontime="+78" swimtime="00:02:30.98" resultid="10095" heatid="14043" lane="2" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="482" swimtime="00:00:37.59" resultid="10096" heatid="14087" lane="6" entrytime="00:00:37.40" />
                <RESULT eventid="1721" points="374" reactiontime="+70" swimtime="00:05:30.65" resultid="10097" heatid="14105" lane="8" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:17.91" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                    <SPLIT distance="200" swimtime="00:02:41.87" />
                    <SPLIT distance="250" swimtime="00:03:23.31" />
                    <SPLIT distance="300" swimtime="00:04:06.39" />
                    <SPLIT distance="350" swimtime="00:04:49.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9571" name="MOSiR KSZO Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="9591">
              <RESULTS>
                <RESULT eventid="1079" points="248" swimtime="00:00:33.26" resultid="9592" heatid="13908" lane="9" entrytime="00:00:33.30" />
                <RESULT eventid="1113" points="151" reactiontime="+90" swimtime="00:03:33.66" resultid="9593" heatid="13923" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:47.01" />
                    <SPLIT distance="150" swimtime="00:02:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="138" reactiontime="+91" swimtime="00:04:05.38" resultid="9594" heatid="13965" lane="8" entrytime="00:03:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:56.70" />
                    <SPLIT distance="150" swimtime="00:03:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="186" reactiontime="+101" swimtime="00:01:22.12" resultid="9595" heatid="13980" lane="3" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="219" swimtime="00:00:37.19" resultid="9596" heatid="14020" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1508" points="139" reactiontime="+103" swimtime="00:03:16.54" resultid="9597" heatid="14046" lane="7" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:26.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="110" reactiontime="+105" swimtime="00:01:43.96" resultid="9598" heatid="14067" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="216" reactiontime="+101" swimtime="00:00:44.00" resultid="9599" heatid="14091" lane="7" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="PDK" clubid="11118" name="MOTYL  MOSiR Stalowa Wola">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Andzrej Chmielewski" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="11590">
              <RESULTS>
                <RESULT eventid="1079" points="449" swimtime="00:00:27.30" resultid="11591" heatid="13915" lane="9" entrytime="00:00:26.92" />
                <RESULT eventid="1113" points="395" reactiontime="+88" swimtime="00:02:35.34" resultid="11592" heatid="13930" lane="7" entrytime="00:02:33.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="475" reactiontime="+75" swimtime="00:00:30.80" resultid="11593" heatid="13958" lane="8" entrytime="00:00:30.31" />
                <RESULT eventid="1273" points="454" reactiontime="+88" swimtime="00:01:01.00" resultid="11594" heatid="13986" lane="6" entrytime="00:01:00.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="382" swimtime="00:00:30.89" resultid="11595" heatid="14023" lane="6" entrytime="00:00:32.10" />
                <RESULT eventid="1474" points="427" reactiontime="+78" swimtime="00:01:08.94" resultid="11596" heatid="14038" lane="1" entrytime="00:01:07.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="377" reactiontime="+79" swimtime="00:02:34.91" resultid="11597" heatid="14082" lane="8" entrytime="00:02:32.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="330" reactiontime="+82" swimtime="00:00:38.23" resultid="11598" heatid="14096" lane="4" entrytime="00:00:34.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="11599">
              <RESULTS>
                <RESULT eventid="1079" points="420" reactiontime="+80" swimtime="00:00:27.91" resultid="11600" heatid="13912" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1205" points="291" swimtime="00:00:36.24" resultid="11601" heatid="13955" lane="2" entrytime="00:00:35.20" />
                <RESULT eventid="1341" points="178" reactiontime="+103" swimtime="00:03:17.90" resultid="11602" heatid="13994" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:31.40" />
                    <SPLIT distance="150" swimtime="00:02:25.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="366" reactiontime="+90" swimtime="00:00:31.35" resultid="11603" heatid="14024" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="11604" heatid="14069" lane="5" entrytime="00:01:16.80" />
                <RESULT eventid="1647" points="237" reactiontime="+78" swimtime="00:03:00.74" resultid="11605" heatid="14080" lane="9" entrytime="00:03:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:13.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-07" firstname="Paweł" gender="M" lastname="Ciurko" nation="POL" athleteid="11615">
              <RESULTS>
                <RESULT eventid="1079" points="220" swimtime="00:00:34.60" resultid="11616" heatid="13907" lane="9" entrytime="00:00:35.30" />
                <RESULT eventid="1113" points="287" reactiontime="+80" swimtime="00:02:52.68" resultid="11617" heatid="13926" lane="2" entrytime="00:02:59.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="150" swimtime="00:02:13.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="300" reactiontime="+86" swimtime="00:03:09.54" resultid="11618" heatid="13967" lane="1" entrytime="00:03:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:32.70" />
                    <SPLIT distance="150" swimtime="00:02:21.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="169" reactiontime="+86" swimtime="00:03:21.54" resultid="11619" heatid="13993" lane="4" entrytime="00:03:19.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:36.47" />
                    <SPLIT distance="150" swimtime="00:02:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="11620" heatid="14009" lane="5" entrytime="00:01:24.17" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="11621" heatid="14060" lane="0" entrytime="00:07:32.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="11582">
              <RESULTS>
                <RESULT eventid="1062" points="299" reactiontime="+94" swimtime="00:00:35.48" resultid="11583" heatid="13899" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1096" points="280" swimtime="00:03:12.61" resultid="11584" heatid="13920" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:02:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="263" reactiontime="+81" swimtime="00:03:36.94" resultid="11585" heatid="13960" lane="4" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:43.28" />
                    <SPLIT distance="150" swimtime="00:02:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="248" reactiontime="+94" swimtime="00:01:42.39" resultid="11586" heatid="14002" lane="7" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="261" reactiontime="+97" swimtime="00:06:59.89" resultid="11587" heatid="14058" lane="0" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:04:24.88" />
                    <SPLIT distance="200" swimtime="00:03:28.94" />
                    <SPLIT distance="250" swimtime="00:06:12.19" />
                    <SPLIT distance="300" swimtime="00:05:22.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="205" reactiontime="+97" swimtime="00:01:34.23" resultid="11588" heatid="14064" lane="0" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="259" swimtime="00:00:46.19" resultid="11589" heatid="14085" lane="9" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="11606">
              <RESULTS>
                <RESULT eventid="1079" points="296" reactiontime="+89" swimtime="00:00:31.37" resultid="11607" heatid="13909" lane="1" entrytime="00:00:31.53" />
                <RESULT eventid="1113" points="263" reactiontime="+89" swimtime="00:02:57.76" resultid="11608" heatid="13926" lane="3" entrytime="00:02:55.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                    <SPLIT distance="150" swimtime="00:02:17.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="269" reactiontime="+76" swimtime="00:00:37.21" resultid="11609" heatid="13953" lane="6" entrytime="00:00:38.50" />
                <RESULT eventid="1273" points="290" reactiontime="+81" swimtime="00:01:10.82" resultid="11610" heatid="13982" lane="6" entrytime="00:01:09.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="256" reactiontime="+81" swimtime="00:01:21.78" resultid="11611" heatid="14035" lane="5" entrytime="00:01:19.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="250" reactiontime="+89" swimtime="00:06:26.81" resultid="11612" heatid="14061" lane="8" entrytime="00:06:24.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:28.49" />
                    <SPLIT distance="150" swimtime="00:02:16.81" />
                    <SPLIT distance="200" swimtime="00:03:05.47" />
                    <SPLIT distance="250" swimtime="00:04:02.36" />
                    <SPLIT distance="300" swimtime="00:04:59.53" />
                    <SPLIT distance="350" swimtime="00:05:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="235" reactiontime="+83" swimtime="00:03:01.34" resultid="11613" heatid="14080" lane="0" entrytime="00:02:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                    <SPLIT distance="100" swimtime="00:01:28.75" />
                    <SPLIT distance="150" swimtime="00:02:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11614" heatid="14110" lane="8" entrytime="00:05:52.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="11622">
              <RESULTS>
                <RESULT eventid="1079" points="463" reactiontime="+77" swimtime="00:00:27.01" resultid="11623" heatid="13909" lane="0" entrytime="00:00:31.99" />
                <RESULT eventid="1113" points="495" reactiontime="+77" swimtime="00:02:24.02" resultid="11624" heatid="13931" lane="1" entrytime="00:02:22.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="395" reactiontime="+72" swimtime="00:00:32.76" resultid="11625" heatid="13956" lane="1" entrytime="00:00:33.99" />
                <RESULT eventid="1273" points="516" reactiontime="+77" swimtime="00:00:58.46" resultid="11626" heatid="13989" lane="0" entrytime="00:00:57.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="462" reactiontime="+76" swimtime="00:01:14.91" resultid="11627" heatid="14013" lane="7" entrytime="00:01:12.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="496" reactiontime="+77" swimtime="00:00:28.33" resultid="11628" heatid="14027" lane="7" entrytime="00:00:27.39" />
                <RESULT eventid="1613" points="543" reactiontime="+76" swimtime="00:01:01.05" resultid="11629" heatid="14071" lane="5" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="494" swimtime="00:00:33.41" resultid="11630" heatid="14097" lane="6" entrytime="00:00:33.49" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="419" reactiontime="+84" swimtime="00:02:04.83" resultid="11631" heatid="13999" lane="0" entrytime="00:02:05.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:37.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11590" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="11615" number="2" />
                    <RELAYPOSITION athleteid="11622" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="11599" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MSWIM" nation="POL" clubid="11043" name="MSWIM Szczecin">
          <CONTACT email="m@mswim.pl" name="Kaczanowski Miłosz" phone="888181234" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-22" firstname="Miłosz" gender="M" lastname="Kaczanowski" nation="POL" athleteid="11055">
              <RESULTS>
                <RESULT eventid="1079" points="429" reactiontime="+77" swimtime="00:00:27.72" resultid="11056" heatid="13914" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1273" points="474" reactiontime="+73" swimtime="00:01:00.14" resultid="11057" heatid="13987" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="487" reactiontime="+75" swimtime="00:00:28.50" resultid="11058" heatid="14026" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="1613" points="462" reactiontime="+81" swimtime="00:01:04.42" resultid="11059" heatid="14070" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="404" reactiontime="+75" swimtime="00:00:35.71" resultid="11060" heatid="14095" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="11051">
              <RESULTS>
                <RESULT eventid="1187" points="253" reactiontime="+88" swimtime="00:00:42.74" resultid="11052" heatid="13946" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1457" points="249" reactiontime="+90" swimtime="00:01:32.26" resultid="11053" heatid="14030" lane="0" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="244" reactiontime="+83" swimtime="00:03:18.43" resultid="11054" heatid="14074" lane="8" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="100" swimtime="00:01:34.76" />
                    <SPLIT distance="150" swimtime="00:02:26.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="11044">
              <RESULTS>
                <RESULT eventid="1205" points="248" reactiontime="+74" swimtime="00:00:38.22" resultid="11045" heatid="13954" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1239" points="223" reactiontime="+108" swimtime="00:03:29.25" resultid="11046" heatid="13967" lane="0" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:38.82" />
                    <SPLIT distance="150" swimtime="00:02:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="226" reactiontime="+79" swimtime="00:01:25.15" resultid="11047" heatid="14035" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="11048" heatid="14048" lane="5" entrytime="00:02:40.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11049" heatid="14079" lane="5" entrytime="00:03:07.00" />
                <RESULT eventid="1681" points="255" reactiontime="+92" swimtime="00:00:41.61" resultid="11050" heatid="14092" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NABAIJI" nation="POL" clubid="12161" name="Nabaiji Team Decathlon">
          <CONTACT city="Toruń" email="filip.wojciechowski@decathlon.com" name="Filip Wojciechowski" phone="503414875" state="KP" street="ul. Żółkiewskiego 15" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="12175">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="12176" heatid="13900" lane="7" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="12177" heatid="13973" lane="5" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="12178" heatid="14042" lane="9" entrytime="00:02:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-04" firstname="Filip" gender="M" lastname="Wojciechowski" nation="POL" athleteid="12169">
              <RESULTS>
                <RESULT eventid="1079" points="517" reactiontime="+76" swimtime="00:00:26.05" resultid="12170" heatid="13917" lane="0" entrytime="00:00:25.73" entrycourse="LCM" />
                <RESULT eventid="1273" points="560" reactiontime="+74" swimtime="00:00:56.88" resultid="12171" heatid="13989" lane="3" entrytime="00:00:55.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="514" swimtime="00:00:27.99" resultid="12172" heatid="14026" lane="6" entrytime="00:00:28.05" entrycourse="LCM" />
                <RESULT eventid="1508" points="496" reactiontime="+76" swimtime="00:02:08.81" resultid="12173" heatid="14053" lane="3" entrytime="00:02:04.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="150" swimtime="00:01:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="491" reactiontime="+76" swimtime="00:04:38.90" resultid="12174" heatid="14114" lane="5" entrytime="00:04:25.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:04.94" />
                    <SPLIT distance="150" swimtime="00:01:40.40" />
                    <SPLIT distance="200" swimtime="00:02:16.62" />
                    <SPLIT distance="250" swimtime="00:02:52.60" />
                    <SPLIT distance="300" swimtime="00:03:29.28" />
                    <SPLIT distance="350" swimtime="00:04:04.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="12165">
              <RESULTS>
                <RESULT eventid="1079" points="458" reactiontime="+79" swimtime="00:00:27.11" resultid="12166" heatid="13913" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1205" points="418" reactiontime="+78" swimtime="00:00:32.15" resultid="12167" heatid="13957" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1681" points="534" reactiontime="+77" swimtime="00:00:32.55" resultid="12168" heatid="14097" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="10735" name="Nereus Zilina">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1959-11-14" firstname="Rastislav" gender="M" lastname="Pavlik" nation="SVK" athleteid="10736">
              <RESULTS>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="10737" heatid="14038" lane="8" entrytime="00:01:09.70" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10738" heatid="14097" lane="7" entrytime="00:00:33.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORS OPOLE" nation="POL" region="OPO" clubid="10877" name="ORS Opole">
          <CONTACT name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="10883">
              <RESULTS>
                <RESULT eventid="1096" points="415" reactiontime="+86" swimtime="00:02:49.02" resultid="10884" heatid="13921" lane="7" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:02:11.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="357" reactiontime="+86" swimtime="00:11:26.59" resultid="10885" heatid="13937" lane="2" entrytime="00:11:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:02:07.49" />
                    <SPLIT distance="200" swimtime="00:02:51.34" />
                    <SPLIT distance="250" swimtime="00:03:34.66" />
                    <SPLIT distance="300" swimtime="00:04:17.64" />
                    <SPLIT distance="350" swimtime="00:05:00.18" />
                    <SPLIT distance="400" swimtime="00:05:44.31" />
                    <SPLIT distance="450" swimtime="00:06:27.82" />
                    <SPLIT distance="500" swimtime="00:07:11.75" />
                    <SPLIT distance="550" swimtime="00:07:55.14" />
                    <SPLIT distance="600" swimtime="00:08:39.31" />
                    <SPLIT distance="650" swimtime="00:09:23.07" />
                    <SPLIT distance="700" swimtime="00:10:06.59" />
                    <SPLIT distance="750" swimtime="00:10:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="392" reactiontime="+82" swimtime="00:06:06.59" resultid="10886" heatid="14058" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                    <SPLIT distance="150" swimtime="00:02:17.33" />
                    <SPLIT distance="200" swimtime="00:03:04.87" />
                    <SPLIT distance="250" swimtime="00:03:56.93" />
                    <SPLIT distance="300" swimtime="00:04:48.42" />
                    <SPLIT distance="350" swimtime="00:05:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="387" reactiontime="+97" swimtime="00:01:16.30" resultid="10887" heatid="14065" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="375" reactiontime="+94" swimtime="00:05:30.33" resultid="10888" heatid="14105" lane="2" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                    <SPLIT distance="200" swimtime="00:02:43.76" />
                    <SPLIT distance="250" swimtime="00:03:26.81" />
                    <SPLIT distance="300" swimtime="00:04:10.45" />
                    <SPLIT distance="350" swimtime="00:04:52.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Wojciech" gender="M" lastname="Stanek" nation="POL" athleteid="10878">
              <RESULTS>
                <RESULT eventid="1113" points="317" reactiontime="+85" swimtime="00:02:47.02" resultid="10879" heatid="13927" lane="4" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="10880" heatid="13966" lane="4" entrytime="00:03:21.80" />
                <RESULT eventid="1508" points="309" reactiontime="+87" swimtime="00:02:30.82" resultid="10881" heatid="14050" lane="0" entrytime="00:02:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:52.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="314" reactiontime="+77" swimtime="00:05:23.71" resultid="10882" heatid="14111" lane="7" entrytime="00:05:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:01:58.32" />
                    <SPLIT distance="200" swimtime="00:02:39.81" />
                    <SPLIT distance="250" swimtime="00:03:21.46" />
                    <SPLIT distance="300" swimtime="00:04:03.33" />
                    <SPLIT distance="350" swimtime="00:04:44.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KPMTV" nation="SVK" clubid="9911" name="OZ Komunita plavania - Turcianski vlci" shortname="OZ Komunita plavania - Turcian">
          <CONTACT city="Martin" email="brani.hakel@turcianskivlci.sk" internet="turcianskivlci.sk" name="Branislav Hakel" phone="+421915437184" street="Cajkovského štvrt 8/10" zip="03601" />
          <ATHLETES>
            <ATHLETE birthdate="1971-10-14" firstname="Andrea" gender="F" lastname="Liptaiova" nation="SVK" license="SVK17930" athleteid="9912">
              <RESULTS>
                <RESULT eventid="1062" points="366" reactiontime="+87" swimtime="00:00:33.16" resultid="9913" heatid="13900" lane="3" entrytime="00:00:32.80" />
                <RESULT eventid="1388" points="277" reactiontime="+94" swimtime="00:01:38.60" resultid="9914" heatid="14004" lane="0" entrytime="00:01:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 10:54)" eventid="1664" reactiontime="+69" status="DSQ" swimtime="00:00:43.33" resultid="9915" heatid="14087" lane="4" entrytime="00:00:36.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="12093" name="Pregel">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="12100">
              <RESULTS>
                <RESULT eventid="1062" points="639" reactiontime="+83" swimtime="00:00:27.54" resultid="12101" heatid="13902" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1147" points="500" reactiontime="+89" swimtime="00:10:13.79" resultid="12102" heatid="13937" lane="5" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:52.21" />
                    <SPLIT distance="200" swimtime="00:02:31.11" />
                    <SPLIT distance="250" swimtime="00:03:10.27" />
                    <SPLIT distance="300" swimtime="00:03:49.20" />
                    <SPLIT distance="350" swimtime="00:04:27.39" />
                    <SPLIT distance="400" swimtime="00:05:05.73" />
                    <SPLIT distance="450" swimtime="00:05:44.46" />
                    <SPLIT distance="500" swimtime="00:06:23.19" />
                    <SPLIT distance="550" swimtime="00:07:02.15" />
                    <SPLIT distance="600" swimtime="00:07:40.55" />
                    <SPLIT distance="650" swimtime="00:08:19.11" />
                    <SPLIT distance="700" swimtime="00:08:57.69" />
                    <SPLIT distance="750" swimtime="00:09:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="636" reactiontime="+83" swimtime="00:01:00.54" resultid="12103" heatid="13976" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="12104" heatid="14017" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="12105" heatid="14043" lane="5" entrytime="00:02:19.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="12094">
              <RESULTS>
                <RESULT eventid="1062" points="296" reactiontime="+106" swimtime="00:00:35.60" resultid="12095" heatid="13899" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1147" points="293" reactiontime="+110" swimtime="00:12:13.56" resultid="12096" heatid="13936" lane="4" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="150" swimtime="00:02:11.90" />
                    <SPLIT distance="200" swimtime="00:02:58.49" />
                    <SPLIT distance="250" swimtime="00:03:45.45" />
                    <SPLIT distance="300" swimtime="00:04:32.13" />
                    <SPLIT distance="350" swimtime="00:05:18.92" />
                    <SPLIT distance="400" swimtime="00:06:05.40" />
                    <SPLIT distance="450" swimtime="00:06:52.22" />
                    <SPLIT distance="500" swimtime="00:07:38.29" />
                    <SPLIT distance="550" swimtime="00:08:24.86" />
                    <SPLIT distance="600" swimtime="00:09:11.24" />
                    <SPLIT distance="650" swimtime="00:09:57.77" />
                    <SPLIT distance="700" swimtime="00:10:44.16" />
                    <SPLIT distance="750" swimtime="00:11:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="294" reactiontime="+116" swimtime="00:01:18.22" resultid="12097" heatid="13974" lane="2" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="12098" heatid="14041" lane="2" entrytime="00:02:52.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="12099" heatid="14104" lane="1" entrytime="00:05:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="12106">
              <RESULTS>
                <RESULT eventid="1079" points="230" reactiontime="+95" swimtime="00:00:34.12" resultid="12107" heatid="13907" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1205" points="190" reactiontime="+83" swimtime="00:00:41.77" resultid="12108" heatid="13952" lane="0" entrytime="00:00:42.80" />
                <RESULT eventid="1406" points="201" reactiontime="+89" swimtime="00:01:38.73" resultid="12109" heatid="14007" lane="8" entrytime="00:01:40.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="12110" heatid="14091" lane="4" entrytime="00:00:42.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Victor" gender="M" lastname="Lyubavin" nation="RUS" athleteid="12111">
              <RESULTS>
                <RESULT eventid="1113" points="266" reactiontime="+91" swimtime="00:02:57.18" resultid="12112" heatid="13927" lane="1" entrytime="00:02:51.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="150" swimtime="00:02:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="311" reactiontime="+91" swimtime="00:03:07.35" resultid="12113" heatid="13968" lane="8" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:30.87" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="381" reactiontime="+81" swimtime="00:01:04.70" resultid="12114" heatid="13984" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="322" reactiontime="+84" swimtime="00:01:24.48" resultid="12115" heatid="14010" lane="7" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="12116" heatid="14022" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="12117" heatid="14094" lane="2" entrytime="00:00:37.50" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="12118" heatid="14111" lane="3" entrytime="00:05:19.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="14186" heatid="14100" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:15.92" />
                    <SPLIT distance="100" swimtime="00:02:02.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12100" number="1" />
                    <RELAYPOSITION athleteid="12106" number="2" />
                    <RELAYPOSITION athleteid="12111" number="3" />
                    <RELAYPOSITION athleteid="12094" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="12120" heatid="13933" lane="4" entrytime="00:02:09.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12100" number="1" />
                    <RELAYPOSITION athleteid="12111" number="2" />
                    <RELAYPOSITION athleteid="12106" number="3" />
                    <RELAYPOSITION athleteid="12094" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="11913" name="Redeco Wrocław">
          <CONTACT name="Wolny Dariusz" phone="603630870" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="11924">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1474" points="380" reactiontime="+80" swimtime="00:01:11.70" resultid="11925" heatid="14037" lane="1" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1647" points="358" reactiontime="+76" swimtime="00:02:37.61" resultid="11926" heatid="14081" lane="2" entrytime="00:02:35.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-31" firstname="Agata" gender="F" lastname="Szydło" nation="POL" athleteid="11936">
              <RESULTS>
                <RESULT eventid="1147" points="184" reactiontime="+104" swimtime="00:14:15.93" resultid="11937" heatid="13935" lane="4" entrytime="00:14:39.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:31.59" />
                    <SPLIT distance="100" swimtime="00:01:37.86" />
                    <SPLIT distance="150" swimtime="00:04:20.44" />
                    <SPLIT distance="200" swimtime="00:03:25.75" />
                    <SPLIT distance="250" swimtime="00:06:09.89" />
                    <SPLIT distance="300" swimtime="00:05:14.91" />
                    <SPLIT distance="350" swimtime="00:07:59.13" />
                    <SPLIT distance="400" swimtime="00:07:04.30" />
                    <SPLIT distance="450" swimtime="00:09:48.07" />
                    <SPLIT distance="500" swimtime="00:08:53.63" />
                    <SPLIT distance="550" swimtime="00:11:36.62" />
                    <SPLIT distance="600" swimtime="00:10:42.26" />
                    <SPLIT distance="650" swimtime="00:13:24.16" />
                    <SPLIT distance="700" swimtime="00:12:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="217" reactiontime="+110" swimtime="00:03:51.28" resultid="11938" heatid="13960" lane="2" entrytime="00:03:56.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="100" swimtime="00:01:52.10" />
                    <SPLIT distance="150" swimtime="00:02:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="173" reactiontime="+102" swimtime="00:01:33.32" resultid="11939" heatid="13971" lane="6" entrytime="00:01:41.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="195" reactiontime="+101" swimtime="00:01:50.88" resultid="11940" heatid="14001" lane="2" entrytime="00:01:50.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="172" swimtime="00:03:22.95" resultid="11941" heatid="14040" lane="9" entrytime="00:03:29.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:37.38" />
                    <SPLIT distance="150" swimtime="00:02:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="178" swimtime="00:00:52.31" resultid="11942" heatid="14084" lane="9" entrytime="00:00:52.99" />
                <RESULT eventid="1721" points="170" reactiontime="+103" swimtime="00:07:09.95" resultid="11943" heatid="14103" lane="8" entrytime="00:06:59.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:42.00" />
                    <SPLIT distance="150" swimtime="00:02:36.12" />
                    <SPLIT distance="200" swimtime="00:03:31.44" />
                    <SPLIT distance="250" swimtime="00:04:26.66" />
                    <SPLIT distance="300" swimtime="00:05:22.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Joanna" gender="F" lastname="Chojcan" nation="POL" athleteid="11927">
              <RESULTS>
                <RESULT eventid="1096" points="282" reactiontime="+86" swimtime="00:03:12.22" resultid="11928" heatid="13920" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:27.74" />
                    <SPLIT distance="150" swimtime="00:02:26.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="244" reactiontime="+89" swimtime="00:12:59.54" resultid="11929" heatid="13936" lane="6" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.56" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                    <SPLIT distance="200" swimtime="00:02:59.16" />
                    <SPLIT distance="250" swimtime="00:03:47.94" />
                    <SPLIT distance="300" swimtime="00:04:38.29" />
                    <SPLIT distance="350" swimtime="00:05:28.52" />
                    <SPLIT distance="400" swimtime="00:06:18.99" />
                    <SPLIT distance="450" swimtime="00:07:09.33" />
                    <SPLIT distance="500" swimtime="00:08:00.49" />
                    <SPLIT distance="550" swimtime="00:08:51.38" />
                    <SPLIT distance="600" swimtime="00:09:42.34" />
                    <SPLIT distance="650" swimtime="00:10:32.51" />
                    <SPLIT distance="700" swimtime="00:11:22.35" />
                    <SPLIT distance="750" swimtime="00:12:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="276" reactiontime="+66" swimtime="00:00:41.53" resultid="11930" heatid="13947" lane="8" entrytime="00:00:37.90" />
                <RESULT eventid="1324" points="171" reactiontime="+88" swimtime="00:03:39.07" resultid="11931" heatid="13991" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                    <SPLIT distance="100" swimtime="00:01:38.43" />
                    <SPLIT distance="150" swimtime="00:02:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="262" reactiontime="+73" swimtime="00:01:30.80" resultid="11932" heatid="14031" lane="9" entrytime="00:01:20.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="262" reactiontime="+91" swimtime="00:06:59.47" resultid="11933" heatid="14058" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                    <SPLIT distance="200" swimtime="00:03:24.90" />
                    <SPLIT distance="250" swimtime="00:04:25.10" />
                    <SPLIT distance="300" swimtime="00:05:25.82" />
                    <SPLIT distance="350" swimtime="00:06:13.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="219" reactiontime="+87" swimtime="00:01:32.22" resultid="11934" heatid="14065" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="274" reactiontime="+75" swimtime="00:03:10.87" resultid="11935" heatid="14074" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:32.22" />
                    <SPLIT distance="150" swimtime="00:02:21.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-14" firstname="Anna" gender="F" lastname="Jaśkiewicz" nation="POL" athleteid="11944">
              <RESULTS>
                <RESULT eventid="1062" points="321" reactiontime="+89" swimtime="00:00:34.65" resultid="11945" heatid="13899" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1147" points="209" reactiontime="+91" swimtime="00:13:40.50" resultid="11946" heatid="13936" lane="8" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:04:02.48" />
                    <SPLIT distance="200" swimtime="00:03:10.35" />
                    <SPLIT distance="250" swimtime="00:05:48.22" />
                    <SPLIT distance="300" swimtime="00:04:55.35" />
                    <SPLIT distance="350" swimtime="00:07:35.08" />
                    <SPLIT distance="400" swimtime="00:06:41.36" />
                    <SPLIT distance="450" swimtime="00:09:21.75" />
                    <SPLIT distance="500" swimtime="00:08:28.56" />
                    <SPLIT distance="550" swimtime="00:11:06.99" />
                    <SPLIT distance="600" swimtime="00:10:14.19" />
                    <SPLIT distance="700" swimtime="00:12:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="306" reactiontime="+98" swimtime="00:03:26.42" resultid="11947" heatid="13961" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:39.07" />
                    <SPLIT distance="150" swimtime="00:02:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="290" reactiontime="+95" swimtime="00:01:18.60" resultid="11948" heatid="13974" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="247" reactiontime="+89" swimtime="00:02:59.84" resultid="11949" heatid="14040" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="150" swimtime="00:02:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="302" reactiontime="+94" swimtime="00:00:43.93" resultid="11950" heatid="14085" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1721" points="220" reactiontime="+91" swimtime="00:06:34.70" resultid="11951" heatid="14103" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                    <SPLIT distance="200" swimtime="00:03:11.06" />
                    <SPLIT distance="250" swimtime="00:04:02.92" />
                    <SPLIT distance="300" swimtime="00:04:54.75" />
                    <SPLIT distance="350" swimtime="00:05:46.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMKS" nation="POL" region="SLA" clubid="11061" name="Rmks Rybnik">
          <CONTACT city="rybnik" email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" state="SLA" street="orzepowicka 22a/37" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="11062">
              <RESULTS>
                <RESULT eventid="1256" points="485" reactiontime="+81" swimtime="00:01:06.23" resultid="12377" heatid="13975" lane="5" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="418" reactiontime="+92" swimtime="00:00:32.65" resultid="12378" heatid="14017" lane="0" entrytime="00:00:33.50" />
                <RESULT eventid="1664" points="422" reactiontime="+90" swimtime="00:00:39.30" resultid="12379" heatid="14087" lane="1" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="11063">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1062" points="600" reactiontime="+79" swimtime="00:00:28.12" resultid="11064" heatid="13902" lane="4" entrytime="00:00:28.45" />
                <RESULT comment="Rekord Polski" eventid="1096" points="461" reactiontime="+86" swimtime="00:02:43.18" resultid="11065" heatid="13921" lane="3" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="413" reactiontime="+66" swimtime="00:00:36.31" resultid="11066" heatid="13946" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1324" points="311" reactiontime="+90" swimtime="00:02:59.70" resultid="11067" heatid="13991" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="150" swimtime="00:02:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1423" points="549" reactiontime="+83" swimtime="00:00:29.82" resultid="11068" heatid="14017" lane="4" entrytime="00:00:29.86" />
                <RESULT comment="Rekord Polski" eventid="1555" points="418" reactiontime="+92" swimtime="00:05:58.83" resultid="11069" heatid="14058" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="150" swimtime="00:02:05.56" />
                    <SPLIT distance="250" swimtime="00:03:48.43" />
                    <SPLIT distance="350" swimtime="00:05:21.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1595" points="516" reactiontime="+79" swimtime="00:01:09.33" resultid="11070" heatid="14065" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="406" reactiontime="+80" swimtime="00:00:39.80" resultid="11071" heatid="14085" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9861" name="Rydułtowska Akademia Aktywnego Seniora 60+" shortname="Rydułtowska Akademia Aktywnego">
          <CONTACT email="otelom.080966@interia.pl" name="OTLIK MARIAN" phone="692112775" state="SLONS" street="Wodzisław Śląski" zip="44300" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="9877">
              <RESULTS>
                <RESULT eventid="1079" points="76" reactiontime="+107" swimtime="00:00:49.28" resultid="9878" heatid="13904" lane="6" entrytime="00:00:46.00" />
                <RESULT comment="Z3 - Płynięcie podczas odcinku stylu dowolnego stylu grzbietowym, klasycznym lub motylkowym (Time: 17:19)" eventid="1113" reactiontime="+97" status="DSQ" swimtime="00:05:08.13" resultid="9879" heatid="13923" lane="8" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.20" />
                    <SPLIT distance="100" swimtime="00:02:24.06" />
                    <SPLIT distance="150" swimtime="00:03:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="68" reactiontime="+80" swimtime="00:00:58.69" resultid="9880" heatid="13950" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1341" points="38" reactiontime="+101" swimtime="00:05:29.93" resultid="9881" heatid="13992" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.94" />
                    <SPLIT distance="100" swimtime="00:02:31.52" />
                    <SPLIT distance="150" swimtime="00:04:00.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="48" reactiontime="+102" swimtime="00:01:01.69" resultid="9882" heatid="14019" lane="1" entrytime="00:00:56.00" />
                <RESULT eventid="1578" points="60" reactiontime="+101" swimtime="00:10:21.82" resultid="9883" heatid="14059" lane="6" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.17" />
                    <SPLIT distance="100" swimtime="00:02:37.17" />
                    <SPLIT distance="150" swimtime="00:03:57.89" />
                    <SPLIT distance="200" swimtime="00:05:18.28" />
                    <SPLIT distance="250" swimtime="00:06:41.46" />
                    <SPLIT distance="300" swimtime="00:08:02.53" />
                    <SPLIT distance="350" swimtime="00:09:13.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="40" reactiontime="+102" swimtime="00:02:25.34" resultid="9884" heatid="14066" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="66" reactiontime="+89" swimtime="00:04:36.77" resultid="9885" heatid="14077" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.15" />
                    <SPLIT distance="100" swimtime="00:02:18.51" />
                    <SPLIT distance="150" swimtime="00:03:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-21" firstname="Michał" gender="M" lastname="Kądzioła" nation="POL" athleteid="11758">
              <RESULTS>
                <RESULT eventid="1205" points="359" reactiontime="+74" swimtime="00:00:33.82" resultid="11759" heatid="13956" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1273" points="364" reactiontime="+102" swimtime="00:01:05.68" resultid="11760" heatid="13983" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="375" reactiontime="+88" swimtime="00:00:31.09" resultid="11761" heatid="14024" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="314" reactiontime="+72" swimtime="00:01:16.36" resultid="11762" heatid="14036" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11763" heatid="14081" lane="9" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="9886">
              <RESULTS>
                <RESULT eventid="1079" points="79" reactiontime="+116" swimtime="00:00:48.61" resultid="9887" heatid="13904" lane="7" entrytime="00:00:47.00" />
                <RESULT eventid="1113" points="61" reactiontime="+119" swimtime="00:04:49.16" resultid="9888" heatid="13922" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.30" />
                    <SPLIT distance="100" swimtime="00:02:26.75" />
                    <SPLIT distance="150" swimtime="00:03:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="66" reactiontime="+95" swimtime="00:00:59.22" resultid="9889" heatid="13949" lane="1" />
                <RESULT eventid="1273" points="65" swimtime="00:01:56.27" resultid="9890" heatid="13978" lane="9" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="71" reactiontime="+101" swimtime="00:02:19.40" resultid="9891" heatid="14005" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="51" reactiontime="+115" swimtime="00:04:34.07" resultid="9892" heatid="14045" lane="2" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.22" />
                    <SPLIT distance="100" swimtime="00:02:09.64" />
                    <SPLIT distance="150" swimtime="00:03:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="54" reactiontime="+82" swimtime="00:04:56.05" resultid="9893" heatid="14077" lane="8" entrytime="00:04:43.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.75" />
                    <SPLIT distance="100" swimtime="00:02:22.65" />
                    <SPLIT distance="150" swimtime="00:03:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="87" reactiontime="+82" swimtime="00:00:59.42" resultid="9894" heatid="14089" lane="7" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="9895">
              <RESULTS>
                <RESULT eventid="1079" points="326" reactiontime="+75" swimtime="00:00:30.37" resultid="9896" heatid="13911" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="216" reactiontime="+75" swimtime="00:03:09.82" resultid="9897" heatid="13925" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:29.81" />
                    <SPLIT distance="150" swimtime="00:02:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="184" reactiontime="+75" swimtime="00:03:43.19" resultid="9898" heatid="13963" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.10" />
                    <SPLIT distance="100" swimtime="00:01:45.76" />
                    <SPLIT distance="150" swimtime="00:02:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="303" reactiontime="+81" swimtime="00:01:09.82" resultid="9899" heatid="13982" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="236" reactiontime="+74" swimtime="00:00:36.26" resultid="9900" heatid="14021" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1578" points="183" reactiontime="+81" swimtime="00:07:08.95" resultid="9901" heatid="14059" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                    <SPLIT distance="150" swimtime="00:02:27.89" />
                    <SPLIT distance="200" swimtime="00:03:25.43" />
                    <SPLIT distance="250" swimtime="00:04:28.90" />
                    <SPLIT distance="300" swimtime="00:05:33.86" />
                    <SPLIT distance="350" swimtime="00:06:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="186" swimtime="00:01:27.26" resultid="9902" heatid="14066" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="200" reactiontime="+79" swimtime="00:00:45.12" resultid="9903" heatid="14091" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="9862">
              <RESULTS>
                <RESULT eventid="1113" points="161" reactiontime="+97" swimtime="00:03:29.17" resultid="9863" heatid="13924" lane="2" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="188" reactiontime="+99" swimtime="00:25:19.68" resultid="9864" heatid="13940" lane="3" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:32.01" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                    <SPLIT distance="200" swimtime="00:03:13.27" />
                    <SPLIT distance="250" swimtime="00:04:04.14" />
                    <SPLIT distance="300" swimtime="00:04:55.56" />
                    <SPLIT distance="350" swimtime="00:05:46.42" />
                    <SPLIT distance="400" swimtime="00:06:38.34" />
                    <SPLIT distance="450" swimtime="00:07:29.54" />
                    <SPLIT distance="500" swimtime="00:08:21.73" />
                    <SPLIT distance="550" swimtime="00:09:12.68" />
                    <SPLIT distance="600" swimtime="00:10:04.13" />
                    <SPLIT distance="650" swimtime="00:10:55.53" />
                    <SPLIT distance="700" swimtime="00:11:47.31" />
                    <SPLIT distance="750" swimtime="00:12:38.41" />
                    <SPLIT distance="800" swimtime="00:13:29.90" />
                    <SPLIT distance="850" swimtime="00:14:21.02" />
                    <SPLIT distance="900" swimtime="00:15:12.75" />
                    <SPLIT distance="950" swimtime="00:16:03.91" />
                    <SPLIT distance="1000" swimtime="00:16:55.15" />
                    <SPLIT distance="1050" swimtime="00:17:46.73" />
                    <SPLIT distance="1100" swimtime="00:18:38.69" />
                    <SPLIT distance="1150" swimtime="00:19:29.99" />
                    <SPLIT distance="1200" swimtime="00:20:21.39" />
                    <SPLIT distance="1250" swimtime="00:21:11.55" />
                    <SPLIT distance="1300" swimtime="00:22:02.62" />
                    <SPLIT distance="1350" swimtime="00:22:52.64" />
                    <SPLIT distance="1400" swimtime="00:23:43.29" />
                    <SPLIT distance="1450" swimtime="00:24:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="166" reactiontime="+85" swimtime="00:00:43.69" resultid="9865" heatid="13951" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1341" points="102" reactiontime="+92" swimtime="00:03:57.94" resultid="9866" heatid="13993" lane="0" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:48.19" />
                    <SPLIT distance="150" swimtime="00:02:52.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="9867" heatid="14034" lane="2" entrytime="00:01:33.00" />
                <RESULT eventid="1578" points="155" reactiontime="+95" swimtime="00:07:33.59" resultid="9868" heatid="14060" lane="8" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:46.25" />
                    <SPLIT distance="150" swimtime="00:04:49.73" />
                    <SPLIT distance="200" swimtime="00:03:43.95" />
                    <SPLIT distance="250" swimtime="00:06:44.35" />
                    <SPLIT distance="300" swimtime="00:05:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="152" reactiontime="+89" swimtime="00:01:33.15" resultid="9869" heatid="14067" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="133" reactiontime="+81" swimtime="00:03:39.02" resultid="9870" heatid="14079" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:46.68" />
                    <SPLIT distance="150" swimtime="00:02:44.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="9871">
              <RESULTS>
                <RESULT eventid="1205" points="12" reactiontime="+89" swimtime="00:01:42.73" resultid="9872" heatid="13949" lane="6" />
                <RESULT eventid="1273" points="30" reactiontime="+121" swimtime="00:02:30.83" resultid="9873" heatid="13977" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="12" reactiontime="+82" swimtime="00:03:44.84" resultid="9874" heatid="14032" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="28" reactiontime="+130" swimtime="00:05:34.21" resultid="9875" heatid="14045" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.57" />
                    <SPLIT distance="100" swimtime="00:02:36.65" />
                    <SPLIT distance="150" swimtime="00:04:06.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="16" reactiontime="+95" swimtime="00:07:23.14" resultid="9876" heatid="14076" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.59" />
                    <SPLIT distance="100" swimtime="00:03:38.08" />
                    <SPLIT distance="150" swimtime="00:05:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9653" name="Sikret Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@wp.pl" internet="www.sikret-plywanie.pl" name="Joanna Zagała" phone="601427257" street="Jagielońska 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="9661">
              <RESULTS>
                <RESULT eventid="1062" points="178" reactiontime="+80" swimtime="00:00:42.18" resultid="9662" heatid="13898" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1222" points="194" reactiontime="+84" swimtime="00:04:00.17" resultid="9663" heatid="13960" lane="8" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:01:57.90" />
                    <SPLIT distance="150" swimtime="00:03:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="45" reactiontime="+83" swimtime="00:05:40.52" resultid="9664" heatid="13990" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.67" />
                    <SPLIT distance="100" swimtime="00:02:20.29" />
                    <SPLIT distance="150" swimtime="00:03:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="173" reactiontime="+85" swimtime="00:01:55.27" resultid="9665" heatid="14001" lane="1" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="121" reactiontime="+96" swimtime="00:09:02.44" resultid="9666" heatid="14057" lane="3" entrytime="00:09:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:03:44.21" />
                    <SPLIT distance="200" swimtime="00:05:00.01" />
                    <SPLIT distance="250" swimtime="00:06:05.18" />
                    <SPLIT distance="300" swimtime="00:07:06.91" />
                    <SPLIT distance="350" swimtime="00:08:06.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="72" reactiontime="+82" swimtime="00:02:13.27" resultid="9667" heatid="14063" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="205" reactiontime="+80" swimtime="00:00:49.93" resultid="9668" heatid="14084" lane="0" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-03-14" firstname="Tomasz" gender="M" lastname="Bartosik" nation="POL" athleteid="9692">
              <RESULTS>
                <RESULT eventid="1079" points="402" reactiontime="+79" swimtime="00:00:28.31" resultid="9693" heatid="13913" lane="3" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="9685">
              <RESULTS>
                <RESULT eventid="1079" points="351" swimtime="00:00:29.63" resultid="9686" heatid="13911" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="250" reactiontime="+95" swimtime="00:03:00.82" resultid="9687" heatid="13925" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:18.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="9688" heatid="13955" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1440" points="356" reactiontime="+82" swimtime="00:00:31.64" resultid="9689" heatid="14022" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="9690" heatid="14035" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1744" points="251" reactiontime="+83" swimtime="00:05:48.45" resultid="9691" heatid="14109" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="200" swimtime="00:02:49.49" />
                    <SPLIT distance="300" swimtime="00:04:19.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="9669">
              <RESULTS>
                <RESULT eventid="1062" points="236" reactiontime="+76" swimtime="00:00:38.38" resultid="9670" heatid="13898" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1096" points="167" reactiontime="+84" swimtime="00:03:49.02" resultid="9671" heatid="13919" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                    <SPLIT distance="100" swimtime="00:01:57.13" />
                    <SPLIT distance="150" swimtime="00:02:59.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="183" swimtime="00:00:47.60" resultid="9672" heatid="13944" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1256" points="222" reactiontime="+76" swimtime="00:01:25.96" resultid="9673" heatid="13973" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="155" reactiontime="+80" swimtime="00:01:48.18" resultid="9674" heatid="14029" lane="1" entrytime="00:02:00.00" />
                <RESULT eventid="1491" points="199" reactiontime="+80" swimtime="00:03:13.41" resultid="9675" heatid="14039" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="150" swimtime="00:02:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="165" reactiontime="+87" swimtime="00:03:46.00" resultid="9676" heatid="14073" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                    <SPLIT distance="100" swimtime="00:03:46.23" />
                    <SPLIT distance="150" swimtime="00:02:50.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="202" reactiontime="+87" swimtime="00:00:50.24" resultid="9677" heatid="14083" lane="7" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="9654">
              <RESULTS>
                <RESULT eventid="1062" points="206" swimtime="00:00:40.17" resultid="9655" heatid="13898" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1222" points="223" reactiontime="+100" swimtime="00:03:49.39" resultid="9656" heatid="13960" lane="7" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.65" />
                    <SPLIT distance="100" swimtime="00:01:51.34" />
                    <SPLIT distance="150" swimtime="00:02:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="172" reactiontime="+103" swimtime="00:01:33.56" resultid="9657" heatid="13972" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="201" reactiontime="+100" swimtime="00:01:49.68" resultid="9658" heatid="14001" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="160" reactiontime="+100" swimtime="00:03:27.99" resultid="9659" heatid="14039" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:39.48" />
                    <SPLIT distance="150" swimtime="00:02:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="184" reactiontime="+102" swimtime="00:00:51.82" resultid="9660" heatid="14084" lane="8" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="9694">
              <RESULTS>
                <RESULT eventid="1079" points="205" reactiontime="+113" swimtime="00:00:35.43" resultid="9695" heatid="13906" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1205" points="171" reactiontime="+90" swimtime="00:00:43.30" resultid="9696" heatid="13953" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1273" points="189" reactiontime="+93" swimtime="00:01:21.67" resultid="9697" heatid="13979" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="153" reactiontime="+87" swimtime="00:01:37.06" resultid="9698" heatid="14034" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-15" firstname="Mieczysław" gender="M" lastname="Mydłowski" nation="POL" athleteid="9678">
              <RESULTS>
                <RESULT eventid="1079" points="284" reactiontime="+97" swimtime="00:00:31.81" resultid="9679" heatid="13908" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1205" points="232" reactiontime="+76" swimtime="00:00:39.08" resultid="9680" heatid="13953" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1273" points="281" reactiontime="+87" swimtime="00:01:11.54" resultid="9681" heatid="13981" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="259" reactiontime="+85" swimtime="00:01:30.76" resultid="9682" heatid="14008" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="200" reactiontime="+132" swimtime="00:01:28.71" resultid="9683" heatid="14035" lane="0" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="281" reactiontime="+86" swimtime="00:00:40.33" resultid="9684" heatid="14092" lane="0" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="285" reactiontime="+71" swimtime="00:02:21.96" resultid="9701" heatid="13998" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                    <SPLIT distance="100" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:01:53.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9694" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="9678" number="2" />
                    <RELAYPOSITION athleteid="9685" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="9692" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="329" reactiontime="+84" swimtime="00:02:02.89" resultid="9702" heatid="14055" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:33.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9692" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="9678" number="2" />
                    <RELAYPOSITION athleteid="9694" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="9685" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="204" reactiontime="+89" swimtime="00:02:24.03" resultid="9699" heatid="13933" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:01:55.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9678" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="9661" number="2" />
                    <RELAYPOSITION athleteid="9669" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="9692" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="172" reactiontime="+90" swimtime="00:02:47.68" resultid="9700" heatid="14100" lane="0" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.53" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:19.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9669" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="9661" number="2" />
                    <RELAYPOSITION athleteid="9678" number="3" reactiontime="-64" />
                    <RELAYPOSITION athleteid="9692" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11663" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="os. Stefana Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-01" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="11664">
              <RESULTS>
                <RESULT eventid="1062" points="353" reactiontime="+89" swimtime="00:00:33.57" resultid="11665" heatid="13899" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1147" points="278" reactiontime="+100" swimtime="00:12:26.01" resultid="11666" heatid="13936" lane="7" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:02:11.77" />
                    <SPLIT distance="200" swimtime="00:02:58.79" />
                    <SPLIT distance="250" swimtime="00:03:45.28" />
                    <SPLIT distance="300" swimtime="00:04:32.30" />
                    <SPLIT distance="350" swimtime="00:05:18.77" />
                    <SPLIT distance="400" swimtime="00:06:06.23" />
                    <SPLIT distance="450" swimtime="00:06:53.87" />
                    <SPLIT distance="500" swimtime="00:07:41.55" />
                    <SPLIT distance="550" swimtime="00:08:29.34" />
                    <SPLIT distance="600" swimtime="00:09:17.21" />
                    <SPLIT distance="650" swimtime="00:10:05.13" />
                    <SPLIT distance="750" swimtime="00:11:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="338" reactiontime="+96" swimtime="00:01:14.72" resultid="11667" heatid="13972" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="194" reactiontime="+100" swimtime="00:03:30.06" resultid="11668" heatid="13991" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:42.68" />
                    <SPLIT distance="150" swimtime="00:02:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="304" reactiontime="+94" swimtime="00:00:36.30" resultid="11669" heatid="14015" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1491" points="309" reactiontime="+96" swimtime="00:02:46.98" resultid="11670" heatid="14041" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:21.53" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="190" reactiontime="+103" swimtime="00:01:36.78" resultid="11671" heatid="14064" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="271" swimtime="00:06:08.19" resultid="11672" heatid="14104" lane="9" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                    <SPLIT distance="200" swimtime="00:03:04.06" />
                    <SPLIT distance="250" swimtime="00:03:50.18" />
                    <SPLIT distance="300" swimtime="00:04:37.60" />
                    <SPLIT distance="350" swimtime="00:05:23.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-01" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="11673">
              <RESULTS>
                <RESULT eventid="1096" points="407" reactiontime="+100" swimtime="00:02:50.11" resultid="11674" heatid="13921" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:02:09.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="354" reactiontime="+94" swimtime="00:11:28.74" resultid="11675" heatid="13937" lane="8" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:01.82" />
                    <SPLIT distance="200" swimtime="00:02:45.34" />
                    <SPLIT distance="250" swimtime="00:03:29.09" />
                    <SPLIT distance="300" swimtime="00:04:12.95" />
                    <SPLIT distance="350" swimtime="00:04:56.76" />
                    <SPLIT distance="400" swimtime="00:05:40.94" />
                    <SPLIT distance="450" swimtime="00:06:24.78" />
                    <SPLIT distance="500" swimtime="00:07:08.78" />
                    <SPLIT distance="550" swimtime="00:07:53.05" />
                    <SPLIT distance="600" swimtime="00:08:37.50" />
                    <SPLIT distance="650" swimtime="00:09:21.49" />
                    <SPLIT distance="700" swimtime="00:10:05.51" />
                    <SPLIT distance="750" swimtime="00:10:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="422" reactiontime="+79" swimtime="00:00:36.07" resultid="11676" heatid="13948" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1256" points="429" swimtime="00:01:09.02" resultid="11677" heatid="13976" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="439" reactiontime="+77" swimtime="00:01:16.45" resultid="11678" heatid="14029" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="401" reactiontime="+94" swimtime="00:02:33.15" resultid="11679" heatid="14042" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="150" swimtime="00:01:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="444" reactiontime="+76" swimtime="00:02:42.58" resultid="11680" heatid="14075" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:01.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="384" reactiontime="+96" swimtime="00:05:27.67" resultid="11681" heatid="14104" lane="4" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                    <SPLIT distance="150" swimtime="00:01:59.98" />
                    <SPLIT distance="200" swimtime="00:02:42.28" />
                    <SPLIT distance="250" swimtime="00:03:24.75" />
                    <SPLIT distance="300" swimtime="00:04:07.16" />
                    <SPLIT distance="350" swimtime="00:04:48.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-01" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="11682">
              <RESULTS>
                <RESULT eventid="1079" points="445" swimtime="00:00:27.38" resultid="11683" heatid="13914" lane="9" entrytime="00:00:27.50" />
                <RESULT eventid="1113" points="415" reactiontime="+83" swimtime="00:02:32.72" resultid="11684" heatid="13930" lane="6" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:13.25" />
                    <SPLIT distance="150" swimtime="00:01:58.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="501" reactiontime="+80" swimtime="00:00:59.04" resultid="11685" heatid="13988" lane="0" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="445" reactiontime="+81" swimtime="00:02:13.51" resultid="11686" heatid="14052" lane="5" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="366" reactiontime="+88" swimtime="00:05:40.75" resultid="11687" heatid="14062" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                    <SPLIT distance="200" swimtime="00:02:46.35" />
                    <SPLIT distance="250" swimtime="00:03:36.72" />
                    <SPLIT distance="300" swimtime="00:04:28.21" />
                    <SPLIT distance="350" swimtime="00:05:05.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="448" reactiontime="+69" swimtime="00:04:47.60" resultid="11688" heatid="14113" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:47.72" />
                    <SPLIT distance="200" swimtime="00:02:24.97" />
                    <SPLIT distance="250" swimtime="00:03:01.11" />
                    <SPLIT distance="300" swimtime="00:03:37.64" />
                    <SPLIT distance="350" swimtime="00:04:13.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-01" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="11698">
              <RESULTS>
                <RESULT eventid="1079" points="495" reactiontime="+78" swimtime="00:00:26.42" resultid="11699" heatid="13913" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="11700" heatid="13930" lane="0" entrytime="00:02:35.00" />
                <RESULT eventid="1205" points="457" reactiontime="+76" swimtime="00:00:31.19" resultid="11701" heatid="13956" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="518" reactiontime="+79" swimtime="00:00:58.38" resultid="11702" heatid="13986" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="503" reactiontime="+79" swimtime="00:00:28.19" resultid="11703" heatid="14019" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1474" points="451" swimtime="00:01:07.68" resultid="11704" heatid="14037" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="463" swimtime="00:01:04.39" resultid="11705" heatid="14068" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11706" heatid="14082" lane="9" entrytime="00:02:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-06-01" firstname="Łukasz" gender="M" lastname="Beszterda" nation="POL" athleteid="11689">
              <RESULTS>
                <RESULT eventid="1079" points="403" reactiontime="+104" swimtime="00:00:28.30" resultid="11690" heatid="13913" lane="7" entrytime="00:00:28.00" />
                <RESULT comment="(Time: 21:28), Przekroczony regulaminowy limit czasu." eventid="1165" reactiontime="+115" status="OTL" swimtime="00:20:10.58" resultid="11691" heatid="13943" lane="8" entrytime="00:19:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:46.91" />
                    <SPLIT distance="200" swimtime="00:02:25.73" />
                    <SPLIT distance="250" swimtime="00:03:04.87" />
                    <SPLIT distance="300" swimtime="00:03:45.02" />
                    <SPLIT distance="350" swimtime="00:04:25.31" />
                    <SPLIT distance="400" swimtime="00:05:05.78" />
                    <SPLIT distance="450" swimtime="00:05:46.98" />
                    <SPLIT distance="500" swimtime="00:06:27.93" />
                    <SPLIT distance="550" swimtime="00:07:08.99" />
                    <SPLIT distance="600" swimtime="00:07:50.08" />
                    <SPLIT distance="650" swimtime="00:08:30.85" />
                    <SPLIT distance="700" swimtime="00:09:12.33" />
                    <SPLIT distance="750" swimtime="00:09:53.69" />
                    <SPLIT distance="800" swimtime="00:10:34.84" />
                    <SPLIT distance="850" swimtime="00:11:16.35" />
                    <SPLIT distance="900" swimtime="00:11:57.90" />
                    <SPLIT distance="950" swimtime="00:12:39.31" />
                    <SPLIT distance="1000" swimtime="00:13:20.82" />
                    <SPLIT distance="1050" swimtime="00:14:01.62" />
                    <SPLIT distance="1100" swimtime="00:14:42.98" />
                    <SPLIT distance="1150" swimtime="00:15:24.26" />
                    <SPLIT distance="1200" swimtime="00:16:06.04" />
                    <SPLIT distance="1250" swimtime="00:16:47.42" />
                    <SPLIT distance="1300" swimtime="00:17:28.34" />
                    <SPLIT distance="1350" swimtime="00:18:09.63" />
                    <SPLIT distance="1400" swimtime="00:18:50.58" />
                    <SPLIT distance="1450" swimtime="00:19:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="294" reactiontime="+71" swimtime="00:00:36.14" resultid="11692" heatid="13957" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="399" reactiontime="+108" swimtime="00:01:03.67" resultid="11693" heatid="13987" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="326" reactiontime="+99" swimtime="00:00:32.56" resultid="11694" heatid="14023" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1508" points="368" swimtime="00:02:22.28" resultid="11695" heatid="14053" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="328" reactiontime="+101" swimtime="00:00:38.29" resultid="11696" heatid="14096" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1744" points="374" reactiontime="+102" swimtime="00:05:05.33" resultid="11697" heatid="14114" lane="8" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:49.23" />
                    <SPLIT distance="200" swimtime="00:02:28.71" />
                    <SPLIT distance="250" swimtime="00:03:08.81" />
                    <SPLIT distance="300" swimtime="00:03:49.22" />
                    <SPLIT distance="350" swimtime="00:04:28.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="11102" name="Steef">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" phone="500388374" state="DOL" street="Edyty Stein 6" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="11111">
              <RESULTS>
                <RESULT eventid="1165" points="190" reactiontime="+109" swimtime="00:25:15.01" resultid="11112" heatid="13940" lane="1" entrytime="00:25:26.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:33.79" />
                    <SPLIT distance="150" swimtime="00:02:23.30" />
                    <SPLIT distance="200" swimtime="00:03:12.86" />
                    <SPLIT distance="250" swimtime="00:04:02.99" />
                    <SPLIT distance="300" swimtime="00:04:52.19" />
                    <SPLIT distance="350" swimtime="00:05:42.34" />
                    <SPLIT distance="400" swimtime="00:06:33.85" />
                    <SPLIT distance="450" swimtime="00:07:23.98" />
                    <SPLIT distance="500" swimtime="00:08:14.00" />
                    <SPLIT distance="550" swimtime="00:09:04.63" />
                    <SPLIT distance="600" swimtime="00:09:55.99" />
                    <SPLIT distance="650" swimtime="00:10:49.60" />
                    <SPLIT distance="700" swimtime="00:11:40.23" />
                    <SPLIT distance="750" swimtime="00:12:32.47" />
                    <SPLIT distance="800" swimtime="00:13:24.05" />
                    <SPLIT distance="850" swimtime="00:14:16.12" />
                    <SPLIT distance="900" swimtime="00:15:06.13" />
                    <SPLIT distance="950" swimtime="00:15:56.67" />
                    <SPLIT distance="1000" swimtime="00:16:47.60" />
                    <SPLIT distance="1050" swimtime="00:17:38.82" />
                    <SPLIT distance="1100" swimtime="00:18:29.76" />
                    <SPLIT distance="1150" swimtime="00:19:21.64" />
                    <SPLIT distance="1200" swimtime="00:20:12.76" />
                    <SPLIT distance="1250" swimtime="00:21:05.04" />
                    <SPLIT distance="1300" swimtime="00:21:56.49" />
                    <SPLIT distance="1350" swimtime="00:22:47.01" />
                    <SPLIT distance="1400" swimtime="00:23:37.37" />
                    <SPLIT distance="1450" swimtime="00:24:28.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="126" reactiontime="+102" swimtime="00:03:42.23" resultid="11113" heatid="13993" lane="5" entrytime="00:03:30.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                    <SPLIT distance="100" swimtime="00:01:45.19" />
                    <SPLIT distance="150" swimtime="00:02:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="206" reactiontime="+106" swimtime="00:02:52.60" resultid="11114" heatid="14047" lane="6" entrytime="00:02:50.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                    <SPLIT distance="150" swimtime="00:02:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="153" reactiontime="+106" swimtime="00:07:35.74" resultid="11115" heatid="14060" lane="3" entrytime="00:06:45.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.16" />
                    <SPLIT distance="100" swimtime="00:01:45.41" />
                    <SPLIT distance="150" swimtime="00:02:48.48" />
                    <SPLIT distance="200" swimtime="00:03:49.06" />
                    <SPLIT distance="250" swimtime="00:04:52.33" />
                    <SPLIT distance="300" swimtime="00:05:56.81" />
                    <SPLIT distance="350" swimtime="00:06:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="128" swimtime="00:01:38.75" resultid="11116" heatid="14068" lane="9" entrytime="00:01:30.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="209" reactiontime="+110" swimtime="00:06:10.55" resultid="11117" heatid="14109" lane="2" entrytime="00:06:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:29.24" />
                    <SPLIT distance="150" swimtime="00:02:17.74" />
                    <SPLIT distance="200" swimtime="00:03:06.55" />
                    <SPLIT distance="250" swimtime="00:03:52.27" />
                    <SPLIT distance="300" swimtime="00:04:39.12" />
                    <SPLIT distance="350" swimtime="00:05:26.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="11103">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1096" points="330" reactiontime="+90" swimtime="00:03:02.46" resultid="11104" heatid="13920" lane="6" entrytime="00:03:04.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="286" swimtime="00:12:19.36" resultid="11105" heatid="13937" lane="9" entrytime="00:12:13.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:11.00" />
                    <SPLIT distance="200" swimtime="00:02:56.91" />
                    <SPLIT distance="250" swimtime="00:03:43.74" />
                    <SPLIT distance="300" swimtime="00:04:30.41" />
                    <SPLIT distance="350" swimtime="00:05:16.97" />
                    <SPLIT distance="400" swimtime="00:06:03.58" />
                    <SPLIT distance="450" swimtime="00:06:50.87" />
                    <SPLIT distance="500" swimtime="00:07:38.36" />
                    <SPLIT distance="550" swimtime="00:08:24.94" />
                    <SPLIT distance="600" swimtime="00:09:12.43" />
                    <SPLIT distance="650" swimtime="00:09:59.47" />
                    <SPLIT distance="700" swimtime="00:10:46.88" />
                    <SPLIT distance="750" swimtime="00:11:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1324" points="224" reactiontime="+102" swimtime="00:03:20.37" resultid="11106" heatid="13991" lane="7" entrytime="00:03:19.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                    <SPLIT distance="150" swimtime="00:02:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="306" reactiontime="+80" swimtime="00:01:26.21" resultid="11107" heatid="14030" lane="6" entrytime="00:01:26.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="318" reactiontime="+101" swimtime="00:06:33.20" resultid="11108" heatid="14058" lane="1" entrytime="00:06:21.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:33.08" />
                    <SPLIT distance="150" swimtime="00:02:22.43" />
                    <SPLIT distance="200" swimtime="00:03:11.96" />
                    <SPLIT distance="250" swimtime="00:04:07.63" />
                    <SPLIT distance="300" swimtime="00:05:03.74" />
                    <SPLIT distance="350" swimtime="00:05:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="304" reactiontime="+80" swimtime="00:03:04.33" resultid="11109" heatid="14074" lane="6" entrytime="00:03:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:17.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="269" reactiontime="+98" swimtime="00:06:08.91" resultid="11110" heatid="14104" lane="5" entrytime="00:05:51.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:02:12.29" />
                    <SPLIT distance="200" swimtime="00:02:59.95" />
                    <SPLIT distance="250" swimtime="00:03:47.24" />
                    <SPLIT distance="300" swimtime="00:04:34.01" />
                    <SPLIT distance="350" swimtime="00:05:21.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" nation="POL" region="KR" clubid="11490" name="Straż Miejska Miasta Kraków">
          <CONTACT city="KRAKÓW" name="JAWIEŃ" phone="505593911" state="MAŁ" street="kRZYSZTOF" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-11" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="11505">
              <RESULTS>
                <RESULT eventid="1113" points="294" swimtime="00:02:51.32" resultid="11506" heatid="13927" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:07.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="327" reactiontime="+85" swimtime="00:03:04.29" resultid="11507" heatid="13964" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:28.25" />
                    <SPLIT distance="150" swimtime="00:02:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="208" reactiontime="+87" swimtime="00:03:07.97" resultid="11508" heatid="13995" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="331" reactiontime="+80" swimtime="00:01:23.67" resultid="11509" heatid="14011" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="292" reactiontime="+76" swimtime="00:06:07.35" resultid="11510" heatid="14061" lane="7" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:18.16" />
                    <SPLIT distance="150" swimtime="00:02:09.54" />
                    <SPLIT distance="200" swimtime="00:03:00.03" />
                    <SPLIT distance="250" swimtime="00:03:48.65" />
                    <SPLIT distance="300" swimtime="00:04:39.57" />
                    <SPLIT distance="350" swimtime="00:05:24.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="280" reactiontime="+77" swimtime="00:01:16.14" resultid="11511" heatid="14066" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 11:02)" eventid="1681" reactiontime="+68" status="DSQ" swimtime="00:00:38.21" resultid="11512" heatid="14094" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WA" clubid="12313" name="Swimmers St. Pływackie">
          <CONTACT city="WARSZAWA" email="REMOG@SWIMMERSTEAM.PL" internet="WWW.SWIMMERSTEAM.PL" name="GOŁĘBIOWSKI REMIGIUSZ" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-27" firstname="Remigiusz" gender="M" lastname="Miklewski" nation="POL" athleteid="12331">
              <RESULTS>
                <RESULT eventid="1079" points="356" reactiontime="+72" swimtime="00:00:29.48" resultid="12332" heatid="13912" lane="2" entrytime="00:00:28.70" />
                <RESULT eventid="1273" points="281" reactiontime="+76" swimtime="00:01:11.57" resultid="12333" heatid="13982" lane="0" entrytime="00:01:10.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="288" reactiontime="+79" swimtime="00:00:33.94" resultid="12334" heatid="14023" lane="8" entrytime="00:00:32.70" />
                <RESULT eventid="1681" points="252" reactiontime="+79" swimtime="00:00:41.81" resultid="12335" heatid="14093" lane="2" entrytime="00:00:38.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="12314">
              <RESULTS>
                <RESULT eventid="1079" points="472" reactiontime="+75" swimtime="00:00:26.85" resultid="12315" heatid="13915" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1165" points="467" reactiontime="+83" swimtime="00:18:42.59" resultid="12316" heatid="13943" lane="6" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:45.13" />
                    <SPLIT distance="200" swimtime="00:02:21.82" />
                    <SPLIT distance="250" swimtime="00:02:58.78" />
                    <SPLIT distance="300" swimtime="00:03:35.52" />
                    <SPLIT distance="350" swimtime="00:04:12.11" />
                    <SPLIT distance="400" swimtime="00:04:48.74" />
                    <SPLIT distance="450" swimtime="00:05:25.32" />
                    <SPLIT distance="500" swimtime="00:06:02.39" />
                    <SPLIT distance="550" swimtime="00:06:39.27" />
                    <SPLIT distance="600" swimtime="00:07:16.89" />
                    <SPLIT distance="650" swimtime="00:07:54.19" />
                    <SPLIT distance="700" swimtime="00:08:32.10" />
                    <SPLIT distance="750" swimtime="00:09:10.14" />
                    <SPLIT distance="800" swimtime="00:09:48.82" />
                    <SPLIT distance="850" swimtime="00:10:26.93" />
                    <SPLIT distance="900" swimtime="00:11:05.53" />
                    <SPLIT distance="950" swimtime="00:11:43.69" />
                    <SPLIT distance="1000" swimtime="00:12:22.72" />
                    <SPLIT distance="1050" swimtime="00:13:00.90" />
                    <SPLIT distance="1100" swimtime="00:13:39.47" />
                    <SPLIT distance="1150" swimtime="00:14:17.67" />
                    <SPLIT distance="1200" swimtime="00:14:56.31" />
                    <SPLIT distance="1250" swimtime="00:15:34.42" />
                    <SPLIT distance="1300" swimtime="00:16:12.83" />
                    <SPLIT distance="1350" swimtime="00:16:50.69" />
                    <SPLIT distance="1400" swimtime="00:17:28.82" />
                    <SPLIT distance="1450" swimtime="00:18:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="494" reactiontime="+74" swimtime="00:00:59.32" resultid="12317" heatid="13988" lane="6" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="498" swimtime="00:00:28.29" resultid="12318" heatid="14027" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1508" points="464" reactiontime="+78" swimtime="00:02:11.67" resultid="12319" heatid="14053" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="470" reactiontime="+75" swimtime="00:01:04.07" resultid="12320" heatid="14071" lane="1" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="469" reactiontime="+76" swimtime="00:04:43.23" resultid="12321" heatid="14114" lane="7" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:43.40" />
                    <SPLIT distance="200" swimtime="00:02:20.14" />
                    <SPLIT distance="250" swimtime="00:02:56.92" />
                    <SPLIT distance="300" swimtime="00:03:33.17" />
                    <SPLIT distance="350" swimtime="00:04:09.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brozyna" nation="POL" athleteid="12336">
              <RESULTS>
                <RESULT eventid="1205" points="340" reactiontime="+78" swimtime="00:00:34.44" resultid="12337" heatid="13956" lane="2" entrytime="00:00:33.70" />
                <RESULT eventid="1474" points="325" reactiontime="+79" swimtime="00:01:15.53" resultid="12338" heatid="14037" lane="9" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="313" reactiontime="+65" swimtime="00:02:44.81" resultid="12339" heatid="14081" lane="8" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:19.26" />
                    <SPLIT distance="150" swimtime="00:02:02.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="12360">
              <RESULTS>
                <RESULT eventid="1113" points="563" reactiontime="+70" swimtime="00:02:17.98" resultid="12361" heatid="13931" lane="5" entrytime="00:02:17.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="639" reactiontime="+71" swimtime="00:02:27.41" resultid="12362" heatid="13970" lane="4" entrytime="00:02:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="588" reactiontime="+71" swimtime="00:01:09.13" resultid="12363" heatid="14013" lane="5" entrytime="00:01:08.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="533" reactiontime="+78" swimtime="00:05:00.67" resultid="12364" heatid="14062" lane="6" entrytime="00:05:14.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:52.21" />
                    <SPLIT distance="200" swimtime="00:02:33.85" />
                    <SPLIT distance="250" swimtime="00:03:12.73" />
                    <SPLIT distance="300" swimtime="00:03:51.76" />
                    <SPLIT distance="350" swimtime="00:04:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="576" reactiontime="+58" swimtime="00:00:31.75" resultid="12365" heatid="14098" lane="3" entrytime="00:00:30.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-03" firstname="Bolesław" gender="M" lastname="Porolniczak" nation="POL" athleteid="12349">
              <RESULTS>
                <RESULT eventid="1079" points="450" reactiontime="+83" swimtime="00:00:27.28" resultid="12350" heatid="13913" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1205" points="259" reactiontime="+78" swimtime="00:00:37.67" resultid="12351" heatid="13955" lane="3" entrytime="00:00:34.70" />
                <RESULT eventid="1273" points="431" reactiontime="+87" swimtime="00:01:02.09" resultid="12352" heatid="13985" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="366" reactiontime="+87" swimtime="00:00:31.35" resultid="12353" heatid="14025" lane="8" entrytime="00:00:30.70" />
                <RESULT eventid="1508" points="348" reactiontime="+102" swimtime="00:02:24.99" resultid="12354" heatid="14052" lane="1" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:10.07" />
                    <SPLIT distance="150" swimtime="00:01:47.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba" nation="POL" athleteid="12355">
              <RESULTS>
                <RESULT eventid="1062" points="418" reactiontime="+84" swimtime="00:00:31.72" resultid="12356" heatid="13901" lane="5" entrytime="00:00:31.35" />
                <RESULT eventid="1256" points="354" reactiontime="+85" swimtime="00:01:13.57" resultid="12357" heatid="13975" lane="2" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="336" reactiontime="+88" swimtime="00:00:35.13" resultid="12358" heatid="14016" lane="3" entrytime="00:00:35.78" />
                <RESULT eventid="1595" points="221" reactiontime="+94" swimtime="00:01:31.91" resultid="12359" heatid="14064" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-11" firstname="Mikołaj" gender="M" lastname="Tusiński" nation="POL" athleteid="12340">
              <RESULTS>
                <RESULT eventid="1079" points="427" reactiontime="+85" swimtime="00:00:27.75" resultid="12341" heatid="13914" lane="0" entrytime="00:00:27.40" />
                <RESULT comment="(Time: 21:07), Przekroczony regulaminowy limit czasu." eventid="1165" status="OTL" swimtime="00:21:34.56" resultid="12342" heatid="13942" lane="9" entrytime="00:21:55.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:58.50" />
                    <SPLIT distance="200" swimtime="00:02:41.06" />
                    <SPLIT distance="250" swimtime="00:03:25.65" />
                    <SPLIT distance="300" swimtime="00:04:09.94" />
                    <SPLIT distance="350" swimtime="00:04:54.96" />
                    <SPLIT distance="400" swimtime="00:05:39.96" />
                    <SPLIT distance="450" swimtime="00:06:25.09" />
                    <SPLIT distance="500" swimtime="00:07:09.82" />
                    <SPLIT distance="550" swimtime="00:07:55.10" />
                    <SPLIT distance="600" swimtime="00:08:40.31" />
                    <SPLIT distance="650" swimtime="00:09:25.52" />
                    <SPLIT distance="700" swimtime="00:10:10.11" />
                    <SPLIT distance="750" swimtime="00:10:54.55" />
                    <SPLIT distance="800" swimtime="00:11:38.70" />
                    <SPLIT distance="850" swimtime="00:12:20.74" />
                    <SPLIT distance="900" swimtime="00:13:03.10" />
                    <SPLIT distance="950" swimtime="00:13:45.54" />
                    <SPLIT distance="1000" swimtime="00:14:29.49" />
                    <SPLIT distance="1050" swimtime="00:15:12.83" />
                    <SPLIT distance="1100" swimtime="00:15:56.16" />
                    <SPLIT distance="1150" swimtime="00:16:39.24" />
                    <SPLIT distance="1200" swimtime="00:17:24.30" />
                    <SPLIT distance="1250" swimtime="00:18:08.15" />
                    <SPLIT distance="1300" swimtime="00:18:49.48" />
                    <SPLIT distance="1350" swimtime="00:19:34.02" />
                    <SPLIT distance="1400" swimtime="00:20:17.12" />
                    <SPLIT distance="1450" swimtime="00:20:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="12343" heatid="13955" lane="6" entrytime="00:00:34.89" />
                <RESULT eventid="1273" points="451" reactiontime="+86" swimtime="00:01:01.17" resultid="12344" heatid="13987" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="413" swimtime="00:00:30.10" resultid="12345" heatid="14024" lane="6" entrytime="00:00:31.15" />
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 18:58)" eventid="1508" reactiontime="+54" status="DSQ" swimtime="00:02:19.81" resultid="12346" heatid="14052" lane="3" entrytime="00:02:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="12347" heatid="14070" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="12348" heatid="14113" lane="2" entrytime="00:04:54.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="12366">
              <RESULTS>
                <RESULT eventid="1079" points="503" reactiontime="+71" swimtime="00:00:26.28" resultid="12367" heatid="13916" lane="5" entrytime="00:00:25.85" />
                <RESULT eventid="1113" points="312" reactiontime="+89" swimtime="00:02:47.91" resultid="12368" heatid="13926" lane="0" entrytime="00:03:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="320" reactiontime="+73" swimtime="00:00:35.12" resultid="12369" heatid="13954" lane="7" entrytime="00:00:36.53" />
                <RESULT eventid="1273" points="485" swimtime="00:00:59.67" resultid="12370" heatid="13988" lane="9" entrytime="00:00:58.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="441" reactiontime="+80" swimtime="00:00:29.46" resultid="12371" heatid="14025" lane="4" entrytime="00:00:29.15" />
                <RESULT eventid="1508" points="331" reactiontime="+83" swimtime="00:02:27.41" resultid="12372" heatid="14051" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="12373" heatid="14071" lane="0" entrytime="00:01:03.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="12374" heatid="14095" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="Tchorzewski" nation="POL" athleteid="12322">
              <RESULTS>
                <RESULT eventid="1113" points="254" reactiontime="+94" swimtime="00:02:59.83" resultid="12323" heatid="13926" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:23.38" />
                    <SPLIT distance="150" swimtime="00:02:20.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="242" reactiontime="+117" swimtime="00:23:16.41" resultid="12324" heatid="13941" lane="3" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:21.67" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                    <SPLIT distance="200" swimtime="00:02:51.40" />
                    <SPLIT distance="250" swimtime="00:03:37.74" />
                    <SPLIT distance="300" swimtime="00:04:24.60" />
                    <SPLIT distance="350" swimtime="00:05:11.62" />
                    <SPLIT distance="400" swimtime="00:05:58.78" />
                    <SPLIT distance="450" swimtime="00:06:45.88" />
                    <SPLIT distance="500" swimtime="00:07:32.50" />
                    <SPLIT distance="550" swimtime="00:08:20.28" />
                    <SPLIT distance="600" swimtime="00:09:07.75" />
                    <SPLIT distance="650" swimtime="00:09:55.83" />
                    <SPLIT distance="700" swimtime="00:10:44.06" />
                    <SPLIT distance="750" swimtime="00:11:30.87" />
                    <SPLIT distance="800" swimtime="00:12:17.16" />
                    <SPLIT distance="850" swimtime="00:13:04.70" />
                    <SPLIT distance="900" swimtime="00:13:51.53" />
                    <SPLIT distance="950" swimtime="00:14:39.95" />
                    <SPLIT distance="1000" swimtime="00:15:27.45" />
                    <SPLIT distance="1050" swimtime="00:16:15.66" />
                    <SPLIT distance="1100" swimtime="00:17:03.28" />
                    <SPLIT distance="1150" swimtime="00:17:51.19" />
                    <SPLIT distance="1200" swimtime="00:18:38.98" />
                    <SPLIT distance="1250" swimtime="00:19:25.94" />
                    <SPLIT distance="1300" swimtime="00:20:14.01" />
                    <SPLIT distance="1350" swimtime="00:21:01.27" />
                    <SPLIT distance="1400" swimtime="00:21:48.58" />
                    <SPLIT distance="1450" swimtime="00:22:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="309" reactiontime="+90" swimtime="00:01:09.33" resultid="12325" heatid="13982" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="182" reactiontime="+91" swimtime="00:03:16.76" resultid="12326" heatid="13994" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:02:21.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="265" reactiontime="+99" swimtime="00:02:38.63" resultid="12327" heatid="14049" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:00.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="208" reactiontime="+113" swimtime="00:06:51.31" resultid="12328" heatid="14060" lane="2" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:33.03" />
                    <SPLIT distance="150" swimtime="00:02:27.66" />
                    <SPLIT distance="200" swimtime="00:03:25.62" />
                    <SPLIT distance="250" swimtime="00:04:27.21" />
                    <SPLIT distance="300" swimtime="00:05:26.41" />
                    <SPLIT distance="350" swimtime="00:06:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="221" reactiontime="+64" swimtime="00:01:22.28" resultid="12329" heatid="14069" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="259" reactiontime="+100" swimtime="00:05:44.96" resultid="12330" heatid="14111" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="150" swimtime="00:02:03.85" />
                    <SPLIT distance="200" swimtime="00:02:48.16" />
                    <SPLIT distance="250" swimtime="00:03:33.30" />
                    <SPLIT distance="300" swimtime="00:04:19.17" />
                    <SPLIT distance="350" swimtime="00:05:05.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="402" reactiontime="+76" swimtime="00:02:06.58" resultid="12375" heatid="13999" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="150" swimtime="00:01:39.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12336" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="12366" number="2" />
                    <RELAYPOSITION athleteid="12314" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="12349" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="441" reactiontime="+85" swimtime="00:01:51.41" resultid="12376" heatid="14056" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="100" swimtime="00:00:54.58" />
                    <SPLIT distance="150" swimtime="00:01:25.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12314" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="12349" number="2" />
                    <RELAYPOSITION athleteid="12322" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="12366" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10104" name="Swimming Masters Team Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="10114">
              <RESULTS>
                <RESULT eventid="1079" points="315" reactiontime="+81" swimtime="00:00:30.71" resultid="10115" heatid="13910" lane="7" entrytime="00:00:30.61" entrycourse="LCM" />
                <RESULT eventid="1273" points="268" reactiontime="+76" swimtime="00:01:12.74" resultid="10116" heatid="13980" lane="6" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="203" reactiontime="+88" swimtime="00:02:53.55" resultid="10117" heatid="14047" lane="0" entrytime="00:02:55.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:23.09" />
                    <SPLIT distance="150" swimtime="00:02:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="182" swimtime="00:06:28.07" resultid="10118" heatid="14109" lane="9" entrytime="00:06:29.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                    <SPLIT distance="200" swimtime="00:03:04.96" />
                    <SPLIT distance="250" swimtime="00:03:55.93" />
                    <SPLIT distance="300" swimtime="00:04:48.53" />
                    <SPLIT distance="350" swimtime="00:05:40.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="10119">
              <RESULTS>
                <RESULT eventid="1079" points="432" reactiontime="+82" swimtime="00:00:27.64" resultid="10120" heatid="13910" lane="3" entrytime="00:00:30.50" entrycourse="LCM" />
                <RESULT eventid="1273" points="404" reactiontime="+81" swimtime="00:01:03.42" resultid="10121" heatid="13983" lane="5" entrytime="00:01:05.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="397" reactiontime="+84" swimtime="00:00:30.51" resultid="10122" heatid="14022" lane="2" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1613" points="304" reactiontime="+89" swimtime="00:01:14.04" resultid="10123" heatid="14070" lane="2" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="426" swimtime="00:00:35.10" resultid="10124" heatid="14095" lane="6" entrytime="00:00:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="10132">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="10133" heatid="13902" lane="7" entrytime="00:00:29.30" entrycourse="LCM" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="10134" heatid="13921" lane="2" entrytime="00:02:45.00" entrycourse="LCM" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="10135" heatid="13948" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="10136" heatid="14031" lane="5" entrytime="00:01:12.00" entrycourse="LCM" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="10137" heatid="14075" lane="3" entrytime="00:02:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-07" firstname="Marta" gender="F" lastname="Pachuc" nation="POL" athleteid="10152">
              <RESULTS>
                <RESULT eventid="1062" points="356" swimtime="00:00:33.48" resultid="10153" heatid="13901" lane="9" entrytime="00:00:32.08" entrycourse="LCM" />
                <RESULT eventid="1187" points="305" reactiontime="+77" swimtime="00:00:40.19" resultid="10154" heatid="13947" lane="4" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="326" swimtime="00:01:15.58" resultid="10155" heatid="13974" lane="9" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="255" reactiontime="+94" swimtime="00:01:41.39" resultid="10156" heatid="14002" lane="1" entrytime="00:01:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="255" reactiontime="+86" swimtime="00:00:46.45" resultid="10157" heatid="14085" lane="5" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="10145">
              <RESULTS>
                <RESULT eventid="1079" points="481" reactiontime="+79" swimtime="00:00:26.67" resultid="10146" heatid="13915" lane="6" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1113" points="418" reactiontime="+86" swimtime="00:02:32.45" resultid="10147" heatid="13930" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="512" reactiontime="+82" swimtime="00:00:58.60" resultid="10148" heatid="13988" lane="3" entrytime="00:00:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="443" reactiontime="+80" swimtime="00:00:29.42" resultid="10149" heatid="14025" lane="7" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1578" points="358" reactiontime="+86" swimtime="00:05:43.10" resultid="10150" heatid="14062" lane="8" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:58.54" />
                    <SPLIT distance="200" swimtime="00:02:43.52" />
                    <SPLIT distance="250" swimtime="00:03:32.97" />
                    <SPLIT distance="300" swimtime="00:04:24.07" />
                    <SPLIT distance="350" swimtime="00:05:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="393" reactiontime="+88" swimtime="00:05:00.31" resultid="10151" heatid="14112" lane="3" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:08.89" />
                    <SPLIT distance="150" swimtime="00:01:46.24" />
                    <SPLIT distance="200" swimtime="00:02:24.48" />
                    <SPLIT distance="250" swimtime="00:03:03.27" />
                    <SPLIT distance="300" swimtime="00:03:42.73" />
                    <SPLIT distance="350" swimtime="00:04:22.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-11-03" firstname="Agnieszka" gender="F" lastname="Suwiczak" nation="POL" athleteid="10125">
              <RESULTS>
                <RESULT eventid="1062" points="468" swimtime="00:00:30.56" resultid="10126" heatid="13902" lane="9" entrytime="00:00:29.80" entrycourse="LCM" />
                <RESULT eventid="1187" points="356" reactiontime="+82" swimtime="00:00:38.17" resultid="10127" heatid="13948" lane="8" entrytime="00:00:35.10" entrycourse="LCM" />
                <RESULT eventid="1256" points="450" reactiontime="+85" swimtime="00:01:07.94" resultid="10128" heatid="13976" lane="1" entrytime="00:01:06.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="336" reactiontime="+85" swimtime="00:01:32.50" resultid="10129" heatid="14004" lane="7" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="10130" heatid="14042" lane="5" entrytime="00:02:35.00" entrycourse="LCM" />
                <RESULT eventid="1664" points="325" reactiontime="+81" swimtime="00:00:42.84" resultid="10131" heatid="14087" lane="2" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-21" firstname="Michał" gender="M" lastname="Krysiak" nation="POL" athleteid="10105">
              <RESULTS>
                <RESULT eventid="1079" points="443" reactiontime="+80" swimtime="00:00:27.42" resultid="10106" heatid="13914" lane="2" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="323" reactiontime="+87" swimtime="00:02:46.14" resultid="10107" heatid="13928" lane="0" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:08.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="442" reactiontime="+81" swimtime="00:01:01.54" resultid="10108" heatid="13987" lane="0" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="334" reactiontime="+80" swimtime="00:02:40.66" resultid="10109" heatid="13995" lane="7" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:02:00.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="436" reactiontime="+87" swimtime="00:00:29.57" resultid="10110" heatid="14026" lane="0" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1508" points="320" reactiontime="+85" swimtime="00:02:29.12" resultid="10111" heatid="14049" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="451" reactiontime="+80" swimtime="00:01:04.93" resultid="10112" heatid="14070" lane="5" entrytime="00:01:06.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="321" reactiontime="+89" swimtime="00:05:21.08" resultid="10113" heatid="14112" lane="0" entrytime="00:05:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                    <SPLIT distance="150" swimtime="00:01:56.17" />
                    <SPLIT distance="200" swimtime="00:02:37.68" />
                    <SPLIT distance="250" swimtime="00:03:18.89" />
                    <SPLIT distance="300" swimtime="00:04:01.17" />
                    <SPLIT distance="350" swimtime="00:04:42.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-21" firstname="Wiktoria" gender="F" lastname="Podkowińska" nation="POL" athleteid="10138">
              <RESULTS>
                <RESULT eventid="1096" points="392" swimtime="00:02:52.32" resultid="10139" heatid="13921" lane="9" entrytime="00:02:56.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="464" reactiontime="+74" swimtime="00:01:07.25" resultid="10140" heatid="13976" lane="0" entrytime="00:01:07.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="371" swimtime="00:00:33.97" resultid="10141" heatid="14017" lane="9" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1555" points="397" reactiontime="+76" swimtime="00:06:05.05" resultid="10142" heatid="14058" lane="6" entrytime="00:06:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="150" swimtime="00:02:14.21" />
                    <SPLIT distance="200" swimtime="00:03:02.70" />
                    <SPLIT distance="250" swimtime="00:03:54.32" />
                    <SPLIT distance="300" swimtime="00:04:45.95" />
                    <SPLIT distance="350" swimtime="00:05:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="337" reactiontime="+83" swimtime="00:01:19.91" resultid="10143" heatid="14065" lane="1" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="316" reactiontime="+81" swimtime="00:00:43.28" resultid="10144" heatid="14086" lane="0" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="398" reactiontime="+47" swimtime="00:02:06.98" resultid="10162" heatid="13998" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="150" swimtime="00:01:36.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10145" number="1" reactiontime="+47" />
                    <RELAYPOSITION athleteid="10119" number="2" />
                    <RELAYPOSITION athleteid="10105" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="10114" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="444" reactiontime="+75" swimtime="00:01:51.18" resultid="10163" heatid="14056" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:00:58.11" />
                    <SPLIT distance="150" swimtime="00:01:25.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10114" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="10105" number="2" />
                    <RELAYPOSITION athleteid="10119" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10145" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="10160" heatid="13996" lane="4" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10132" number="1" />
                    <RELAYPOSITION athleteid="10125" number="2" />
                    <RELAYPOSITION athleteid="10138" number="3" />
                    <RELAYPOSITION athleteid="10152" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="10161" heatid="14054" lane="4" entrytime="00:02:02.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10132" number="1" />
                    <RELAYPOSITION athleteid="10152" number="2" />
                    <RELAYPOSITION athleteid="10138" number="3" />
                    <RELAYPOSITION athleteid="10125" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1130" points="362" reactiontime="+80" swimtime="00:01:59.00" resultid="10158" heatid="13934" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="100" swimtime="00:01:01.08" />
                    <SPLIT distance="150" swimtime="00:01:31.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10105" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="10152" number="2" />
                    <RELAYPOSITION athleteid="10125" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="10119" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="309" reactiontime="+52" swimtime="00:02:18.15" resultid="10159" heatid="14101" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:44.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10145" number="1" reactiontime="+52" />
                    <RELAYPOSITION athleteid="10119" number="2" />
                    <RELAYPOSITION athleteid="10138" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="10152" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9925" name="Szczecineckie Towarzystwo Pływackie MASTERS" shortname="Szczecineckie Towarzystwo Pływ">
          <CONTACT name="a" />
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10997" name="T.P. Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="11023">
              <RESULTS>
                <RESULT eventid="1079" points="493" reactiontime="+74" swimtime="00:00:26.46" resultid="11024" heatid="13916" lane="6" entrytime="00:00:25.99" />
                <RESULT eventid="1113" points="506" reactiontime="+90" swimtime="00:02:22.98" resultid="11025" heatid="13929" lane="0" entrytime="00:02:40.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:07.99" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="473" reactiontime="+76" swimtime="00:05:12.93" resultid="11026" heatid="14061" lane="4" entrytime="00:05:50.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                    <SPLIT distance="250" swimtime="00:03:13.95" />
                    <SPLIT distance="350" swimtime="00:04:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11027" heatid="14081" lane="7" entrytime="00:02:36.70" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="11028" heatid="14112" lane="1" entrytime="00:05:10.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="11016">
              <RESULTS>
                <RESULT eventid="1079" points="146" swimtime="00:00:39.68" resultid="11017" heatid="13906" lane="9" entrytime="00:00:39.50" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="11018" heatid="13950" lane="7" entrytime="00:00:57.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="11019" heatid="13979" lane="9" entrytime="00:01:39.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="11020" heatid="14033" lane="7" entrytime="00:02:05.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11021" heatid="14077" lane="5" entrytime="00:04:20.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="11022" heatid="14089" lane="3" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="11011">
              <RESULTS>
                <RESULT eventid="1079" points="419" swimtime="00:00:27.94" resultid="11012" heatid="13910" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1113" points="379" reactiontime="+87" swimtime="00:02:37.46" resultid="11013" heatid="13928" lane="4" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="406" reactiontime="+61" swimtime="00:00:32.44" resultid="11014" heatid="13957" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1273" points="434" reactiontime="+85" swimtime="00:01:01.94" resultid="11015" heatid="13985" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="11005">
              <RESULTS>
                <RESULT eventid="1079" points="283" reactiontime="+95" swimtime="00:00:31.82" resultid="11006" heatid="13909" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1113" points="184" reactiontime="+95" swimtime="00:03:20.37" resultid="11007" heatid="13924" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:37.22" />
                    <SPLIT distance="150" swimtime="00:02:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="261" swimtime="00:01:13.35" resultid="11008" heatid="13982" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="224" reactiontime="+93" swimtime="00:00:36.92" resultid="11009" heatid="14021" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1613" points="159" reactiontime="+101" swimtime="00:01:31.88" resultid="11010" heatid="14067" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="11029">
              <RESULTS>
                <RESULT eventid="1239" points="202" reactiontime="+98" swimtime="00:03:36.42" resultid="11030" heatid="13966" lane="6" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:41.64" />
                    <SPLIT distance="150" swimtime="00:02:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="217" swimtime="00:01:36.37" resultid="11031" heatid="14008" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="261" swimtime="00:00:41.32" resultid="11032" heatid="14092" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5130" nation="GER" region="17" clubid="9389" name="TG Lage">
          <CONTACT city="Lage" email="tg-schwimmen@gmx.de" name="Lange Ute" state="NO" street="Ringstrasse 3" zip="32791" />
          <ATHLETES>
            <ATHLETE birthdate="1968-04-07" firstname="Konstantin" gender="M" lastname="Sklyar" nation="GER" license="321129" athleteid="9390">
              <RESULTS>
                <RESULT eventid="1165" points="310" reactiontime="+98" swimtime="00:21:26.57" resultid="9391" heatid="13942" lane="4" entrytime="00:20:49.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:01:59.52" />
                    <SPLIT distance="200" swimtime="00:02:41.96" />
                    <SPLIT distance="250" swimtime="00:03:25.13" />
                    <SPLIT distance="300" swimtime="00:04:07.68" />
                    <SPLIT distance="350" swimtime="00:04:51.13" />
                    <SPLIT distance="400" swimtime="00:05:34.53" />
                    <SPLIT distance="450" swimtime="00:06:18.56" />
                    <SPLIT distance="500" swimtime="00:07:02.51" />
                    <SPLIT distance="550" swimtime="00:07:46.56" />
                    <SPLIT distance="600" swimtime="00:08:30.51" />
                    <SPLIT distance="650" swimtime="00:09:14.96" />
                    <SPLIT distance="700" swimtime="00:09:59.36" />
                    <SPLIT distance="750" swimtime="00:10:43.15" />
                    <SPLIT distance="800" swimtime="00:11:26.27" />
                    <SPLIT distance="850" swimtime="00:12:09.41" />
                    <SPLIT distance="900" swimtime="00:12:52.34" />
                    <SPLIT distance="950" swimtime="00:13:35.54" />
                    <SPLIT distance="1000" swimtime="00:14:18.85" />
                    <SPLIT distance="1050" swimtime="00:15:02.03" />
                    <SPLIT distance="1100" swimtime="00:15:45.68" />
                    <SPLIT distance="1150" swimtime="00:16:28.89" />
                    <SPLIT distance="1200" swimtime="00:17:12.62" />
                    <SPLIT distance="1250" swimtime="00:17:55.13" />
                    <SPLIT distance="1300" swimtime="00:18:38.86" />
                    <SPLIT distance="1350" swimtime="00:19:21.98" />
                    <SPLIT distance="1400" swimtime="00:20:03.54" />
                    <SPLIT distance="1450" swimtime="00:20:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="299" reactiontime="+90" swimtime="00:03:09.88" resultid="9392" heatid="13968" lane="3" entrytime="00:02:59.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                    <SPLIT distance="100" swimtime="00:01:31.14" />
                    <SPLIT distance="150" swimtime="00:02:21.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="231" reactiontime="+94" swimtime="00:03:01.50" resultid="9393" heatid="13995" lane="8" entrytime="00:02:49.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="271" reactiontime="+93" swimtime="00:01:29.42" resultid="9394" heatid="14010" lane="2" entrytime="00:01:21.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="290" reactiontime="+95" swimtime="00:06:08.14" resultid="9395" heatid="14061" lane="6" entrytime="00:05:58.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:21.69" />
                    <SPLIT distance="150" swimtime="00:03:55.69" />
                    <SPLIT distance="200" swimtime="00:03:01.97" />
                    <SPLIT distance="300" swimtime="00:04:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="303" reactiontime="+89" swimtime="00:01:14.11" resultid="9396" heatid="14070" lane="8" entrytime="00:01:12.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="9990" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="10007">
              <RESULTS>
                <RESULT eventid="1079" points="96" reactiontime="+94" swimtime="00:00:45.58" resultid="10008" heatid="13905" lane="8" entrytime="00:00:42.23" />
                <RESULT eventid="1205" points="98" reactiontime="+73" swimtime="00:00:51.97" resultid="10009" heatid="13951" lane="0" entrytime="00:00:51.09" />
                <RESULT eventid="1239" points="95" reactiontime="+112" swimtime="00:04:37.61" resultid="10010" heatid="13964" lane="3" entrytime="00:04:24.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.76" />
                    <SPLIT distance="100" swimtime="00:02:12.89" />
                    <SPLIT distance="150" swimtime="00:03:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="97" reactiontime="+122" swimtime="00:02:05.87" resultid="10011" heatid="14006" lane="1" entrytime="00:01:59.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="71" reactiontime="+70" swimtime="00:02:05.36" resultid="10012" heatid="14033" lane="8" entrytime="00:02:05.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="128" reactiontime="+114" swimtime="00:00:52.38" resultid="10013" heatid="14090" lane="5" entrytime="00:00:49.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="10037">
              <RESULTS>
                <RESULT eventid="1079" points="313" reactiontime="+81" swimtime="00:00:30.79" resultid="10038" heatid="13908" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1341" points="183" reactiontime="+94" swimtime="00:03:16.15" resultid="10039" heatid="13994" lane="7" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:31.42" />
                    <SPLIT distance="150" swimtime="00:02:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="206" reactiontime="+96" swimtime="00:02:52.52" resultid="10040" heatid="14048" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:02:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="212" reactiontime="+94" swimtime="00:06:48.90" resultid="10041" heatid="14060" lane="4" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="150" swimtime="00:02:27.60" />
                    <SPLIT distance="250" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:06:05.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="256" reactiontime="+89" swimtime="00:01:18.42" resultid="10042" heatid="14069" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="10043" heatid="14110" lane="3" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="10014">
              <RESULTS>
                <RESULT eventid="1079" points="262" reactiontime="+82" swimtime="00:00:32.67" resultid="10015" heatid="13909" lane="8" entrytime="00:00:31.80" />
                <RESULT eventid="1165" points="188" reactiontime="+80" swimtime="00:25:18.07" resultid="10016" heatid="13940" lane="5" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:34.37" />
                    <SPLIT distance="150" swimtime="00:02:26.56" />
                    <SPLIT distance="200" swimtime="00:03:17.69" />
                    <SPLIT distance="250" swimtime="00:04:08.46" />
                    <SPLIT distance="300" swimtime="00:04:59.03" />
                    <SPLIT distance="350" swimtime="00:05:49.84" />
                    <SPLIT distance="400" swimtime="00:06:41.36" />
                    <SPLIT distance="450" swimtime="00:07:32.63" />
                    <SPLIT distance="500" swimtime="00:08:23.79" />
                    <SPLIT distance="550" swimtime="00:09:15.45" />
                    <SPLIT distance="600" swimtime="00:10:07.06" />
                    <SPLIT distance="650" swimtime="00:10:58.21" />
                    <SPLIT distance="700" swimtime="00:11:49.89" />
                    <SPLIT distance="750" swimtime="00:12:41.47" />
                    <SPLIT distance="800" swimtime="00:13:33.18" />
                    <SPLIT distance="850" swimtime="00:14:24.68" />
                    <SPLIT distance="900" swimtime="00:15:15.10" />
                    <SPLIT distance="950" swimtime="00:16:07.71" />
                    <SPLIT distance="1000" swimtime="00:16:57.21" />
                    <SPLIT distance="1050" swimtime="00:17:48.88" />
                    <SPLIT distance="1100" swimtime="00:18:39.35" />
                    <SPLIT distance="1150" swimtime="00:19:30.52" />
                    <SPLIT distance="1200" swimtime="00:20:21.55" />
                    <SPLIT distance="1250" swimtime="00:21:11.33" />
                    <SPLIT distance="1300" swimtime="00:22:03.18" />
                    <SPLIT distance="1350" swimtime="00:22:54.92" />
                    <SPLIT distance="1400" swimtime="00:23:45.57" />
                    <SPLIT distance="1450" swimtime="00:24:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="253" reactiontime="+82" swimtime="00:01:14.15" resultid="10017" heatid="13981" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="201" swimtime="00:00:38.23" resultid="10018" heatid="14021" lane="9" entrytime="00:00:35.50" />
                <RESULT eventid="1508" points="205" reactiontime="+88" swimtime="00:02:52.96" resultid="10019" heatid="14048" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:02:13.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="10020" heatid="14068" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1744" points="197" reactiontime="+81" swimtime="00:06:17.84" resultid="10021" heatid="14109" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:02:14.76" />
                    <SPLIT distance="200" swimtime="00:03:03.77" />
                    <SPLIT distance="250" swimtime="00:03:52.79" />
                    <SPLIT distance="300" swimtime="00:04:43.10" />
                    <SPLIT distance="350" swimtime="00:05:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="10029">
              <RESULTS>
                <RESULT eventid="1079" points="446" reactiontime="+83" swimtime="00:00:27.35" resultid="10030" heatid="13913" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1239" points="429" reactiontime="+87" swimtime="00:02:48.39" resultid="10031" heatid="13969" lane="2" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:01:21.23" />
                    <SPLIT distance="150" swimtime="00:02:05.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="10032" heatid="13986" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1406" points="507" reactiontime="+83" swimtime="00:01:12.61" resultid="10033" heatid="14012" lane="5" entrytime="00:01:15.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="416" reactiontime="+94" swimtime="00:02:16.58" resultid="10034" heatid="14051" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="546" reactiontime="+82" swimtime="00:00:32.32" resultid="10035" heatid="14097" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="10036" heatid="14113" lane="8" entrytime="00:04:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="9996">
              <RESULTS>
                <RESULT eventid="1079" points="38" reactiontime="+142" swimtime="00:01:01.84" resultid="9997" heatid="13904" lane="0" entrytime="00:01:03.40" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="9998" heatid="14089" lane="1" entrytime="00:01:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="10022">
              <RESULTS>
                <RESULT eventid="1096" points="440" reactiontime="+78" swimtime="00:02:45.73" resultid="10023" heatid="13921" lane="6" entrytime="00:02:44.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="418" reactiontime="+79" swimtime="00:03:05.92" resultid="10024" heatid="13962" lane="6" entrytime="00:03:05.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                    <SPLIT distance="150" swimtime="00:02:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="429" reactiontime="+88" swimtime="00:01:25.31" resultid="10025" heatid="14004" lane="1" entrytime="00:01:25.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1555" points="429" reactiontime="+81" swimtime="00:05:55.64" resultid="10026" heatid="14058" lane="5" entrytime="00:06:01.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:08.02" />
                    <SPLIT distance="200" swimtime="00:02:53.61" />
                    <SPLIT distance="250" swimtime="00:03:42.69" />
                    <SPLIT distance="300" swimtime="00:04:32.60" />
                    <SPLIT distance="350" swimtime="00:05:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="357" reactiontime="+78" swimtime="00:01:18.36" resultid="10027" heatid="14063" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="407" reactiontime="+74" swimtime="00:00:39.75" resultid="10028" heatid="14086" lane="5" entrytime="00:00:39.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="10049">
              <RESULTS>
                <RESULT eventid="1113" points="111" reactiontime="+109" swimtime="00:03:56.53" resultid="10050" heatid="13923" lane="2" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                    <SPLIT distance="100" swimtime="00:01:53.74" />
                    <SPLIT distance="150" swimtime="00:02:57.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="91" reactiontime="+97" swimtime="00:00:53.28" resultid="10051" heatid="13951" lane="8" entrytime="00:00:51.00" />
                <RESULT eventid="1406" points="122" reactiontime="+109" swimtime="00:01:56.47" resultid="10052" heatid="14006" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="114" swimtime="00:00:46.20" resultid="10053" heatid="14019" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1681" points="148" reactiontime="+109" swimtime="00:00:49.91" resultid="10054" heatid="14090" lane="4" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="9991">
              <RESULTS>
                <RESULT eventid="1079" points="89" reactiontime="+107" swimtime="00:00:46.68" resultid="9992" heatid="13905" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="9993" heatid="13978" lane="1" entrytime="00:01:46.20" />
                <RESULT eventid="1474" points="41" swimtime="00:02:30.14" resultid="9994" heatid="14032" lane="4" entrytime="00:02:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="9995" heatid="14077" lane="9" entrytime="00:05:08.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="9999">
              <RESULTS>
                <RESULT eventid="1113" points="52" reactiontime="+150" swimtime="00:05:04.00" resultid="10000" heatid="13923" lane="0" entrytime="00:04:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.14" />
                    <SPLIT distance="100" swimtime="00:02:36.26" />
                    <SPLIT distance="150" swimtime="00:04:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="57" reactiontime="+151" swimtime="00:05:29.56" resultid="10001" heatid="13964" lane="6" entrytime="00:04:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.93" />
                    <SPLIT distance="100" swimtime="00:02:42.82" />
                    <SPLIT distance="150" swimtime="00:04:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="33" reactiontime="+151" swimtime="00:05:46.93" resultid="10002" heatid="13992" lane="2" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.03" />
                    <SPLIT distance="100" swimtime="00:02:31.66" />
                    <SPLIT distance="150" swimtime="00:04:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="75" reactiontime="+142" swimtime="00:04:00.88" resultid="10003" heatid="14045" lane="3" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.35" />
                    <SPLIT distance="150" swimtime="00:03:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="55" reactiontime="+152" swimtime="00:10:38.38" resultid="10004" heatid="14059" lane="2" entrytime="00:10:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.13" />
                    <SPLIT distance="100" swimtime="00:02:37.06" />
                    <SPLIT distance="150" swimtime="00:04:06.80" />
                    <SPLIT distance="200" swimtime="00:05:38.55" />
                    <SPLIT distance="250" swimtime="00:07:05.59" />
                    <SPLIT distance="300" swimtime="00:08:36.59" />
                    <SPLIT distance="350" swimtime="00:09:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="33" reactiontime="+128" swimtime="00:02:34.54" resultid="10005" heatid="14066" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="36" reactiontime="+98" swimtime="00:05:38.76" resultid="10006" heatid="14077" lane="1" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.24" />
                    <SPLIT distance="100" swimtime="00:02:49.35" />
                    <SPLIT distance="150" swimtime="00:04:16.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="46" reactiontime="+82" swimtime="00:04:19.13" resultid="10062" heatid="13997" lane="3" entrytime="00:03:43.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.44" />
                    <SPLIT distance="100" swimtime="00:02:27.61" />
                    <SPLIT distance="150" swimtime="00:03:33.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10007" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="9996" number="2" />
                    <RELAYPOSITION athleteid="9999" number="3" reactiontime="+126" />
                    <RELAYPOSITION athleteid="9991" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="76" reactiontime="+130" swimtime="00:03:19.73" resultid="10063" heatid="14055" lane="1" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:45.02" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9999" number="1" reactiontime="+130" />
                    <RELAYPOSITION athleteid="9996" number="2" />
                    <RELAYPOSITION athleteid="10007" number="3" reactiontime="+117" />
                    <RELAYPOSITION athleteid="9991" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="12121" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="12145">
              <RESULTS>
                <RESULT eventid="1113" points="214" swimtime="00:03:10.41" resultid="12146" heatid="13925" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:29.48" />
                    <SPLIT distance="150" swimtime="00:02:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="240" reactiontime="+105" swimtime="00:03:24.15" resultid="12147" heatid="13966" lane="7" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:37.34" />
                    <SPLIT distance="150" swimtime="00:02:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="108" reactiontime="+88" swimtime="00:03:53.51" resultid="12148" heatid="13993" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:47.48" />
                    <SPLIT distance="150" swimtime="00:02:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="234" reactiontime="+90" swimtime="00:01:33.94" resultid="12149" heatid="14007" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="232" reactiontime="+100" swimtime="00:00:36.49" resultid="12150" heatid="14020" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1613" points="158" reactiontime="+87" swimtime="00:01:32.12" resultid="12151" heatid="14067" lane="2" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="283" reactiontime="+90" swimtime="00:00:40.21" resultid="12152" heatid="14092" lane="1" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="12131">
              <RESULTS>
                <RESULT eventid="1079" points="164" reactiontime="+120" swimtime="00:00:38.14" resultid="12132" heatid="13906" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1205" points="154" reactiontime="+85" swimtime="00:00:44.79" resultid="12133" heatid="13952" lane="8" entrytime="00:00:42.50" />
                <RESULT eventid="1474" points="111" reactiontime="+91" swimtime="00:01:47.78" resultid="12134" heatid="14034" lane="0" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="100" reactiontime="+87" swimtime="00:04:00.71" resultid="12135" heatid="14078" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.20" />
                    <SPLIT distance="100" swimtime="00:02:04.50" />
                    <SPLIT distance="150" swimtime="00:03:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="12136" heatid="14107" lane="4" entrytime="00:07:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="12137">
              <RESULTS>
                <RESULT eventid="1113" points="205" swimtime="00:03:13.21" resultid="12138" heatid="13926" lane="9" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                    <SPLIT distance="150" swimtime="00:02:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="178" reactiontime="+77" swimtime="00:00:42.67" resultid="12139" heatid="13952" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="12140" heatid="13993" lane="6" entrytime="00:03:40.00" />
                <RESULT eventid="1474" points="192" reactiontime="+75" swimtime="00:01:29.91" resultid="12141" heatid="14034" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="206" reactiontime="+92" swimtime="00:06:52.22" resultid="12142" heatid="14060" lane="5" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                    <SPLIT distance="100" swimtime="00:01:47.72" />
                    <SPLIT distance="150" swimtime="00:02:38.28" />
                    <SPLIT distance="200" swimtime="00:03:28.01" />
                    <SPLIT distance="250" swimtime="00:04:23.80" />
                    <SPLIT distance="300" swimtime="00:05:20.19" />
                    <SPLIT distance="350" swimtime="00:06:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="200" reactiontime="+80" swimtime="00:03:11.19" resultid="12143" heatid="14079" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                    <SPLIT distance="100" swimtime="00:01:34.91" />
                    <SPLIT distance="150" swimtime="00:02:23.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="12144" heatid="14109" lane="8" entrytime="00:06:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="12153">
              <RESULTS>
                <RESULT eventid="1113" points="270" reactiontime="+81" swimtime="00:02:56.28" resultid="12154" heatid="13926" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="258" reactiontime="+81" swimtime="00:03:19.46" resultid="12155" heatid="13967" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:34.49" />
                    <SPLIT distance="150" swimtime="00:02:18.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="331" reactiontime="+77" swimtime="00:01:23.70" resultid="12156" heatid="14009" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="270" swimtime="00:02:37.71" resultid="12157" heatid="14050" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="232" reactiontime="+85" swimtime="00:01:21.05" resultid="12158" heatid="14069" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="352" reactiontime="+81" swimtime="00:00:37.40" resultid="12159" heatid="14094" lane="4" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="12122">
              <RESULTS>
                <RESULT eventid="1062" points="225" reactiontime="+96" swimtime="00:00:39.01" resultid="12123" heatid="13898" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1096" points="147" reactiontime="+100" swimtime="00:03:58.83" resultid="12124" heatid="13919" lane="8" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.13" />
                    <SPLIT distance="100" swimtime="00:02:01.72" />
                    <SPLIT distance="150" swimtime="00:03:08.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="142" swimtime="00:00:51.78" resultid="12125" heatid="13945" lane="1" entrytime="00:00:52.00" />
                <RESULT eventid="1256" points="168" reactiontime="+102" swimtime="00:01:34.19" resultid="12126" heatid="13971" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="100" reactiontime="+96" swimtime="00:00:52.53" resultid="12127" heatid="14015" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1555" points="141" reactiontime="+117" swimtime="00:08:35.03" resultid="12128" heatid="14057" lane="6" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.78" />
                    <SPLIT distance="100" swimtime="00:02:09.99" />
                    <SPLIT distance="150" swimtime="00:03:20.51" />
                    <SPLIT distance="200" swimtime="00:04:26.00" />
                    <SPLIT distance="250" swimtime="00:05:37.11" />
                    <SPLIT distance="300" swimtime="00:06:47.80" />
                    <SPLIT distance="350" swimtime="00:07:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="95" reactiontime="+106" swimtime="00:02:01.75" resultid="12129" heatid="14063" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="148" reactiontime="+103" swimtime="00:00:55.71" resultid="12130" heatid="14083" lane="4" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="216" reactiontime="+100" swimtime="00:02:35.64" resultid="12160" heatid="13998" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:02:01.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12131" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="12145" number="2" />
                    <RELAYPOSITION athleteid="12153" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="12137" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UKSCI" nation="POL" region="WIE" clubid="10098" name="UKS CITYZEN Poznań">
          <CONTACT name="roszak" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="10099">
              <RESULTS>
                <RESULT eventid="1147" points="258" reactiontime="+98" swimtime="00:12:45.15" resultid="10100" heatid="13936" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:16.26" />
                    <SPLIT distance="200" swimtime="00:03:05.25" />
                    <SPLIT distance="250" swimtime="00:03:54.29" />
                    <SPLIT distance="300" swimtime="00:04:43.08" />
                    <SPLIT distance="350" swimtime="00:05:31.95" />
                    <SPLIT distance="400" swimtime="00:06:20.72" />
                    <SPLIT distance="450" swimtime="00:07:09.06" />
                    <SPLIT distance="500" swimtime="00:07:57.66" />
                    <SPLIT distance="550" swimtime="00:08:46.39" />
                    <SPLIT distance="600" swimtime="00:09:35.39" />
                    <SPLIT distance="650" swimtime="00:10:23.61" />
                    <SPLIT distance="700" swimtime="00:11:12.32" />
                    <SPLIT distance="750" swimtime="00:11:59.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="282" reactiontime="+82" swimtime="00:01:19.40" resultid="10101" heatid="13973" lane="4" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="261" reactiontime="+88" swimtime="00:02:56.68" resultid="10102" heatid="14041" lane="8" entrytime="00:02:53.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                    <SPLIT distance="150" swimtime="00:02:11.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="253" reactiontime="+100" swimtime="00:06:16.49" resultid="10103" heatid="14103" lane="4" entrytime="00:06:09.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                    <SPLIT distance="100" swimtime="00:01:28.20" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                    <SPLIT distance="200" swimtime="00:03:05.37" />
                    <SPLIT distance="250" swimtime="00:03:53.70" />
                    <SPLIT distance="300" swimtime="00:04:42.30" />
                    <SPLIT distance="350" swimtime="00:05:30.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="11826" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="11846">
              <RESULTS>
                <RESULT eventid="1079" points="466" swimtime="00:00:26.96" resultid="11847" heatid="13913" lane="9" entrytime="00:00:28.04" />
                <RESULT eventid="1113" points="410" reactiontime="+88" swimtime="00:02:33.34" resultid="11848" heatid="13928" lane="6" entrytime="00:02:44.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="363" reactiontime="+73" swimtime="00:00:33.68" resultid="11849" heatid="13954" lane="3" entrytime="00:00:36.24" />
                <RESULT eventid="1273" points="490" reactiontime="+85" swimtime="00:00:59.50" resultid="11850" heatid="13986" lane="1" entrytime="00:01:01.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="460" reactiontime="+86" swimtime="00:00:29.05" resultid="11851" heatid="14024" lane="2" entrytime="00:00:31.24" />
                <RESULT eventid="1508" points="431" reactiontime="+91" swimtime="00:02:15.02" resultid="11852" heatid="14051" lane="3" entrytime="00:02:15.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="404" reactiontime="+91" swimtime="00:01:07.35" resultid="11853" heatid="14070" lane="0" entrytime="00:01:14.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="461" reactiontime="+85" swimtime="00:00:34.18" resultid="11854" heatid="14095" lane="2" entrytime="00:00:36.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="11864">
              <RESULTS>
                <RESULT eventid="1079" points="371" reactiontime="+84" swimtime="00:00:29.09" resultid="11865" heatid="13911" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1205" points="319" reactiontime="+63" swimtime="00:00:35.18" resultid="11866" heatid="13955" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="411" reactiontime="+79" swimtime="00:01:03.05" resultid="11867" heatid="13984" lane="7" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="320" reactiontime="+88" swimtime="00:00:32.77" resultid="11868" heatid="14023" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1508" points="347" reactiontime="+82" swimtime="00:02:25.02" resultid="11869" heatid="14050" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="150" swimtime="00:01:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="260" reactiontime="+89" swimtime="00:01:18.01" resultid="11870" heatid="14069" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-03" firstname="Patrycja" gender="F" lastname="Urbaniak" nation="POL" athleteid="11842">
              <RESULTS>
                <RESULT eventid="1324" points="221" reactiontime="+94" swimtime="00:03:21.27" resultid="11843" heatid="13991" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:33.43" />
                    <SPLIT distance="150" swimtime="00:02:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="11844" heatid="14043" lane="0" entrytime="00:02:30.00" />
                <RESULT eventid="1595" points="284" reactiontime="+82" swimtime="00:01:24.56" resultid="11845" heatid="14065" lane="7" entrytime="00:01:18.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="11827">
              <RESULTS>
                <RESULT eventid="1147" points="366" reactiontime="+87" swimtime="00:11:21.31" resultid="11828" heatid="13937" lane="7" entrytime="00:11:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:00.84" />
                    <SPLIT distance="200" swimtime="00:02:44.06" />
                    <SPLIT distance="250" swimtime="00:03:27.08" />
                    <SPLIT distance="300" swimtime="00:04:10.47" />
                    <SPLIT distance="350" swimtime="00:04:53.86" />
                    <SPLIT distance="400" swimtime="00:05:37.39" />
                    <SPLIT distance="450" swimtime="00:06:20.53" />
                    <SPLIT distance="500" swimtime="00:07:03.93" />
                    <SPLIT distance="550" swimtime="00:07:47.36" />
                    <SPLIT distance="600" swimtime="00:08:31.08" />
                    <SPLIT distance="650" swimtime="00:09:14.43" />
                    <SPLIT distance="700" swimtime="00:09:58.13" />
                    <SPLIT distance="750" swimtime="00:10:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="320" reactiontime="+76" swimtime="00:00:39.53" resultid="11829" heatid="13946" lane="3" entrytime="00:00:39.90" />
                <RESULT eventid="1222" points="313" reactiontime="+92" swimtime="00:03:24.79" resultid="11830" heatid="13961" lane="4" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="337" reactiontime="+75" swimtime="00:01:23.48" resultid="11831" heatid="14030" lane="5" entrytime="00:01:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="348" swimtime="00:02:40.51" resultid="11832" heatid="14042" lane="6" entrytime="00:02:40.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="355" reactiontime="+80" swimtime="00:02:55.07" resultid="11833" heatid="14075" lane="8" entrytime="00:02:58.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:11.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="344" reactiontime="+90" swimtime="00:05:40.04" resultid="11834" heatid="14105" lane="0" entrytime="00:05:28.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:05.70" />
                    <SPLIT distance="200" swimtime="00:02:49.24" />
                    <SPLIT distance="250" swimtime="00:03:32.89" />
                    <SPLIT distance="300" swimtime="00:04:16.24" />
                    <SPLIT distance="350" swimtime="00:04:59.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Witold" gender="M" lastname="Flak" nation="POL" athleteid="11899">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:32)" eventid="1079" reactiontime="+66" status="DSQ" swimtime="00:00:29.60" resultid="11900" heatid="13913" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1205" points="270" reactiontime="+67" swimtime="00:00:37.19" resultid="11901" heatid="13954" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1406" points="319" reactiontime="+88" swimtime="00:01:24.75" resultid="11902" heatid="14012" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="379" reactiontime="+103" swimtime="00:00:36.49" resultid="11903" heatid="14095" lane="1" entrytime="00:00:36.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-15" firstname="Paweł" gender="M" lastname="Nowak" nation="POL" athleteid="11882">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="11883" heatid="13979" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1440" points="271" swimtime="00:00:34.66" resultid="11884" heatid="14021" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-04-09" firstname="Zbigniew" gender="M" lastname="Ramos" nation="POL" athleteid="11871">
              <RESULTS>
                <RESULT eventid="1440" points="273" reactiontime="+97" swimtime="00:00:34.56" resultid="11872" heatid="14021" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="11873" heatid="14093" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="11835">
              <RESULTS>
                <RESULT eventid="1062" points="386" reactiontime="+88" swimtime="00:00:32.57" resultid="11836" heatid="13901" lane="0" entrytime="00:00:32.05" />
                <RESULT eventid="1187" points="303" reactiontime="+72" swimtime="00:00:40.27" resultid="11837" heatid="13946" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1256" points="376" reactiontime="+87" swimtime="00:01:12.13" resultid="11838" heatid="13975" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="278" reactiontime="+96" swimtime="00:00:37.39" resultid="11839" heatid="14016" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1491" points="288" reactiontime="+104" swimtime="00:02:50.97" resultid="11840" heatid="14042" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:07.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="244" reactiontime="+96" swimtime="00:01:28.92" resultid="11841" heatid="14064" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="11874">
              <RESULTS>
                <RESULT eventid="1079" points="296" reactiontime="+76" swimtime="00:00:31.36" resultid="11875" heatid="13910" lane="8" entrytime="00:00:30.88" />
                <RESULT comment="(Time: 20:38), Przekroczony regulaminowy limit czasu." eventid="1165" reactiontime="+87" status="OTL" swimtime="00:23:17.69" resultid="11876" heatid="13941" lane="4" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                    <SPLIT distance="200" swimtime="00:02:49.64" />
                    <SPLIT distance="250" swimtime="00:03:34.20" />
                    <SPLIT distance="300" swimtime="00:04:19.12" />
                    <SPLIT distance="350" swimtime="00:05:04.21" />
                    <SPLIT distance="400" swimtime="00:05:49.53" />
                    <SPLIT distance="450" swimtime="00:06:35.72" />
                    <SPLIT distance="500" swimtime="00:07:21.70" />
                    <SPLIT distance="550" swimtime="00:08:07.96" />
                    <SPLIT distance="600" swimtime="00:08:54.90" />
                    <SPLIT distance="650" swimtime="00:09:41.34" />
                    <SPLIT distance="700" swimtime="00:10:28.20" />
                    <SPLIT distance="750" swimtime="00:11:15.36" />
                    <SPLIT distance="800" swimtime="00:12:03.33" />
                    <SPLIT distance="850" swimtime="00:12:51.41" />
                    <SPLIT distance="900" swimtime="00:13:39.91" />
                    <SPLIT distance="950" swimtime="00:14:27.90" />
                    <SPLIT distance="1000" swimtime="00:15:16.70" />
                    <SPLIT distance="1050" swimtime="00:16:05.64" />
                    <SPLIT distance="1100" swimtime="00:16:53.96" />
                    <SPLIT distance="1150" swimtime="00:17:42.59" />
                    <SPLIT distance="1200" swimtime="00:18:31.95" />
                    <SPLIT distance="1250" swimtime="00:19:21.23" />
                    <SPLIT distance="1300" swimtime="00:20:09.93" />
                    <SPLIT distance="1350" swimtime="00:20:59.47" />
                    <SPLIT distance="1400" swimtime="00:21:47.76" />
                    <SPLIT distance="1450" swimtime="00:22:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="305" reactiontime="+74" swimtime="00:01:09.67" resultid="11877" heatid="13982" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="11878" heatid="13993" lane="1" entrytime="00:03:45.00" />
                <RESULT eventid="1508" points="267" reactiontime="+80" swimtime="00:02:38.21" resultid="11879" heatid="14048" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:58.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="225" swimtime="00:06:40.90" resultid="11880" heatid="14061" lane="9" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:29.08" />
                    <SPLIT distance="150" swimtime="00:02:24.41" />
                    <SPLIT distance="200" swimtime="00:03:18.24" />
                    <SPLIT distance="250" swimtime="00:04:16.58" />
                    <SPLIT distance="300" swimtime="00:05:15.11" />
                    <SPLIT distance="350" swimtime="00:05:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="272" reactiontime="+85" swimtime="00:05:39.40" resultid="11881" heatid="14111" lane="1" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                    <SPLIT distance="200" swimtime="00:02:44.66" />
                    <SPLIT distance="250" swimtime="00:03:29.13" />
                    <SPLIT distance="300" swimtime="00:04:14.52" />
                    <SPLIT distance="350" swimtime="00:04:58.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="11855">
              <RESULTS>
                <RESULT eventid="1079" points="346" reactiontime="+78" swimtime="00:00:29.76" resultid="11856" heatid="13907" lane="0" entrytime="00:00:35.10" />
                <RESULT eventid="1113" points="319" reactiontime="+94" swimtime="00:02:46.83" resultid="11857" heatid="13929" lane="1" entrytime="00:02:40.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:02:06.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="244" reactiontime="+72" swimtime="00:00:38.46" resultid="11858" heatid="13953" lane="5" entrytime="00:00:38.10" />
                <RESULT eventid="1239" points="357" reactiontime="+76" swimtime="00:02:58.91" resultid="11859" heatid="13968" lane="5" entrytime="00:02:58.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="400" reactiontime="+75" swimtime="00:01:18.59" resultid="11860" heatid="14011" lane="7" entrytime="00:01:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="11861" heatid="14023" lane="3" entrytime="00:00:32.10" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="11862" heatid="14069" lane="0" entrytime="00:01:20.10" />
                <RESULT eventid="1681" points="402" swimtime="00:00:35.77" resultid="11863" heatid="14094" lane="9" entrytime="00:00:38.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="11885">
              <RESULTS>
                <RESULT eventid="1096" points="329" reactiontime="+75" swimtime="00:03:02.65" resultid="11886" heatid="13920" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:02:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="11887" heatid="13946" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1222" points="326" reactiontime="+83" swimtime="00:03:22.12" resultid="11888" heatid="13961" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                    <SPLIT distance="100" swimtime="00:01:39.34" />
                    <SPLIT distance="150" swimtime="00:02:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="340" reactiontime="+79" swimtime="00:01:32.19" resultid="11889" heatid="14003" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="254" reactiontime="+85" swimtime="00:00:38.57" resultid="11890" heatid="14016" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="11891" heatid="14064" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1664" points="325" reactiontime="+80" swimtime="00:00:42.84" resultid="11892" heatid="14085" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="11893">
              <RESULTS>
                <RESULT eventid="1113" points="366" reactiontime="+91" swimtime="00:02:39.27" resultid="11894" heatid="13927" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="400" reactiontime="+86" swimtime="00:02:52.24" resultid="11895" heatid="13969" lane="8" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="380" swimtime="00:01:19.96" resultid="11896" heatid="14011" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="320" reactiontime="+88" swimtime="00:05:56.39" resultid="11897" heatid="14061" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="150" swimtime="00:02:06.75" />
                    <SPLIT distance="200" swimtime="00:02:56.62" />
                    <SPLIT distance="250" swimtime="00:03:43.57" />
                    <SPLIT distance="300" swimtime="00:04:32.31" />
                    <SPLIT distance="350" swimtime="00:05:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="378" reactiontime="+82" swimtime="00:00:36.52" resultid="11898" heatid="14096" lane="0" entrytime="00:00:35.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="373" reactiontime="+65" swimtime="00:02:09.74" resultid="11910" heatid="13999" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:43.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11864" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="11893" number="2" />
                    <RELAYPOSITION athleteid="11855" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="11846" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="11911" heatid="13998" lane="2" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11882" number="1" />
                    <RELAYPOSITION athleteid="11871" number="2" />
                    <RELAYPOSITION athleteid="11899" number="3" />
                    <RELAYPOSITION athleteid="11874" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="416" reactiontime="+75" swimtime="00:01:53.65" resultid="11912" heatid="14056" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                    <SPLIT distance="150" swimtime="00:01:26.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11855" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="11899" number="2" />
                    <RELAYPOSITION athleteid="11864" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="11846" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="354" reactiontime="+81" swimtime="00:02:30.06" resultid="11908" heatid="13996" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:01:57.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11827" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="11885" number="2" />
                    <RELAYPOSITION athleteid="11842" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="11835" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="396" reactiontime="+83" swimtime="00:02:11.52" resultid="11909" heatid="14054" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                    <SPLIT distance="150" swimtime="00:01:38.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11842" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="11827" number="2" />
                    <RELAYPOSITION athleteid="11885" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="11835" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="341" swimtime="00:02:01.35" resultid="11904" heatid="13934" lane="6" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                    <SPLIT distance="150" swimtime="00:01:34.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11855" number="1" />
                    <RELAYPOSITION athleteid="11835" number="2" />
                    <RELAYPOSITION athleteid="11885" number="3" />
                    <RELAYPOSITION athleteid="11846" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="285" reactiontime="+70" swimtime="00:02:21.88" resultid="11906" heatid="14100" lane="2" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="150" swimtime="00:01:49.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11864" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="11893" number="2" />
                    <RELAYPOSITION athleteid="11835" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="11885" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="335" reactiontime="+89" swimtime="00:02:02.14" resultid="11905" heatid="13934" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:33.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11842" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="11864" number="2" />
                    <RELAYPOSITION athleteid="11827" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="11899" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="313" swimtime="00:02:17.51" resultid="11907" heatid="14100" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:01:50.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11827" number="1" />
                    <RELAYPOSITION athleteid="11855" number="2" />
                    <RELAYPOSITION athleteid="11842" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="11846" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="12062" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="12063">
              <RESULTS>
                <RESULT eventid="1239" points="69" reactiontime="+94" swimtime="00:05:08.51" resultid="12064" heatid="13964" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.79" />
                    <SPLIT distance="100" swimtime="00:02:29.43" />
                    <SPLIT distance="150" swimtime="00:03:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="79" reactiontime="+95" swimtime="00:01:49.29" resultid="12065" heatid="13978" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="61" swimtime="00:02:26.63" resultid="12066" heatid="14006" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="88" reactiontime="+85" swimtime="00:01:56.63" resultid="12067" heatid="14033" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="84" reactiontime="+51" swimtime="00:04:15.03" resultid="12068" heatid="14078" lane="8" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.68" />
                    <SPLIT distance="100" swimtime="00:02:08.12" />
                    <SPLIT distance="150" swimtime="00:03:14.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="12069" heatid="14107" lane="1" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="9406" name="Uks Sp 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański" phone="692076808" state="MAŁ" street="Niepodległości 7 / 46" zip="32500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="9407">
              <RESULTS>
                <RESULT eventid="1079" points="277" reactiontime="+88" swimtime="00:00:32.07" resultid="9408" heatid="13909" lane="2" entrytime="00:00:31.30" />
                <RESULT eventid="1205" points="188" reactiontime="+65" swimtime="00:00:41.92" resultid="9409" heatid="13952" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1273" points="260" reactiontime="+93" swimtime="00:01:13.43" resultid="9410" heatid="13981" lane="4" entrytime="00:01:11.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="172" reactiontime="+95" swimtime="00:01:44.14" resultid="9411" heatid="14007" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="204" reactiontime="+103" swimtime="00:02:53.04" resultid="9412" heatid="14048" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="150" swimtime="00:02:06.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="9413" heatid="14091" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="9414" heatid="14109" lane="1" entrytime="00:06:12.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="SLA" clubid="11952" name="UKS Wodnik 29 Katowice">
          <CONTACT name="Skoczylas Tomasz" />
          <ATHLETES>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="11983">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1096" points="84" reactiontime="+113" swimtime="00:04:47.48" resultid="11984" heatid="13918" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.91" />
                    <SPLIT distance="100" swimtime="00:02:22.91" />
                    <SPLIT distance="150" swimtime="00:03:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="114" reactiontime="+82" swimtime="00:00:55.67" resultid="11985" heatid="13944" lane="7" entrytime="00:01:03.00" />
                <RESULT comment="Rekord Polski" eventid="1324" points="33" reactiontime="+119" swimtime="00:06:17.77" resultid="11986" heatid="13990" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.96" />
                    <SPLIT distance="100" swimtime="00:02:56.13" />
                    <SPLIT distance="150" swimtime="00:04:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1457" points="113" reactiontime="+79" swimtime="00:02:00.14" resultid="11987" heatid="14029" lane="8" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="34" reactiontime="+110" swimtime="00:02:50.70" resultid="11988" heatid="14063" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="111" reactiontime="+92" swimtime="00:04:17.96" resultid="11989" heatid="14073" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                    <SPLIT distance="100" swimtime="00:02:04.66" />
                    <SPLIT distance="150" swimtime="00:03:12.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="11978">
              <RESULTS>
                <RESULT eventid="1079" points="304" reactiontime="+81" swimtime="00:00:31.07" resultid="11979" heatid="13908" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1239" points="321" reactiontime="+87" swimtime="00:03:05.37" resultid="11980" heatid="13967" lane="3" entrytime="00:03:06.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:01:27.53" />
                    <SPLIT distance="150" swimtime="00:02:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="330" reactiontime="+89" swimtime="00:01:23.79" resultid="11981" heatid="14010" lane="1" entrytime="00:01:21.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="405" reactiontime="+84" swimtime="00:00:35.68" resultid="11982" heatid="14096" lane="2" entrytime="00:00:35.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-05" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="11996">
              <RESULTS>
                <RESULT eventid="1079" points="476" reactiontime="+77" swimtime="00:00:26.77" resultid="11997" heatid="13915" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="527" reactiontime="+76" swimtime="00:00:58.05" resultid="11998" heatid="13988" lane="5" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="11999" heatid="14026" lane="1" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="Spławiński" nation="POL" athleteid="11993">
              <RESULTS>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="11994" heatid="14012" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1681" points="543" reactiontime="+86" swimtime="00:00:32.37" resultid="11995" heatid="14098" lane="1" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="11961">
              <RESULTS>
                <RESULT eventid="1079" points="347" reactiontime="+104" swimtime="00:00:29.75" resultid="11962" heatid="13911" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1165" points="300" reactiontime="+103" swimtime="00:21:41.06" resultid="11963" heatid="13941" lane="5" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="150" swimtime="00:02:02.13" />
                    <SPLIT distance="200" swimtime="00:02:45.72" />
                    <SPLIT distance="250" swimtime="00:03:28.82" />
                    <SPLIT distance="300" swimtime="00:04:12.57" />
                    <SPLIT distance="350" swimtime="00:04:56.00" />
                    <SPLIT distance="400" swimtime="00:05:40.24" />
                    <SPLIT distance="450" swimtime="00:06:23.62" />
                    <SPLIT distance="500" swimtime="00:07:07.92" />
                    <SPLIT distance="550" swimtime="00:07:51.19" />
                    <SPLIT distance="600" swimtime="00:08:35.03" />
                    <SPLIT distance="650" swimtime="00:09:18.48" />
                    <SPLIT distance="700" swimtime="00:10:02.37" />
                    <SPLIT distance="750" swimtime="00:10:45.48" />
                    <SPLIT distance="800" swimtime="00:11:29.48" />
                    <SPLIT distance="850" swimtime="00:12:12.83" />
                    <SPLIT distance="900" swimtime="00:12:57.22" />
                    <SPLIT distance="950" swimtime="00:13:41.29" />
                    <SPLIT distance="1000" swimtime="00:14:26.34" />
                    <SPLIT distance="1050" swimtime="00:15:10.34" />
                    <SPLIT distance="1100" swimtime="00:15:55.03" />
                    <SPLIT distance="1150" swimtime="00:16:38.86" />
                    <SPLIT distance="1200" swimtime="00:17:22.61" />
                    <SPLIT distance="1250" swimtime="00:18:05.41" />
                    <SPLIT distance="1300" swimtime="00:18:49.20" />
                    <SPLIT distance="1350" swimtime="00:19:32.79" />
                    <SPLIT distance="1400" swimtime="00:20:17.28" />
                    <SPLIT distance="1450" swimtime="00:20:58.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="357" reactiontime="+100" swimtime="00:01:06.12" resultid="11964" heatid="13983" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="196" reactiontime="+101" swimtime="00:03:11.85" resultid="11965" heatid="13994" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:19.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="264" reactiontime="+97" swimtime="00:01:20.91" resultid="11966" heatid="14036" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="261" reactiontime="+94" swimtime="00:02:39.46" resultid="11967" heatid="14049" lane="2" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                    <SPLIT distance="150" swimtime="00:01:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="222" reactiontime="+87" swimtime="00:01:22.27" resultid="11968" heatid="14069" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="299" reactiontime="+99" swimtime="00:05:29.01" resultid="11969" heatid="14110" lane="4" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="200" swimtime="00:02:39.34" />
                    <SPLIT distance="300" swimtime="00:04:05.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="11970">
              <RESULTS>
                <RESULT eventid="1079" points="100" reactiontime="+101" swimtime="00:00:45.00" resultid="11971" heatid="13904" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1205" points="75" reactiontime="+78" swimtime="00:00:56.99" resultid="11972" heatid="13950" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1239" points="55" reactiontime="+116" swimtime="00:05:32.73" resultid="11973" heatid="13964" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.08" />
                    <SPLIT distance="100" swimtime="00:02:41.59" />
                    <SPLIT distance="150" swimtime="00:04:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="51" reactiontime="+113" swimtime="00:02:36.17" resultid="11974" heatid="14005" lane="5" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="66" reactiontime="+81" swimtime="00:02:08.14" resultid="11975" heatid="14033" lane="9" entrytime="00:02:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="68" swimtime="00:04:33.15" resultid="11976" heatid="14077" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.59" />
                    <SPLIT distance="100" swimtime="00:02:15.16" />
                    <SPLIT distance="150" swimtime="00:03:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="53" reactiontime="+115" swimtime="00:01:10.08" resultid="11977" heatid="14089" lane="5" entrytime="00:01:01.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-10-10" firstname="Katarzyna" gender="F" lastname="Szczepańska" nation="POL" athleteid="11990">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="11991" heatid="13897" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="11992" heatid="14084" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="11953">
              <RESULTS>
                <RESULT eventid="1079" points="246" reactiontime="+95" swimtime="00:00:33.35" resultid="11954" heatid="13907" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1205" points="186" reactiontime="+81" swimtime="00:00:42.09" resultid="11955" heatid="13952" lane="1" entrytime="00:00:42.50" />
                <RESULT eventid="1341" points="110" reactiontime="+104" swimtime="00:03:52.52" resultid="11956" heatid="13993" lane="2" entrytime="00:03:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                    <SPLIT distance="100" swimtime="00:01:49.53" />
                    <SPLIT distance="150" swimtime="00:02:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="283" reactiontime="+93" swimtime="00:00:34.14" resultid="11957" heatid="14021" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="162" swimtime="00:03:06.93" resultid="11958" heatid="14047" lane="9" entrytime="00:03:00.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:01:31.55" />
                    <SPLIT distance="150" swimtime="00:02:21.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="154" reactiontime="+105" swimtime="00:01:32.91" resultid="11959" heatid="14067" lane="4" entrytime="00:01:31.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="150" reactiontime="+108" swimtime="00:06:53.52" resultid="11960" heatid="14108" lane="2" entrytime="00:06:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:38.79" />
                    <SPLIT distance="150" swimtime="00:02:34.31" />
                    <SPLIT distance="200" swimtime="00:03:29.38" />
                    <SPLIT distance="250" swimtime="00:04:24.38" />
                    <SPLIT distance="300" swimtime="00:05:19.00" />
                    <SPLIT distance="350" swimtime="00:06:08.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9636" name="UKS Wodnik Siemianowice Śląskie" shortname="UKS Wodnik Siemianowice Śląski">
          <CONTACT email="bartolomeo863@wp.pl" name="Szymik" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="9637">
              <RESULTS>
                <RESULT eventid="1113" points="233" reactiontime="+95" swimtime="00:03:05.01" resultid="9638" heatid="13925" lane="0" entrytime="00:03:12.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:21.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="252" swimtime="00:22:57.83" resultid="9639" heatid="13941" lane="6" entrytime="00:22:31.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                    <SPLIT distance="150" swimtime="00:02:11.33" />
                    <SPLIT distance="200" swimtime="00:02:56.89" />
                    <SPLIT distance="250" swimtime="00:03:43.06" />
                    <SPLIT distance="300" swimtime="00:04:29.38" />
                    <SPLIT distance="350" swimtime="00:05:15.95" />
                    <SPLIT distance="400" swimtime="00:06:01.44" />
                    <SPLIT distance="450" swimtime="00:06:48.71" />
                    <SPLIT distance="500" swimtime="00:07:34.67" />
                    <SPLIT distance="550" swimtime="00:08:21.56" />
                    <SPLIT distance="600" swimtime="00:09:07.10" />
                    <SPLIT distance="650" swimtime="00:09:54.50" />
                    <SPLIT distance="700" swimtime="00:10:40.94" />
                    <SPLIT distance="750" swimtime="00:11:27.20" />
                    <SPLIT distance="800" swimtime="00:12:13.35" />
                    <SPLIT distance="850" swimtime="00:12:59.37" />
                    <SPLIT distance="900" swimtime="00:13:45.69" />
                    <SPLIT distance="950" swimtime="00:14:32.85" />
                    <SPLIT distance="1000" swimtime="00:15:19.21" />
                    <SPLIT distance="1050" swimtime="00:16:06.29" />
                    <SPLIT distance="1100" swimtime="00:16:52.49" />
                    <SPLIT distance="1150" swimtime="00:17:40.03" />
                    <SPLIT distance="1200" swimtime="00:18:27.43" />
                    <SPLIT distance="1250" swimtime="00:19:14.43" />
                    <SPLIT distance="1300" swimtime="00:19:59.74" />
                    <SPLIT distance="1350" swimtime="00:20:46.55" />
                    <SPLIT distance="1400" swimtime="00:21:32.80" />
                    <SPLIT distance="1450" swimtime="00:22:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="159" swimtime="00:03:25.52" resultid="9640" heatid="13994" lane="9" entrytime="00:03:19.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:37.88" />
                    <SPLIT distance="150" swimtime="00:02:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="218" reactiontime="+86" swimtime="00:00:37.26" resultid="9641" heatid="14021" lane="0" entrytime="00:00:35.24" />
                <RESULT eventid="1578" points="197" reactiontime="+97" swimtime="00:06:58.48" resultid="9642" heatid="14061" lane="0" entrytime="00:06:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:43.67" />
                    <SPLIT distance="150" swimtime="00:02:36.37" />
                    <SPLIT distance="200" swimtime="00:03:28.84" />
                    <SPLIT distance="250" swimtime="00:04:28.93" />
                    <SPLIT distance="300" swimtime="00:05:27.37" />
                    <SPLIT distance="350" swimtime="00:06:13.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="172" reactiontime="+100" swimtime="00:01:29.52" resultid="9643" heatid="14068" lane="1" entrytime="00:01:28.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="234" reactiontime="+98" swimtime="00:05:57.01" resultid="9644" heatid="14110" lane="2" entrytime="00:05:45.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:08.83" />
                    <SPLIT distance="200" swimtime="00:02:55.12" />
                    <SPLIT distance="250" swimtime="00:03:42.45" />
                    <SPLIT distance="300" swimtime="00:04:29.00" />
                    <SPLIT distance="350" swimtime="00:05:14.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="12414" name="Uniwersytet Śląski Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1950-09-19" firstname="Wiesław" gender="M" lastname="Majcher" nation="POL" athleteid="12415">
              <RESULTS>
                <RESULT eventid="1113" points="62" reactiontime="+108" swimtime="00:04:47.14" resultid="12416" heatid="13922" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:02:31.60" />
                    <SPLIT distance="150" swimtime="00:03:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="(Time: 20:11), Przekroczony regulaminowy limit czasu." eventid="1165" status="OTL" swimtime="00:00:00.00" resultid="12417" heatid="13940" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                    <SPLIT distance="100" swimtime="00:01:54.82" />
                    <SPLIT distance="150" swimtime="00:03:05.88" />
                    <SPLIT distance="200" swimtime="00:04:26.92" />
                    <SPLIT distance="250" swimtime="00:05:53.07" />
                    <SPLIT distance="300" swimtime="00:06:55.50" />
                    <SPLIT distance="350" swimtime="00:08:04.50" />
                    <SPLIT distance="400" swimtime="00:09:11.70" />
                    <SPLIT distance="450" swimtime="00:10:38.39" />
                    <SPLIT distance="500" swimtime="00:11:40.66" />
                    <SPLIT distance="550" swimtime="00:12:48.50" />
                    <SPLIT distance="600" swimtime="00:14:08.80" />
                    <SPLIT distance="650" swimtime="00:15:16.79" />
                    <SPLIT distance="700" swimtime="00:16:23.00" />
                    <SPLIT distance="750" swimtime="00:17:29.18" />
                    <SPLIT distance="800" swimtime="00:18:52.41" />
                    <SPLIT distance="850" swimtime="00:19:59.10" />
                    <SPLIT distance="900" swimtime="00:21:07.59" />
                    <SPLIT distance="950" swimtime="00:22:28.51" />
                    <SPLIT distance="1000" swimtime="00:23:40.32" />
                    <SPLIT distance="1050" swimtime="00:24:50.23" />
                    <SPLIT distance="1100" swimtime="00:26:18.42" />
                    <SPLIT distance="1150" swimtime="00:27:29.28" />
                    <SPLIT distance="1200" swimtime="00:28:49.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="61" reactiontime="+100" swimtime="00:01:00.94" resultid="12418" heatid="13950" lane="0" entrytime="00:01:00.16" />
                <RESULT eventid="1239" points="79" reactiontime="+116" swimtime="00:04:55.31" resultid="12419" heatid="13963" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.15" />
                    <SPLIT distance="100" swimtime="00:02:19.38" />
                    <SPLIT distance="150" swimtime="00:03:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="81" reactiontime="+126" swimtime="00:02:13.84" resultid="12420" heatid="14006" lane="0" entrytime="00:02:14.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="47" reactiontime="+109" swimtime="00:01:02.08" resultid="12421" heatid="14019" lane="8" entrytime="00:00:56.89" />
                <RESULT eventid="1681" points="109" reactiontime="+107" swimtime="00:00:55.24" resultid="12422" heatid="14090" lane="0" entrytime="00:00:56.19" />
                <RESULT eventid="1744" reactiontime="+122" status="DNF" swimtime="00:00:00.00" resultid="12423" heatid="14106" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.26" />
                    <SPLIT distance="150" swimtime="00:03:02.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="12191" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1968-06-01" firstname="Robert" gender="M" lastname="Zieliński" nation="POL" athleteid="12211">
              <RESULTS>
                <RESULT eventid="1079" points="254" reactiontime="+85" swimtime="00:00:33.00" resultid="12212" heatid="13908" lane="2" entrytime="00:00:32.89" />
                <RESULT eventid="1113" points="154" reactiontime="+84" swimtime="00:03:32.53" resultid="12213" heatid="13925" lane="5" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="188" reactiontime="+76" swimtime="00:00:41.94" resultid="12214" heatid="13952" lane="3" entrytime="00:00:41.34" />
                <RESULT eventid="1273" points="232" reactiontime="+89" swimtime="00:01:16.29" resultid="12215" heatid="13980" lane="7" entrytime="00:01:17.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="185" reactiontime="+93" swimtime="00:00:39.34" resultid="12216" heatid="14020" lane="0" entrytime="00:00:38.57" />
                <RESULT eventid="1474" points="121" reactiontime="+70" swimtime="00:01:44.92" resultid="12217" heatid="14034" lane="9" entrytime="00:01:39.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="12218" heatid="14078" lane="2" entrytime="00:03:42.27" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="12219" heatid="14091" lane="9" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="12192">
              <RESULTS>
                <RESULT eventid="1113" points="211" reactiontime="+88" swimtime="00:03:11.29" resultid="12193" heatid="13925" lane="3" entrytime="00:03:09.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:35.11" />
                    <SPLIT distance="150" swimtime="00:02:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="259" reactiontime="+95" swimtime="00:03:19.25" resultid="12194" heatid="13967" lane="8" entrytime="00:03:17.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="100" swimtime="00:01:35.33" />
                    <SPLIT distance="150" swimtime="00:02:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="291" reactiontime="+96" swimtime="00:01:27.39" resultid="12195" heatid="14008" lane="4" entrytime="00:01:26.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="335" reactiontime="+94" swimtime="00:00:38.03" resultid="12196" heatid="14094" lane="7" entrytime="00:00:37.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="12197">
              <RESULTS>
                <RESULT eventid="1079" points="314" reactiontime="+91" swimtime="00:00:30.74" resultid="12198" heatid="13911" lane="3" entrytime="00:00:29.30" />
                <RESULT eventid="1205" points="116" reactiontime="+83" swimtime="00:00:49.22" resultid="12199" heatid="13952" lane="2" entrytime="00:00:41.98" />
                <RESULT eventid="1273" points="302" reactiontime="+95" swimtime="00:01:09.87" resultid="12200" heatid="13984" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="240" reactiontime="+91" swimtime="00:00:36.09" resultid="12201" heatid="14022" lane="0" entrytime="00:00:33.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="12202" heatid="14049" lane="6" entrytime="00:02:32.48" />
                <RESULT eventid="1613" points="195" reactiontime="+86" swimtime="00:01:25.88" resultid="12203" heatid="14068" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="228" reactiontime="+102" swimtime="00:06:00.05" resultid="12204" heatid="14107" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:06.92" />
                    <SPLIT distance="200" swimtime="00:02:54.07" />
                    <SPLIT distance="250" swimtime="00:03:41.94" />
                    <SPLIT distance="300" swimtime="00:04:31.08" />
                    <SPLIT distance="350" swimtime="00:05:18.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="Rybarczyk" nation="POL" athleteid="12205">
              <RESULTS>
                <RESULT eventid="1079" points="99" reactiontime="+101" swimtime="00:00:45.15" resultid="12206" heatid="13905" lane="6" entrytime="00:00:41.27" />
                <RESULT eventid="1205" points="78" reactiontime="+102" swimtime="00:00:56.10" resultid="12207" heatid="13951" lane="9" entrytime="00:00:53.84" />
                <RESULT eventid="1406" points="131" reactiontime="+105" swimtime="00:01:53.98" resultid="12208" heatid="14006" lane="6" entrytime="00:01:50.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="60" reactiontime="+94" swimtime="00:02:12.43" resultid="12209" heatid="14033" lane="3" entrytime="00:01:57.99" />
                <RESULT eventid="1681" points="159" reactiontime="+109" swimtime="00:00:48.74" resultid="12210" heatid="14090" lane="2" entrytime="00:00:49.84" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="189" reactiontime="+60" swimtime="00:02:42.56" resultid="12220" heatid="13998" lane="9" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="150" swimtime="00:01:58.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12211" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="12192" number="2" />
                    <RELAYPOSITION athleteid="12197" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="12205" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="232" reactiontime="+81" swimtime="00:02:17.91" resultid="12221" heatid="14055" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:01:47.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12192" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="12205" number="2" />
                    <RELAYPOSITION athleteid="12211" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="12197" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="031" nation="POL" region="LOD" clubid="9472" name="UTW &quot;Masters&quot;Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmai.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="9484">
              <RESULTS>
                <RESULT eventid="1239" points="149" reactiontime="+110" swimtime="00:03:59.46" resultid="9485" heatid="13965" lane="5" entrytime="00:03:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                    <SPLIT distance="100" swimtime="00:01:51.51" />
                    <SPLIT distance="150" swimtime="00:02:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="186" reactiontime="+105" swimtime="00:01:41.31" resultid="9486" heatid="14007" lane="5" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="260" reactiontime="+107" swimtime="00:00:41.35" resultid="9487" heatid="14092" lane="8" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="9533">
              <RESULTS>
                <RESULT eventid="1079" points="550" reactiontime="+71" swimtime="00:00:25.51" resultid="9534" heatid="13917" lane="5" entrytime="00:00:24.70" entrycourse="LCM" />
                <RESULT eventid="1113" points="501" reactiontime="+76" swimtime="00:02:23.47" resultid="9535" heatid="13931" lane="4" entrytime="00:02:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:45.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="559" reactiontime="+73" swimtime="00:00:56.93" resultid="9536" heatid="13989" lane="4" entrytime="00:00:53.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="575" reactiontime="+76" swimtime="00:00:26.97" resultid="9537" heatid="14027" lane="4" entrytime="00:00:25.80" entrycourse="LCM" />
                <RESULT eventid="1508" points="529" reactiontime="+75" swimtime="00:02:06.05" resultid="9538" heatid="14053" lane="4" entrytime="00:01:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="550" reactiontime="+78" swimtime="00:01:00.77" resultid="9539" heatid="14071" lane="4" entrytime="00:00:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="521" reactiontime="+74" swimtime="00:00:32.83" resultid="9540" heatid="14098" lane="4" entrytime="00:00:29.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="9552">
              <RESULTS>
                <RESULT eventid="1062" points="521" reactiontime="+90" swimtime="00:00:29.49" resultid="9553" heatid="13900" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski" eventid="1096" points="511" reactiontime="+68" swimtime="00:02:37.72" resultid="9554" heatid="13920" lane="3" entrytime="00:03:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1187" points="564" reactiontime="+72" swimtime="00:00:32.74" resultid="9555" heatid="13948" lane="6" entrytime="00:00:33.60" entrycourse="LCM" />
                <RESULT eventid="1256" points="478" reactiontime="+91" swimtime="00:01:06.56" resultid="9556" heatid="13976" lane="3" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="457" reactiontime="+83" swimtime="00:00:31.70" resultid="9557" heatid="14017" lane="3" entrytime="00:00:31.70" entrycourse="LCM" />
                <RESULT eventid="1457" points="528" swimtime="00:01:11.87" resultid="9558" heatid="14031" lane="4" entrytime="00:01:09.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="436" reactiontime="+86" swimtime="00:01:13.33" resultid="9559" heatid="14065" lane="4" entrytime="00:01:10.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="428" reactiontime="+88" swimtime="00:02:44.54" resultid="9560" heatid="14075" lane="5" entrytime="00:02:39.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                    <SPLIT distance="150" swimtime="00:02:01.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="9541">
              <RESULTS>
                <RESULT eventid="1096" points="423" reactiontime="+83" swimtime="00:02:47.97" resultid="9542" heatid="13921" lane="5" entrytime="00:02:43.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:07.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="321" reactiontime="+93" swimtime="00:02:57.81" resultid="9543" heatid="13991" lane="4" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="150" swimtime="00:02:05.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="374" reactiontime="+85" swimtime="00:01:29.24" resultid="9544" heatid="14004" lane="8" entrytime="00:01:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="386" reactiontime="+90" swimtime="00:00:33.54" resultid="9545" heatid="14017" lane="1" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1595" points="408" reactiontime="+89" swimtime="00:01:14.97" resultid="9546" heatid="14065" lane="3" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="9504">
              <RESULTS>
                <RESULT eventid="1062" points="368" reactiontime="+93" swimtime="00:00:33.10" resultid="9505" heatid="13900" lane="1" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="338" reactiontime="+78" swimtime="00:00:38.84" resultid="9506" heatid="13947" lane="0" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1324" points="202" reactiontime="+101" swimtime="00:03:27.34" resultid="9507" heatid="13991" lane="0" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:40.02" />
                    <SPLIT distance="150" swimtime="00:02:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="319" reactiontime="+92" swimtime="00:00:35.75" resultid="9508" heatid="14016" lane="4" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1457" points="225" reactiontime="+77" swimtime="00:01:35.49" resultid="9509" heatid="14030" lane="2" entrytime="00:01:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="191" swimtime="00:01:36.53" resultid="9510" heatid="14065" lane="9" entrytime="00:01:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="207" reactiontime="+75" swimtime="00:03:29.40" resultid="9511" heatid="14074" lane="7" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.29" />
                    <SPLIT distance="100" swimtime="00:01:44.22" />
                    <SPLIT distance="150" swimtime="00:02:38.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="9526">
              <RESULTS>
                <RESULT eventid="1079" points="254" reactiontime="+93" swimtime="00:00:32.98" resultid="9527" heatid="13908" lane="7" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="134" reactiontime="+103" swimtime="00:03:42.37" resultid="9528" heatid="13923" lane="6" entrytime="00:03:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:52.52" />
                    <SPLIT distance="150" swimtime="00:02:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="9529" heatid="13980" lane="2" entrytime="00:01:16.00" entrycourse="LCM" />
                <RESULT eventid="1341" points="67" reactiontime="+99" swimtime="00:04:34.46" resultid="9530" heatid="13992" lane="3" entrytime="00:04:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.12" />
                    <SPLIT distance="100" swimtime="00:02:15.48" />
                    <SPLIT distance="150" swimtime="00:03:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="223" reactiontime="+86" swimtime="00:00:36.98" resultid="9531" heatid="14020" lane="7" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1613" points="102" reactiontime="+95" swimtime="00:01:46.53" resultid="9532" heatid="14067" lane="1" entrytime="00:01:44.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-08" firstname="Piotr" gender="M" lastname="Kapczyński" nation="POL" license="503105700043" athleteid="9547">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="9548" heatid="13968" lane="2" entrytime="00:03:00.00" entrycourse="LCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="9549" heatid="14010" lane="9" entrytime="00:01:23.90" entrycourse="LCM" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="9550" heatid="14022" lane="8" entrytime="00:00:33.14" entrycourse="LCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="9551" heatid="14094" lane="5" entrytime="00:00:37.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-11" firstname="Jakub" gender="M" lastname="Jurek" nation="POL" license="503105700048" athleteid="9518">
              <RESULTS>
                <RESULT eventid="1205" points="323" reactiontime="+63" swimtime="00:00:35.01" resultid="9519" heatid="13956" lane="9" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="9520" heatid="14037" lane="0" entrytime="00:01:13.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="9473">
              <RESULTS>
                <RESULT eventid="1205" points="71" reactiontime="+88" swimtime="00:00:58.05" resultid="9474" heatid="13950" lane="5" entrytime="00:00:55.68" entrycourse="LCM" />
                <RESULT eventid="1273" points="140" reactiontime="+90" swimtime="00:01:30.27" resultid="9475" heatid="13979" lane="0" entrytime="00:01:32.05" entrycourse="LCM" />
                <RESULT eventid="1474" points="60" reactiontime="+101" swimtime="00:02:12.27" resultid="9476" heatid="14033" lane="2" entrytime="00:02:03.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="100" reactiontime="+108" swimtime="00:03:39.35" resultid="9477" heatid="14046" lane="0" entrytime="00:03:34.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="59" swimtime="00:04:47.33" resultid="9478" heatid="14077" lane="7" entrytime="00:04:35.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.29" />
                    <SPLIT distance="100" swimtime="00:02:22.75" />
                    <SPLIT distance="150" swimtime="00:03:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="102" reactiontime="+113" swimtime="00:07:50.59" resultid="9479" heatid="14107" lane="7" entrytime="00:07:54.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.56" />
                    <SPLIT distance="200" swimtime="00:03:53.53" />
                    <SPLIT distance="300" swimtime="00:05:56.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Wożniak" nation="POL" license="503105700039" athleteid="9521">
              <RESULTS>
                <RESULT eventid="1113" points="309" swimtime="00:02:48.60" resultid="9522" heatid="13929" lane="9" entrytime="00:02:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                    <SPLIT distance="150" swimtime="00:02:05.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="395" reactiontime="+66" swimtime="00:00:32.75" resultid="9523" heatid="13957" lane="7" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="392" reactiontime="+70" swimtime="00:01:10.96" resultid="9524" heatid="14037" lane="3" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="341" reactiontime="+76" swimtime="00:02:40.15" resultid="9525" heatid="14081" lane="1" entrytime="00:02:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:15.81" />
                    <SPLIT distance="150" swimtime="00:01:58.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="9480">
              <RESULTS>
                <RESULT eventid="1239" points="199" reactiontime="+102" swimtime="00:03:37.40" resultid="9481" heatid="13966" lane="8" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:45.58" />
                    <SPLIT distance="150" swimtime="00:02:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="219" reactiontime="+101" swimtime="00:01:36.07" resultid="9482" heatid="14008" lane="2" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="253" swimtime="00:00:41.72" resultid="9483" heatid="14093" lane="9" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-13" firstname="Mirosława" gender="F" lastname="Rajtar" nation="POL" license="503105600020" athleteid="9497">
              <RESULTS>
                <RESULT eventid="1062" points="234" reactiontime="+99" swimtime="00:00:38.48" resultid="9498" heatid="13898" lane="6" entrytime="00:00:39.20" entrycourse="LCM" />
                <RESULT eventid="1187" points="192" swimtime="00:00:46.84" resultid="9499" heatid="13945" lane="6" entrytime="00:00:48.60" entrycourse="LCM" />
                <RESULT eventid="1256" points="209" reactiontime="+100" swimtime="00:01:27.61" resultid="9500" heatid="13972" lane="6" entrytime="00:01:30.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="163" reactiontime="+93" swimtime="00:00:44.64" resultid="9501" heatid="14015" lane="7" entrytime="00:00:45.80" entrycourse="LCM" />
                <RESULT eventid="1491" points="179" reactiontime="+101" swimtime="00:03:20.10" resultid="9502" heatid="14040" lane="2" entrytime="00:03:20.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="166" reactiontime="+102" swimtime="00:00:53.60" resultid="9503" heatid="14083" lane="5" entrytime="00:00:54.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" license="503105700049" athleteid="10889">
              <RESULTS>
                <RESULT eventid="1079" points="549" reactiontime="+74" swimtime="00:00:25.53" resultid="10890" heatid="13917" lane="4" entrytime="00:00:24.50" entrycourse="LCM" />
                <RESULT eventid="1440" points="554" reactiontime="+70" swimtime="00:00:27.30" resultid="10891" heatid="14027" lane="5" entrytime="00:00:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="9512">
              <RESULTS>
                <RESULT eventid="1062" points="387" reactiontime="+80" swimtime="00:00:32.56" resultid="9513" heatid="13900" lane="0" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="330" reactiontime="+78" swimtime="00:01:15.34" resultid="9514" heatid="13974" lane="8" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="357" reactiontime="+85" swimtime="00:01:30.68" resultid="9515" heatid="14003" lane="7" entrytime="00:01:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="9516" heatid="14040" lane="5" entrytime="00:03:02.00" entrycourse="LCM" />
                <RESULT eventid="1664" points="388" swimtime="00:00:40.41" resultid="9517" heatid="14086" lane="9" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700026" athleteid="9488">
              <RESULTS>
                <RESULT eventid="1079" points="306" reactiontime="+86" swimtime="00:00:31.02" resultid="9489" heatid="13910" lane="2" entrytime="00:00:30.50" entrycourse="LCM" />
                <RESULT eventid="1113" points="265" reactiontime="+86" swimtime="00:02:57.30" resultid="9490" heatid="13926" lane="6" entrytime="00:02:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="294" reactiontime="+75" swimtime="00:00:36.15" resultid="9491" heatid="13954" lane="2" entrytime="00:00:36.50" entrycourse="LCM" />
                <RESULT eventid="1341" points="198" reactiontime="+87" swimtime="00:03:11.07" resultid="9492" heatid="13994" lane="5" entrytime="00:03:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="150" swimtime="00:02:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="311" swimtime="00:00:33.09" resultid="9493" heatid="14022" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="9494" heatid="14049" lane="5" entrytime="00:02:32.00" entrycourse="LCM" />
                <RESULT eventid="1613" points="227" reactiontime="+86" swimtime="00:01:21.61" resultid="9495" heatid="14069" lane="7" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="9496" heatid="14110" lane="5" entrytime="00:05:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="9561" heatid="13998" lane="5" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9521" number="1" />
                    <RELAYPOSITION athleteid="9484" number="2" />
                    <RELAYPOSITION athleteid="9533" number="3" />
                    <RELAYPOSITION athleteid="9547" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="9562" heatid="14056" lane="9" entrytime="00:02:03.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9547" number="1" />
                    <RELAYPOSITION athleteid="9484" number="2" />
                    <RELAYPOSITION athleteid="9521" number="3" />
                    <RELAYPOSITION athleteid="9533" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="263" reactiontime="+63" swimtime="00:02:25.78" resultid="9563" heatid="13998" lane="6" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:16.48" />
                    <SPLIT distance="150" swimtime="00:01:51.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9518" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="9480" number="2" />
                    <RELAYPOSITION athleteid="9488" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9526" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="268" reactiontime="+75" swimtime="00:02:11.57" resultid="9564" heatid="14055" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:06.45" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9518" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9480" number="2" />
                    <RELAYPOSITION athleteid="9526" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="9488" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1358" points="419" reactiontime="+68" swimtime="00:02:21.93" resultid="9569" heatid="13996" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9552" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="9512" number="2" />
                    <RELAYPOSITION athleteid="9541" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="9504" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1525" points="449" reactiontime="+85" swimtime="00:02:06.07" resultid="9570" heatid="14054" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9541" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="9504" number="2" />
                    <RELAYPOSITION athleteid="9512" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="9552" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="374" reactiontime="+75" swimtime="00:01:57.74" resultid="9565" heatid="13934" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.34" />
                    <SPLIT distance="100" swimtime="00:00:56.65" />
                    <SPLIT distance="150" swimtime="00:01:28.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10889" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9541" number="2" />
                    <RELAYPOSITION athleteid="9488" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="9552" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1698" points="382" reactiontime="+69" swimtime="00:02:08.67" resultid="9566" heatid="14101" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9552" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="9533" number="2" />
                    <RELAYPOSITION athleteid="9541" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="9488" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="228" reactiontime="+94" swimtime="00:02:18.87" resultid="9567" heatid="13933" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:11.59" />
                    <SPLIT distance="150" swimtime="00:01:46.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9504" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="9480" number="2" />
                    <RELAYPOSITION athleteid="9526" number="3" reactiontime="+83" />
                    <RELAYPOSITION athleteid="9512" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="220" reactiontime="+73" swimtime="00:02:34.56" resultid="9568" heatid="14101" lane="8" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9504" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="9480" number="2" />
                    <RELAYPOSITION athleteid="9512" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="9526" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="9825" name="Victory Masters Elbąg">
          <CONTACT city="Elbląg" email="lateccy@o2.pl" name="Latecki" phone="606147184" state="WM" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="9833">
              <RESULTS>
                <RESULT eventid="1062" points="159" reactiontime="+104" swimtime="00:00:43.72" resultid="9834" heatid="13897" lane="6" entrytime="00:00:44.00" />
                <RESULT comment="(Time: 18:49), Przekroczony regulaminowy limit czasu." eventid="1147" reactiontime="+112" status="OTL" swimtime="00:15:16.12" resultid="9835" heatid="13936" lane="2" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                    <SPLIT distance="100" swimtime="00:01:50.17" />
                    <SPLIT distance="150" swimtime="00:02:48.02" />
                    <SPLIT distance="200" swimtime="00:03:47.33" />
                    <SPLIT distance="250" swimtime="00:04:46.36" />
                    <SPLIT distance="300" swimtime="00:05:46.38" />
                    <SPLIT distance="350" swimtime="00:06:44.46" />
                    <SPLIT distance="400" swimtime="00:07:43.74" />
                    <SPLIT distance="450" swimtime="00:08:41.61" />
                    <SPLIT distance="500" swimtime="00:09:40.05" />
                    <SPLIT distance="550" swimtime="00:10:37.02" />
                    <SPLIT distance="600" swimtime="00:11:35.13" />
                    <SPLIT distance="650" swimtime="00:12:32.29" />
                    <SPLIT distance="700" swimtime="00:13:28.73" />
                    <SPLIT distance="750" swimtime="00:14:23.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="156" swimtime="00:01:36.55" resultid="9836" heatid="13972" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="153" reactiontime="+98" swimtime="00:03:31.11" resultid="9837" heatid="14040" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                    <SPLIT distance="100" swimtime="00:01:46.10" />
                    <SPLIT distance="150" swimtime="00:02:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="151" reactiontime="+109" swimtime="00:07:27.01" resultid="9838" heatid="14103" lane="1" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.39" />
                    <SPLIT distance="100" swimtime="00:01:51.63" />
                    <SPLIT distance="150" swimtime="00:02:50.21" />
                    <SPLIT distance="200" swimtime="00:03:48.79" />
                    <SPLIT distance="250" swimtime="00:04:46.03" />
                    <SPLIT distance="300" swimtime="00:05:42.77" />
                    <SPLIT distance="350" swimtime="00:06:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="9839">
              <RESULTS>
                <RESULT eventid="1096" points="115" reactiontime="+109" swimtime="00:04:18.68" resultid="9840" heatid="13919" lane="0" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.29" />
                    <SPLIT distance="100" swimtime="00:02:10.46" />
                    <SPLIT distance="150" swimtime="00:03:24.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="162" swimtime="00:14:52.89" resultid="9841" heatid="13936" lane="9" entrytime="00:14:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.64" />
                    <SPLIT distance="100" swimtime="00:01:46.36" />
                    <SPLIT distance="150" swimtime="00:02:42.83" />
                    <SPLIT distance="200" swimtime="00:03:39.59" />
                    <SPLIT distance="250" swimtime="00:04:36.22" />
                    <SPLIT distance="300" swimtime="00:05:33.46" />
                    <SPLIT distance="350" swimtime="00:06:30.34" />
                    <SPLIT distance="400" swimtime="00:07:27.29" />
                    <SPLIT distance="450" swimtime="00:08:24.05" />
                    <SPLIT distance="500" swimtime="00:09:21.37" />
                    <SPLIT distance="550" swimtime="00:10:17.83" />
                    <SPLIT distance="600" swimtime="00:11:13.88" />
                    <SPLIT distance="650" swimtime="00:12:09.38" />
                    <SPLIT distance="700" swimtime="00:13:04.67" />
                    <SPLIT distance="750" swimtime="00:13:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="135" reactiontime="+103" swimtime="00:01:41.27" resultid="9842" heatid="13972" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="98" reactiontime="+107" swimtime="00:04:23.59" resultid="9843" heatid="13990" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.95" />
                    <SPLIT distance="100" swimtime="00:02:04.53" />
                    <SPLIT distance="150" swimtime="00:03:14.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 18:07)" eventid="1491" reactiontime="+79" status="DSQ" swimtime="00:03:33.51" resultid="9844" heatid="14040" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:44.33" />
                    <SPLIT distance="150" swimtime="00:02:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="123" reactiontime="+130" swimtime="00:08:58.39" resultid="9845" heatid="14057" lane="4" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.02" />
                    <SPLIT distance="150" swimtime="00:03:23.77" />
                    <SPLIT distance="250" swimtime="00:05:52.00" />
                    <SPLIT distance="350" swimtime="00:08:05.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="95" reactiontime="+124" swimtime="00:02:01.86" resultid="9846" heatid="14063" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="168" reactiontime="+119" swimtime="00:07:11.96" resultid="9847" heatid="14102" lane="4" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.97" />
                    <SPLIT distance="100" swimtime="00:01:44.17" />
                    <SPLIT distance="150" swimtime="00:02:39.14" />
                    <SPLIT distance="200" swimtime="00:03:34.23" />
                    <SPLIT distance="250" swimtime="00:04:29.77" />
                    <SPLIT distance="300" swimtime="00:05:24.89" />
                    <SPLIT distance="350" swimtime="00:06:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="9848">
              <RESULTS>
                <RESULT eventid="1062" points="71" reactiontime="+137" swimtime="00:00:57.05" resultid="9849" heatid="13896" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="1147" reactiontime="+113" status="DNF" swimtime="00:00:00.00" resultid="9850" heatid="13935" lane="2" entrytime="00:18:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.22" />
                    <SPLIT distance="100" swimtime="00:02:11.09" />
                    <SPLIT distance="150" swimtime="00:03:28.05" />
                    <SPLIT distance="200" swimtime="00:04:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="66" reactiontime="+75" swimtime="00:01:06.77" resultid="9851" heatid="13944" lane="8" entrytime="00:01:05.00" />
                <RESULT eventid="1222" points="71" reactiontime="+110" swimtime="00:05:35.79" resultid="9852" heatid="13959" lane="5" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.24" />
                    <SPLIT distance="100" swimtime="00:02:47.83" />
                    <SPLIT distance="150" swimtime="00:04:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="61" reactiontime="+106" swimtime="00:02:42.67" resultid="9853" heatid="14000" lane="3" entrytime="00:02:36.00" />
                <RESULT eventid="1457" points="60" reactiontime="+111" swimtime="00:02:28.20" resultid="9854" heatid="14028" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="54" reactiontime="+103" swimtime="00:05:27.58" resultid="9855" heatid="14072" lane="4" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.85" />
                    <SPLIT distance="100" swimtime="00:02:31.42" />
                    <SPLIT distance="150" swimtime="00:03:58.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" reactiontime="+112" status="DNF" swimtime="00:00:00.00" resultid="9856" heatid="14102" lane="6" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.19" />
                    <SPLIT distance="100" swimtime="00:02:18.77" />
                    <SPLIT distance="150" swimtime="00:03:37.49" />
                    <SPLIT distance="200" swimtime="00:04:57.04" />
                    <SPLIT distance="250" swimtime="00:06:16.93" />
                    <SPLIT distance="300" swimtime="00:07:37.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="9826">
              <RESULTS>
                <RESULT eventid="1079" points="423" reactiontime="+85" swimtime="00:00:27.85" resultid="9827" heatid="13911" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="390" reactiontime="+82" swimtime="00:02:35.91" resultid="9828" heatid="13928" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="390" reactiontime="+66" swimtime="00:00:32.89" resultid="9829" heatid="13955" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="9830" heatid="13984" lane="1" entrytime="00:01:04.50" />
                <RESULT eventid="1440" points="472" reactiontime="+83" swimtime="00:00:28.79" resultid="9831" heatid="14024" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1578" points="331" reactiontime="+103" swimtime="00:05:52.46" resultid="9832" heatid="14061" lane="1" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                    <SPLIT distance="200" swimtime="00:02:54.02" />
                    <SPLIT distance="250" swimtime="00:03:44.05" />
                    <SPLIT distance="300" swimtime="00:04:34.84" />
                    <SPLIT distance="350" swimtime="00:05:14.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="10164" name="Warsaw Masters team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 4444" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="10275">
              <RESULTS>
                <RESULT eventid="1062" points="384" reactiontime="+68" swimtime="00:00:32.62" resultid="10276" heatid="13900" lane="4" entrytime="00:00:32.40" />
                <RESULT eventid="1222" points="288" reactiontime="+69" swimtime="00:03:30.60" resultid="10277" heatid="13961" lane="7" entrytime="00:03:25.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                    <SPLIT distance="100" swimtime="00:01:42.53" />
                    <SPLIT distance="150" swimtime="00:02:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="325" reactiontime="+72" swimtime="00:01:33.54" resultid="10278" heatid="14003" lane="1" entrytime="00:01:32.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="373" reactiontime="+63" swimtime="00:00:40.94" resultid="10279" heatid="14086" lane="2" entrytime="00:00:40.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-31" firstname="Katharina" gender="F" lastname="Szymańska" nation="POL" athleteid="10341">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="10342" heatid="13898" lane="5" entrytime="00:00:38.50" />
                <RESULT eventid="1096" points="207" reactiontime="+87" swimtime="00:03:32.87" resultid="10343" heatid="13919" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:45.09" />
                    <SPLIT distance="150" swimtime="00:02:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="225" reactiontime="+89" swimtime="00:01:25.61" resultid="10344" heatid="13973" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="10345" heatid="14015" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="10210">
              <RESULTS>
                <RESULT eventid="1079" points="360" reactiontime="+94" swimtime="00:00:29.37" resultid="10211" heatid="13912" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="310" reactiontime="+97" swimtime="00:02:48.27" resultid="10212" heatid="13927" lane="8" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:11.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="243" reactiontime="+92" swimtime="00:00:38.50" resultid="10213" heatid="13954" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1273" points="366" swimtime="00:01:05.58" resultid="10214" heatid="13984" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="10215" heatid="14021" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1508" points="360" reactiontime="+86" swimtime="00:02:23.33" resultid="10216" heatid="14050" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10217" heatid="14092" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1744" points="344" swimtime="00:05:13.86" resultid="10218" heatid="14111" lane="6" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:52.42" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:13.81" />
                    <SPLIT distance="300" swimtime="00:03:55.40" />
                    <SPLIT distance="350" swimtime="00:04:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="10337">
              <RESULTS>
                <RESULT eventid="1079" points="452" reactiontime="+79" swimtime="00:00:27.23" resultid="10338" heatid="13915" lane="0" entrytime="00:00:26.70" />
                <RESULT eventid="1113" points="413" reactiontime="+87" swimtime="00:02:33.05" resultid="10339" heatid="13931" lane="0" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" reactiontime="+101" status="DSQ" swimtime="00:19:30.13" resultid="10340" heatid="13939" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:52.35" />
                    <SPLIT distance="200" swimtime="00:02:31.57" />
                    <SPLIT distance="250" swimtime="00:03:10.95" />
                    <SPLIT distance="300" swimtime="00:03:50.58" />
                    <SPLIT distance="350" swimtime="00:04:29.73" />
                    <SPLIT distance="400" swimtime="00:05:09.37" />
                    <SPLIT distance="450" swimtime="00:05:47.56" />
                    <SPLIT distance="500" swimtime="00:06:26.09" />
                    <SPLIT distance="550" swimtime="00:07:05.03" />
                    <SPLIT distance="600" swimtime="00:07:44.32" />
                    <SPLIT distance="650" swimtime="00:08:23.27" />
                    <SPLIT distance="700" swimtime="00:09:02.37" />
                    <SPLIT distance="750" swimtime="00:09:41.77" />
                    <SPLIT distance="800" swimtime="00:10:21.32" />
                    <SPLIT distance="850" swimtime="00:11:00.33" />
                    <SPLIT distance="900" swimtime="00:11:39.78" />
                    <SPLIT distance="950" swimtime="00:12:19.14" />
                    <SPLIT distance="1000" swimtime="00:12:58.39" />
                    <SPLIT distance="1050" swimtime="00:13:37.40" />
                    <SPLIT distance="1100" swimtime="00:14:16.81" />
                    <SPLIT distance="1150" swimtime="00:14:56.42" />
                    <SPLIT distance="1200" swimtime="00:15:36.45" />
                    <SPLIT distance="1250" swimtime="00:16:15.82" />
                    <SPLIT distance="1300" swimtime="00:16:54.87" />
                    <SPLIT distance="1350" swimtime="00:17:33.72" />
                    <SPLIT distance="1400" swimtime="00:18:13.26" />
                    <SPLIT distance="1450" swimtime="00:18:51.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="10315">
              <RESULTS>
                <RESULT eventid="1113" points="408" reactiontime="+95" swimtime="00:02:33.62" resultid="10316" heatid="13930" lane="1" entrytime="00:02:33.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                    <SPLIT distance="150" swimtime="00:01:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="332" reactiontime="+109" swimtime="00:20:57.31" resultid="10317" heatid="13942" lane="5" entrytime="00:21:08.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:01:59.12" />
                    <SPLIT distance="200" swimtime="00:02:41.41" />
                    <SPLIT distance="250" swimtime="00:03:23.94" />
                    <SPLIT distance="300" swimtime="00:04:06.09" />
                    <SPLIT distance="350" swimtime="00:04:48.64" />
                    <SPLIT distance="400" swimtime="00:05:31.08" />
                    <SPLIT distance="450" swimtime="00:06:13.24" />
                    <SPLIT distance="500" swimtime="00:06:55.55" />
                    <SPLIT distance="550" swimtime="00:07:37.66" />
                    <SPLIT distance="600" swimtime="00:08:20.00" />
                    <SPLIT distance="650" swimtime="00:09:02.38" />
                    <SPLIT distance="700" swimtime="00:09:44.60" />
                    <SPLIT distance="750" swimtime="00:10:26.86" />
                    <SPLIT distance="800" swimtime="00:11:08.82" />
                    <SPLIT distance="850" swimtime="00:11:51.21" />
                    <SPLIT distance="900" swimtime="00:12:33.29" />
                    <SPLIT distance="950" swimtime="00:13:15.38" />
                    <SPLIT distance="1000" swimtime="00:13:57.72" />
                    <SPLIT distance="1050" swimtime="00:14:39.96" />
                    <SPLIT distance="1100" swimtime="00:15:21.93" />
                    <SPLIT distance="1150" swimtime="00:16:03.91" />
                    <SPLIT distance="1200" swimtime="00:16:46.69" />
                    <SPLIT distance="1250" swimtime="00:17:28.78" />
                    <SPLIT distance="1300" swimtime="00:18:10.95" />
                    <SPLIT distance="1350" swimtime="00:18:53.44" />
                    <SPLIT distance="1400" swimtime="00:19:35.95" />
                    <SPLIT distance="1450" swimtime="00:20:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="10318" heatid="14070" lane="1" entrytime="00:01:11.98" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="10319" heatid="14112" lane="8" entrytime="00:05:11.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-03" firstname="Katarzyna" gender="F" lastname="Nikelewska" nation="POL" athleteid="10284">
              <RESULTS>
                <RESULT eventid="1222" points="207" reactiontime="+93" swimtime="00:03:55.03" resultid="10285" heatid="13962" lane="2" entrytime="00:03:07.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:50.50" />
                    <SPLIT distance="150" swimtime="00:02:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="211" swimtime="00:01:48.01" resultid="10286" heatid="14004" lane="3" entrytime="00:01:22.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="246" reactiontime="+86" swimtime="00:00:46.99" resultid="10287" heatid="14086" lane="4" entrytime="00:00:39.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="10181">
              <RESULTS>
                <RESULT eventid="1079" points="157" reactiontime="+85" swimtime="00:00:38.70" resultid="10182" heatid="13906" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1165" points="94" reactiontime="+103" swimtime="00:31:50.50" resultid="10183" heatid="13939" lane="6" entrytime="00:31:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:44.35" />
                    <SPLIT distance="150" swimtime="00:02:43.54" />
                    <SPLIT distance="200" swimtime="00:03:44.30" />
                    <SPLIT distance="250" swimtime="00:04:46.90" />
                    <SPLIT distance="300" swimtime="00:05:50.63" />
                    <SPLIT distance="350" swimtime="00:06:51.88" />
                    <SPLIT distance="400" swimtime="00:07:54.11" />
                    <SPLIT distance="450" swimtime="00:08:56.57" />
                    <SPLIT distance="500" swimtime="00:10:00.29" />
                    <SPLIT distance="550" swimtime="00:11:03.78" />
                    <SPLIT distance="600" swimtime="00:12:07.86" />
                    <SPLIT distance="650" swimtime="00:13:12.97" />
                    <SPLIT distance="700" swimtime="00:14:17.89" />
                    <SPLIT distance="750" swimtime="00:15:23.02" />
                    <SPLIT distance="800" swimtime="00:16:29.24" />
                    <SPLIT distance="850" swimtime="00:17:32.47" />
                    <SPLIT distance="900" swimtime="00:18:37.69" />
                    <SPLIT distance="950" swimtime="00:19:43.12" />
                    <SPLIT distance="1000" swimtime="00:20:49.00" />
                    <SPLIT distance="1050" swimtime="00:21:54.81" />
                    <SPLIT distance="1100" swimtime="00:23:00.92" />
                    <SPLIT distance="1150" swimtime="00:24:06.51" />
                    <SPLIT distance="1200" swimtime="00:25:13.81" />
                    <SPLIT distance="1250" swimtime="00:26:20.70" />
                    <SPLIT distance="1300" swimtime="00:27:28.11" />
                    <SPLIT distance="1350" swimtime="00:28:34.88" />
                    <SPLIT distance="1400" swimtime="00:29:42.79" />
                    <SPLIT distance="1450" swimtime="00:30:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="107" reactiontime="+67" swimtime="00:00:50.52" resultid="10184" heatid="13951" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1273" points="149" reactiontime="+87" swimtime="00:01:28.34" resultid="10185" heatid="13979" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="100" reactiontime="+83" swimtime="00:01:51.89" resultid="10186" heatid="14033" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="124" reactiontime="+101" swimtime="00:03:24.47" resultid="10187" heatid="14046" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:34.88" />
                    <SPLIT distance="150" swimtime="00:02:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="90" reactiontime="+77" swimtime="00:04:09.11" resultid="10188" heatid="14078" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:02:00.31" />
                    <SPLIT distance="150" swimtime="00:03:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="111" reactiontime="+87" swimtime="00:07:36.88" resultid="10189" heatid="14106" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                    <SPLIT distance="100" swimtime="00:01:42.30" />
                    <SPLIT distance="150" swimtime="00:02:39.61" />
                    <SPLIT distance="200" swimtime="00:03:39.42" />
                    <SPLIT distance="250" swimtime="00:04:39.28" />
                    <SPLIT distance="300" swimtime="00:05:39.76" />
                    <SPLIT distance="350" swimtime="00:06:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="10190">
              <RESULTS>
                <RESULT eventid="1273" points="495" reactiontime="+77" swimtime="00:00:59.28" resultid="10191" heatid="13987" lane="7" entrytime="00:00:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="457" reactiontime="+79" swimtime="00:02:12.41" resultid="10192" heatid="14052" lane="6" entrytime="00:02:11.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1744" points="437" swimtime="00:04:49.84" resultid="10193" heatid="14113" lane="6" entrytime="00:04:53.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:47.96" />
                    <SPLIT distance="200" swimtime="00:02:25.59" />
                    <SPLIT distance="250" swimtime="00:03:02.45" />
                    <SPLIT distance="300" swimtime="00:03:39.19" />
                    <SPLIT distance="350" swimtime="00:04:15.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="10354">
              <RESULTS>
                <RESULT eventid="1273" points="523" reactiontime="+71" swimtime="00:00:58.19" resultid="10355" heatid="13988" lane="4" entrytime="00:00:57.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="507" reactiontime="+84" swimtime="00:02:07.91" resultid="10356" heatid="14053" lane="1" entrytime="00:02:08.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="431" reactiontime="+80" swimtime="00:04:51.27" resultid="10357" heatid="14114" lane="1" entrytime="00:04:38.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                    <SPLIT distance="200" swimtime="00:02:22.17" />
                    <SPLIT distance="250" swimtime="00:02:59.96" />
                    <SPLIT distance="300" swimtime="00:03:37.33" />
                    <SPLIT distance="350" swimtime="00:04:14.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="10194">
              <RESULTS>
                <RESULT eventid="1239" points="427" reactiontime="+76" swimtime="00:02:48.64" resultid="10195" heatid="13969" lane="5" entrytime="00:02:49.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="462" swimtime="00:01:14.92" resultid="10196" heatid="14012" lane="6" entrytime="00:01:16.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="391" reactiontime="+82" swimtime="00:02:19.44" resultid="10197" heatid="14051" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10198" heatid="14097" lane="2" entrytime="00:00:33.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="10280">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="10281" heatid="13969" lane="9" entrytime="00:02:54.50" />
                <RESULT eventid="1406" points="421" reactiontime="+87" swimtime="00:01:17.22" resultid="10282" heatid="14012" lane="0" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="444" reactiontime="+87" swimtime="00:00:34.63" resultid="10283" heatid="14098" lane="0" entrytime="00:00:32.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="10350">
              <RESULTS>
                <RESULT eventid="1239" points="454" reactiontime="+91" swimtime="00:02:45.19" resultid="10351" heatid="13970" lane="0" entrytime="00:02:46.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="544" reactiontime="+89" swimtime="00:01:10.91" resultid="10352" heatid="14013" lane="2" entrytime="00:01:12.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="555" reactiontime="+80" swimtime="00:00:32.13" resultid="10353" heatid="14098" lane="8" entrytime="00:00:31.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="10219">
              <RESULTS>
                <RESULT eventid="1079" points="401" reactiontime="+86" swimtime="00:00:28.35" resultid="10220" heatid="13911" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="372" swimtime="00:02:38.37" resultid="10221" heatid="13929" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="368" reactiontime="+76" swimtime="00:00:33.54" resultid="10222" heatid="13957" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="419" reactiontime="+88" swimtime="00:01:02.65" resultid="10223" heatid="13984" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="381" reactiontime="+80" swimtime="00:01:11.64" resultid="10224" heatid="14038" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="376" reactiontime="+89" swimtime="00:02:21.32" resultid="10225" heatid="14051" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="342" reactiontime="+83" swimtime="00:02:39.94" resultid="10226" heatid="14081" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:01:59.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="10227">
              <RESULTS>
                <RESULT eventid="1079" points="451" reactiontime="+76" swimtime="00:00:27.26" resultid="10228" heatid="13912" lane="5" entrytime="00:00:28.05" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 10:18)" eventid="1239" reactiontime="+84" status="DSQ" swimtime="00:02:55.04" resultid="10229" heatid="13965" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:01:23.56" />
                    <SPLIT distance="150" swimtime="00:02:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="437" swimtime="00:01:01.78" resultid="10230" heatid="13987" lane="9" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="383" reactiontime="+88" swimtime="00:01:19.70" resultid="10231" heatid="14012" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="421" reactiontime="+80" swimtime="00:00:29.91" resultid="10232" heatid="14025" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1681" points="434" reactiontime="+76" swimtime="00:00:34.87" resultid="10233" heatid="14095" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-17" firstname="Waldemar" gender="M" lastname="de Makay" nation="POL" athleteid="10248">
              <RESULTS>
                <RESULT eventid="1079" points="254" reactiontime="+107" swimtime="00:00:33.00" resultid="10249" heatid="13908" lane="8" entrytime="00:00:33.00" />
                <RESULT comment="Rekord Polski" eventid="1165" points="267" reactiontime="+111" swimtime="00:22:31.71" resultid="10250" heatid="13941" lane="7" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="150" swimtime="00:02:10.00" />
                    <SPLIT distance="200" swimtime="00:02:55.82" />
                    <SPLIT distance="250" swimtime="00:03:41.75" />
                    <SPLIT distance="300" swimtime="00:04:27.99" />
                    <SPLIT distance="350" swimtime="00:05:13.95" />
                    <SPLIT distance="400" swimtime="00:06:00.04" />
                    <SPLIT distance="450" swimtime="00:06:45.34" />
                    <SPLIT distance="500" swimtime="00:07:31.11" />
                    <SPLIT distance="550" swimtime="00:08:16.75" />
                    <SPLIT distance="600" swimtime="00:09:02.53" />
                    <SPLIT distance="650" swimtime="00:09:48.34" />
                    <SPLIT distance="700" swimtime="00:10:34.20" />
                    <SPLIT distance="750" swimtime="00:11:19.26" />
                    <SPLIT distance="800" swimtime="00:12:04.27" />
                    <SPLIT distance="850" swimtime="00:12:48.75" />
                    <SPLIT distance="900" swimtime="00:13:34.09" />
                    <SPLIT distance="950" swimtime="00:14:19.90" />
                    <SPLIT distance="1000" swimtime="00:15:05.53" />
                    <SPLIT distance="1050" swimtime="00:15:50.43" />
                    <SPLIT distance="1100" swimtime="00:16:36.03" />
                    <SPLIT distance="1150" swimtime="00:17:20.81" />
                    <SPLIT distance="1200" swimtime="00:18:06.24" />
                    <SPLIT distance="1250" swimtime="00:18:50.55" />
                    <SPLIT distance="1300" swimtime="00:19:36.16" />
                    <SPLIT distance="1350" swimtime="00:20:20.76" />
                    <SPLIT distance="1400" swimtime="00:21:05.72" />
                    <SPLIT distance="1450" swimtime="00:21:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="180" reactiontime="+72" swimtime="00:00:42.57" resultid="10251" heatid="13952" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1273" points="262" reactiontime="+118" swimtime="00:01:13.22" resultid="10252" heatid="13981" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="178" reactiontime="+73" swimtime="00:01:32.17" resultid="10253" heatid="14034" lane="8" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="243" reactiontime="+116" swimtime="00:02:43.44" resultid="10254" heatid="14049" lane="1" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="161" reactiontime="+80" swimtime="00:03:25.45" resultid="10255" heatid="14079" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                    <SPLIT distance="100" swimtime="00:01:40.07" />
                    <SPLIT distance="150" swimtime="00:02:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="259" swimtime="00:05:45.21" resultid="10256" heatid="14111" lane="9" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                    <SPLIT distance="200" swimtime="00:02:50.38" />
                    <SPLIT distance="250" swimtime="00:03:34.65" />
                    <SPLIT distance="300" swimtime="00:04:19.50" />
                    <SPLIT distance="350" swimtime="00:05:03.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="10199">
              <RESULTS>
                <RESULT eventid="1165" points="359" reactiontime="+79" swimtime="00:20:25.52" resultid="10200" heatid="13942" lane="8" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="150" swimtime="00:01:55.79" />
                    <SPLIT distance="200" swimtime="00:02:36.29" />
                    <SPLIT distance="250" swimtime="00:03:17.32" />
                    <SPLIT distance="300" swimtime="00:03:58.59" />
                    <SPLIT distance="350" swimtime="00:04:39.58" />
                    <SPLIT distance="400" swimtime="00:05:20.85" />
                    <SPLIT distance="450" swimtime="00:06:02.17" />
                    <SPLIT distance="500" swimtime="00:06:43.91" />
                    <SPLIT distance="550" swimtime="00:07:24.89" />
                    <SPLIT distance="600" swimtime="00:08:06.23" />
                    <SPLIT distance="650" swimtime="00:08:47.56" />
                    <SPLIT distance="700" swimtime="00:09:29.26" />
                    <SPLIT distance="750" swimtime="00:10:10.46" />
                    <SPLIT distance="800" swimtime="00:10:51.85" />
                    <SPLIT distance="850" swimtime="00:11:33.29" />
                    <SPLIT distance="900" swimtime="00:12:15.17" />
                    <SPLIT distance="950" swimtime="00:12:57.33" />
                    <SPLIT distance="1000" swimtime="00:13:38.74" />
                    <SPLIT distance="1050" swimtime="00:14:19.98" />
                    <SPLIT distance="1100" swimtime="00:15:01.88" />
                    <SPLIT distance="1150" swimtime="00:15:43.08" />
                    <SPLIT distance="1200" swimtime="00:16:24.71" />
                    <SPLIT distance="1250" swimtime="00:17:06.57" />
                    <SPLIT distance="1300" swimtime="00:17:47.39" />
                    <SPLIT distance="1350" swimtime="00:18:28.69" />
                    <SPLIT distance="1400" swimtime="00:19:08.95" />
                    <SPLIT distance="1450" swimtime="00:19:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="385" reactiontime="+81" swimtime="00:01:04.44" resultid="10201" heatid="13983" lane="6" entrytime="00:01:06.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="328" reactiontime="+92" swimtime="00:00:32.51" resultid="10202" heatid="14023" lane="2" entrytime="00:00:32.33" />
                <RESULT eventid="1508" points="363" reactiontime="+87" swimtime="00:02:22.95" resultid="10203" heatid="14050" lane="8" entrytime="00:02:27.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="383" reactiontime="+80" swimtime="00:05:02.96" resultid="10204" heatid="14111" lane="4" entrytime="00:05:18.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:48.25" />
                    <SPLIT distance="200" swimtime="00:02:27.65" />
                    <SPLIT distance="250" swimtime="00:03:06.62" />
                    <SPLIT distance="300" swimtime="00:03:46.50" />
                    <SPLIT distance="350" swimtime="00:04:26.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-18" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="10288">
              <RESULTS>
                <RESULT eventid="1062" points="234" reactiontime="+104" swimtime="00:00:38.48" resultid="10289" heatid="13898" lane="2" entrytime="00:00:39.69" />
                <RESULT eventid="1187" points="187" reactiontime="+81" swimtime="00:00:47.31" resultid="10290" heatid="13945" lane="3" entrytime="00:00:47.73" />
                <RESULT eventid="1256" points="140" reactiontime="+121" swimtime="00:01:40.07" resultid="10291" heatid="13971" lane="3" entrytime="00:01:40.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="144" reactiontime="+88" swimtime="00:01:50.66" resultid="10292" heatid="14029" lane="2" entrytime="00:01:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="133" reactiontime="+77" swimtime="00:04:02.59" resultid="10293" heatid="14072" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.47" />
                    <SPLIT distance="150" swimtime="00:03:01.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="10257">
              <RESULTS>
                <RESULT eventid="1256" points="222" reactiontime="+105" swimtime="00:01:25.96" resultid="10258" heatid="13973" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="222" reactiontime="+91" swimtime="00:01:35.93" resultid="10259" heatid="14030" lane="9" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="205" reactiontime="+100" swimtime="00:03:11.30" resultid="10260" heatid="14040" lane="3" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                    <SPLIT distance="150" swimtime="00:02:22.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="226" reactiontime="+106" swimtime="00:03:23.43" resultid="10261" heatid="14074" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:39.49" />
                    <SPLIT distance="150" swimtime="00:02:32.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="10262">
              <RESULTS>
                <RESULT eventid="1079" points="180" reactiontime="+114" swimtime="00:00:37.03" resultid="10263" heatid="13906" lane="3" entrytime="00:00:36.84" />
                <RESULT eventid="1239" points="228" reactiontime="+120" swimtime="00:03:27.82" resultid="10264" heatid="13966" lane="2" entrytime="00:03:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                    <SPLIT distance="100" swimtime="00:01:40.81" />
                    <SPLIT distance="150" swimtime="00:02:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="220" swimtime="00:01:35.82" resultid="10265" heatid="14007" lane="6" entrytime="00:01:36.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="145" swimtime="00:07:43.58" resultid="10266" heatid="14060" lane="9" entrytime="00:07:44.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:45.26" />
                    <SPLIT distance="150" swimtime="00:02:54.66" />
                    <SPLIT distance="200" swimtime="00:04:04.88" />
                    <SPLIT distance="250" swimtime="00:04:58.04" />
                    <SPLIT distance="300" swimtime="00:05:55.43" />
                    <SPLIT distance="350" swimtime="00:06:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="125" swimtime="00:01:39.55" resultid="10267" heatid="14067" lane="6" entrytime="00:01:36.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="219" swimtime="00:00:43.78" resultid="10268" heatid="14091" lane="6" entrytime="00:00:43.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="10326">
              <RESULTS>
                <RESULT eventid="1165" points="308" reactiontime="+86" swimtime="00:21:29.56" resultid="10327" heatid="13942" lane="0" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:02:36.04" />
                    <SPLIT distance="250" swimtime="00:03:18.07" />
                    <SPLIT distance="300" swimtime="00:04:00.18" />
                    <SPLIT distance="350" swimtime="00:04:42.15" />
                    <SPLIT distance="400" swimtime="00:05:25.19" />
                    <SPLIT distance="450" swimtime="00:06:08.11" />
                    <SPLIT distance="500" swimtime="00:06:51.38" />
                    <SPLIT distance="550" swimtime="00:07:34.65" />
                    <SPLIT distance="600" swimtime="00:08:18.26" />
                    <SPLIT distance="650" swimtime="00:09:02.17" />
                    <SPLIT distance="700" swimtime="00:09:46.39" />
                    <SPLIT distance="750" swimtime="00:10:30.30" />
                    <SPLIT distance="800" swimtime="00:11:14.86" />
                    <SPLIT distance="850" swimtime="00:11:58.67" />
                    <SPLIT distance="900" swimtime="00:12:43.04" />
                    <SPLIT distance="950" swimtime="00:14:55.62" />
                    <SPLIT distance="1000" swimtime="00:14:12.35" />
                    <SPLIT distance="1050" swimtime="00:16:24.13" />
                    <SPLIT distance="1100" swimtime="00:15:40.18" />
                    <SPLIT distance="1150" swimtime="00:19:23.02" />
                    <SPLIT distance="1200" swimtime="00:17:09.14" />
                    <SPLIT distance="1250" swimtime="00:20:49.74" />
                    <SPLIT distance="1300" swimtime="00:18:38.59" />
                    <SPLIT distance="1400" swimtime="00:20:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="397" reactiontime="+81" swimtime="00:01:03.78" resultid="10328" heatid="13985" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="334" reactiontime="+97" swimtime="00:01:23.43" resultid="10329" heatid="14009" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="369" reactiontime="+83" swimtime="00:02:22.11" resultid="10330" heatid="14050" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="340" swimtime="00:00:37.83" resultid="10331" heatid="14095" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="10205">
              <RESULTS>
                <RESULT eventid="1113" points="310" reactiontime="+104" swimtime="00:02:48.36" resultid="10206" heatid="13927" lane="3" entrytime="00:02:48.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="370" reactiontime="+94" swimtime="00:01:05.30" resultid="10207" heatid="13983" lane="0" entrytime="00:01:07.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="313" reactiontime="+73" swimtime="00:01:16.49" resultid="10208" heatid="14036" lane="8" entrytime="00:01:17.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="312" reactiontime="+71" swimtime="00:02:44.85" resultid="10209" heatid="14080" lane="5" entrytime="00:02:47.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="150" swimtime="00:02:02.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="10234">
              <RESULTS>
                <RESULT eventid="1079" points="141" reactiontime="+111" swimtime="00:00:40.09" resultid="10235" heatid="13905" lane="4" entrytime="00:00:39.60" />
                <RESULT comment="Przekroczony regulaminowy limit czasu." eventid="1165" reactiontime="+114" status="OTL" swimtime="00:27:23.17" resultid="10236" heatid="13940" lane="8" entrytime="00:26:29.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:33.50" />
                    <SPLIT distance="200" swimtime="00:03:28.62" />
                    <SPLIT distance="250" swimtime="00:04:24.90" />
                    <SPLIT distance="300" swimtime="00:05:19.98" />
                    <SPLIT distance="350" swimtime="00:06:16.25" />
                    <SPLIT distance="400" swimtime="00:07:12.06" />
                    <SPLIT distance="450" swimtime="00:08:07.40" />
                    <SPLIT distance="500" swimtime="00:09:01.91" />
                    <SPLIT distance="550" swimtime="00:09:56.97" />
                    <SPLIT distance="600" swimtime="00:10:51.33" />
                    <SPLIT distance="650" swimtime="00:11:46.07" />
                    <SPLIT distance="700" swimtime="00:12:41.59" />
                    <SPLIT distance="750" swimtime="00:13:36.99" />
                    <SPLIT distance="800" swimtime="00:14:32.32" />
                    <SPLIT distance="850" swimtime="00:15:27.54" />
                    <SPLIT distance="900" swimtime="00:16:23.16" />
                    <SPLIT distance="950" swimtime="00:17:18.50" />
                    <SPLIT distance="1000" swimtime="00:18:13.60" />
                    <SPLIT distance="1050" swimtime="00:19:09.26" />
                    <SPLIT distance="1100" swimtime="00:20:05.06" />
                    <SPLIT distance="1150" swimtime="00:22:52.97" />
                    <SPLIT distance="1200" swimtime="00:21:56.96" />
                    <SPLIT distance="1250" swimtime="00:24:44.29" />
                    <SPLIT distance="1300" swimtime="00:23:49.34" />
                    <SPLIT distance="1350" swimtime="00:26:33.19" />
                    <SPLIT distance="1400" swimtime="00:25:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="74" reactiontime="+86" swimtime="00:00:57.04" resultid="10237" heatid="13950" lane="6" entrytime="00:00:56.21" />
                <RESULT eventid="1273" points="138" reactiontime="+118" swimtime="00:01:30.68" resultid="10238" heatid="13979" lane="2" entrytime="00:01:28.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="140" reactiontime="+117" swimtime="00:03:16.33" resultid="10239" heatid="14046" lane="2" entrytime="00:03:13.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="100" swimtime="00:01:35.82" />
                    <SPLIT distance="150" swimtime="00:02:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="74" reactiontime="+120" swimtime="00:01:58.22" resultid="10240" heatid="14066" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="152" reactiontime="+112" swimtime="00:06:51.74" resultid="10241" heatid="14108" lane="8" entrytime="00:06:48.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="150" swimtime="00:02:31.75" />
                    <SPLIT distance="250" swimtime="00:04:19.33" />
                    <SPLIT distance="300" swimtime="00:05:12.54" />
                    <SPLIT distance="350" swimtime="00:06:03.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-10" firstname="Anna" gender="F" lastname="Turczyn" nation="POL" athleteid="10310">
              <RESULTS>
                <RESULT eventid="1096" points="139" reactiontime="+110" swimtime="00:04:03.29" resultid="10311" heatid="13918" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.41" />
                    <SPLIT distance="100" swimtime="00:02:05.78" />
                    <SPLIT distance="150" swimtime="00:03:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="198" reactiontime="+134" swimtime="00:03:58.55" resultid="10312" heatid="13960" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.30" />
                    <SPLIT distance="100" swimtime="00:01:53.48" />
                    <SPLIT distance="150" swimtime="00:02:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="209" reactiontime="+101" swimtime="00:01:48.43" resultid="10313" heatid="14002" lane="9" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="10314" heatid="14084" lane="6" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="10300">
              <RESULTS>
                <RESULT eventid="1113" points="419" reactiontime="+71" swimtime="00:02:32.29" resultid="10301" heatid="13930" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="489" reactiontime="+72" swimtime="00:02:41.19" resultid="10303" heatid="13970" lane="7" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:01:58.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="449" reactiontime="+78" swimtime="00:01:15.60" resultid="10304" heatid="14013" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="10269">
              <RESULTS>
                <RESULT eventid="1079" points="234" reactiontime="+83" swimtime="00:00:33.89" resultid="10270" heatid="13909" lane="5" entrytime="00:00:31.20" />
                <RESULT eventid="1205" points="168" reactiontime="+71" swimtime="00:00:43.52" resultid="10271" heatid="13953" lane="9" entrytime="00:00:40.86" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="10272" heatid="13981" lane="7" entrytime="00:01:12.11" />
                <RESULT eventid="1406" points="231" reactiontime="+91" swimtime="00:01:34.33" resultid="10273" heatid="14008" lane="6" entrytime="00:01:29.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="10274" heatid="14047" lane="2" entrytime="00:02:54.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="10332">
              <RESULTS>
                <RESULT eventid="1147" points="107" reactiontime="+98" swimtime="00:17:06.07" resultid="10333" heatid="13935" lane="6" entrytime="00:17:05.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.34" />
                    <SPLIT distance="100" swimtime="00:01:58.53" />
                    <SPLIT distance="150" swimtime="00:03:04.78" />
                    <SPLIT distance="200" swimtime="00:04:09.43" />
                    <SPLIT distance="250" swimtime="00:05:15.04" />
                    <SPLIT distance="300" swimtime="00:06:19.98" />
                    <SPLIT distance="350" swimtime="00:07:25.58" />
                    <SPLIT distance="400" swimtime="00:08:30.74" />
                    <SPLIT distance="450" swimtime="00:09:36.97" />
                    <SPLIT distance="500" swimtime="00:10:41.63" />
                    <SPLIT distance="550" swimtime="00:11:45.75" />
                    <SPLIT distance="600" swimtime="00:12:51.03" />
                    <SPLIT distance="650" swimtime="00:13:55.24" />
                    <SPLIT distance="700" swimtime="00:15:00.71" />
                    <SPLIT distance="750" swimtime="00:16:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="10334" heatid="13971" lane="1" entrytime="00:01:55.00" />
                <RESULT eventid="1491" points="91" reactiontime="+98" swimtime="00:04:10.97" resultid="10335" heatid="14039" lane="2" entrytime="00:04:12.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.19" />
                    <SPLIT distance="100" swimtime="00:02:00.54" />
                    <SPLIT distance="150" swimtime="00:03:09.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="95" reactiontime="+104" swimtime="00:08:41.55" resultid="10336" heatid="14102" lane="5" entrytime="00:07:22.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                    <SPLIT distance="100" swimtime="00:02:03.38" />
                    <SPLIT distance="150" swimtime="00:03:12.61" />
                    <SPLIT distance="200" swimtime="00:04:20.67" />
                    <SPLIT distance="250" swimtime="00:05:27.40" />
                    <SPLIT distance="300" swimtime="00:06:34.58" />
                    <SPLIT distance="350" swimtime="00:07:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="10242">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1222" points="373" reactiontime="+83" swimtime="00:03:13.18" resultid="10243" heatid="13962" lane="1" entrytime="00:03:14.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:02:24.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="359" swimtime="00:01:30.51" resultid="10244" heatid="14003" lane="3" entrytime="00:01:30.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="285" reactiontime="+82" swimtime="00:02:51.51" resultid="10245" heatid="14041" lane="1" entrytime="00:02:52.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:09.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="355" reactiontime="+80" swimtime="00:00:41.63" resultid="10246" heatid="14086" lane="1" entrytime="00:00:41.41" />
                <RESULT eventid="1721" points="284" swimtime="00:06:02.36" resultid="10247" heatid="14104" lane="3" entrytime="00:05:54.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:02:15.88" />
                    <SPLIT distance="200" swimtime="00:03:03.03" />
                    <SPLIT distance="250" swimtime="00:03:47.27" />
                    <SPLIT distance="300" swimtime="00:04:32.87" />
                    <SPLIT distance="350" swimtime="00:05:19.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-11" firstname="Bolesław" gender="M" lastname="Szuter" nation="POL" athleteid="10178">
              <RESULTS>
                <RESULT eventid="1273" points="595" reactiontime="+82" swimtime="00:00:55.75" resultid="10179" heatid="13989" lane="7" entrytime="00:00:56.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1508" points="540" reactiontime="+89" swimtime="00:02:05.18" resultid="10180" heatid="14053" lane="2" entrytime="00:02:06.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="150" swimtime="00:01:33.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="10346">
              <RESULTS>
                <RESULT eventid="1079" points="562" reactiontime="+73" swimtime="00:00:25.33" resultid="10347" heatid="13917" lane="6" entrytime="00:00:24.96" />
                <RESULT eventid="1205" points="558" reactiontime="+72" swimtime="00:00:29.19" resultid="10348" heatid="13958" lane="6" entrytime="00:00:29.13" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="10349" heatid="14027" lane="2" entrytime="00:00:27.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="10294">
              <RESULTS>
                <RESULT eventid="1079" points="528" reactiontime="+72" swimtime="00:00:25.86" resultid="10295" heatid="13917" lane="8" entrytime="00:00:25.60" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="10296" heatid="13977" lane="8" />
                <RESULT eventid="1440" points="590" reactiontime="+73" swimtime="00:00:26.74" resultid="10297" heatid="14027" lane="3" entrytime="00:00:26.80" />
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 20:20), Z-2" eventid="1578" reactiontime="+78" status="DSQ" swimtime="00:05:29.66" resultid="10298" heatid="14062" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:34.79" />
                    <SPLIT distance="250" swimtime="00:03:23.17" />
                    <SPLIT distance="300" swimtime="00:04:11.87" />
                    <SPLIT distance="350" swimtime="00:04:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="495" swimtime="00:01:02.96" resultid="10299" heatid="14071" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="10305">
              <RESULTS>
                <RESULT eventid="1256" points="276" reactiontime="+89" swimtime="00:01:19.91" resultid="10306" heatid="13974" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="245" reactiontime="+91" swimtime="00:00:39.00" resultid="10307" heatid="14016" lane="0" entrytime="00:00:38.50" />
                <RESULT eventid="1491" points="246" reactiontime="+96" swimtime="00:03:00.08" resultid="10308" heatid="14042" lane="8" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:27.32" />
                    <SPLIT distance="150" swimtime="00:02:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="247" reactiontime="+82" swimtime="00:06:19.49" resultid="10309" heatid="14103" lane="3" entrytime="00:06:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:30.07" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                    <SPLIT distance="200" swimtime="00:03:07.57" />
                    <SPLIT distance="250" swimtime="00:03:57.13" />
                    <SPLIT distance="300" swimtime="00:04:46.04" />
                    <SPLIT distance="350" swimtime="00:05:34.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="456" reactiontime="+79" swimtime="00:02:01.37" resultid="10360" heatid="13999" lane="3" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:06.43" />
                    <SPLIT distance="150" swimtime="00:01:36.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10219" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="10280" number="2" />
                    <RELAYPOSITION athleteid="10300" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="10178" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="542" reactiontime="+78" swimtime="00:01:54.56" resultid="10361" heatid="13999" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="100" swimtime="00:01:00.85" />
                    <SPLIT distance="150" swimtime="00:01:28.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10346" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="10350" number="2" />
                    <RELAYPOSITION athleteid="10354" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="10194" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1548" points="561" reactiontime="+73" swimtime="00:01:42.84" resultid="10363" heatid="14056" lane="5" entrytime="00:01:44.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.45" />
                    <SPLIT distance="100" swimtime="00:00:51.36" />
                    <SPLIT distance="150" swimtime="00:01:16.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10294" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="10194" number="2" />
                    <RELAYPOSITION athleteid="10178" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="10354" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1548" points="386" reactiontime="+91" swimtime="00:01:56.49" resultid="10366" heatid="14056" lane="7" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:00:58.19" />
                    <SPLIT distance="150" swimtime="00:01:27.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10210" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="10350" number="2" />
                    <RELAYPOSITION athleteid="10199" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="10326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="1358" points="280" reactiontime="+76" swimtime="00:02:42.38" resultid="10362" heatid="13996" lane="1" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:05.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10257" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="10275" number="2" />
                    <RELAYPOSITION athleteid="10305" number="3" reactiontime="+86" />
                    <RELAYPOSITION athleteid="10341" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="7">
              <RESULTS>
                <RESULT eventid="1525" points="281" reactiontime="+77" swimtime="00:02:27.47" resultid="10364" heatid="14054" lane="1" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10275" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="10288" number="2" />
                    <RELAYPOSITION athleteid="10257" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="10305" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="325" reactiontime="+81" swimtime="00:02:03.39" resultid="10358" heatid="13934" lane="7" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="150" swimtime="00:01:35.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10346" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="10275" number="2" />
                    <RELAYPOSITION athleteid="10341" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="10300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="238" swimtime="00:02:16.77" resultid="10359" heatid="13934" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10294" number="1" />
                    <RELAYPOSITION athleteid="10257" number="2" />
                    <RELAYPOSITION athleteid="10310" number="3" />
                    <RELAYPOSITION athleteid="10210" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1698" points="338" reactiontime="+75" swimtime="00:02:14.07" resultid="10365" heatid="14101" lane="6" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:39.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10354" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="10275" number="2" />
                    <RELAYPOSITION athleteid="10294" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="10305" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="10694" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁPODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="502611200008" athleteid="10718">
              <RESULTS>
                <RESULT eventid="1079" points="287" reactiontime="+92" swimtime="00:00:31.68" resultid="10719" heatid="13910" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1205" points="213" reactiontime="+67" swimtime="00:00:40.22" resultid="10720" heatid="13954" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1474" points="198" reactiontime="+71" swimtime="00:01:29.09" resultid="10721" heatid="14035" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="10722" heatid="14079" lane="2" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611" athleteid="10702">
              <RESULTS>
                <RESULT eventid="1239" points="197" swimtime="00:03:38.21" resultid="10703" heatid="13966" lane="9" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:46.92" />
                    <SPLIT distance="150" swimtime="00:02:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1406" points="189" reactiontime="+99" swimtime="00:01:40.76" resultid="10704" heatid="14007" lane="0" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="10723">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="10724" heatid="13897" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="10725" heatid="13972" lane="7" entrytime="00:01:35.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="10726" heatid="14039" lane="6" entrytime="00:03:40.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="10727" heatid="14073" lane="6" entrytime="00:04:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" license="502611200001" athleteid="10711">
              <RESULTS>
                <RESULT eventid="1079" points="318" reactiontime="+89" swimtime="00:00:30.61" resultid="10712" heatid="13911" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1341" points="225" swimtime="00:03:03.31" resultid="10713" heatid="13995" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:01:27.18" />
                    <SPLIT distance="150" swimtime="00:02:15.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="333" reactiontime="+88" swimtime="00:00:32.36" resultid="10714" heatid="14022" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1613" points="285" swimtime="00:01:15.67" resultid="10715" heatid="14070" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="10728">
              <RESULTS>
                <RESULT eventid="1147" points="446" reactiontime="+81" swimtime="00:10:37.72" resultid="10729" heatid="13937" lane="3" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:01:54.02" />
                    <SPLIT distance="200" swimtime="00:02:34.11" />
                    <SPLIT distance="250" swimtime="00:03:13.83" />
                    <SPLIT distance="300" swimtime="00:03:54.04" />
                    <SPLIT distance="350" swimtime="00:04:34.17" />
                    <SPLIT distance="400" swimtime="00:05:14.40" />
                    <SPLIT distance="450" swimtime="00:05:54.53" />
                    <SPLIT distance="500" swimtime="00:06:35.26" />
                    <SPLIT distance="550" swimtime="00:07:15.45" />
                    <SPLIT distance="600" swimtime="00:07:56.11" />
                    <SPLIT distance="650" swimtime="00:08:36.28" />
                    <SPLIT distance="700" swimtime="00:09:17.58" />
                    <SPLIT distance="750" swimtime="00:09:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1222" points="427" reactiontime="+84" swimtime="00:03:04.71" resultid="10730" heatid="13962" lane="3" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1388" points="446" reactiontime="+93" swimtime="00:01:24.17" resultid="10731" heatid="14004" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="440" reactiontime="+88" swimtime="00:02:28.49" resultid="10732" heatid="14043" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="427" swimtime="00:00:39.12" resultid="10733" heatid="14087" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1721" points="442" reactiontime="+74" swimtime="00:05:12.75" resultid="10734" heatid="14105" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:52.78" />
                    <SPLIT distance="200" swimtime="00:02:33.20" />
                    <SPLIT distance="250" swimtime="00:03:13.42" />
                    <SPLIT distance="300" swimtime="00:03:54.28" />
                    <SPLIT distance="350" swimtime="00:04:34.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="12310">
              <RESULTS>
                <RESULT eventid="1388" points="103" reactiontime="+103" swimtime="00:02:16.91" resultid="12311" heatid="14000" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="123" reactiontime="+105" swimtime="00:00:59.26" resultid="12312" heatid="14083" lane="0" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-04" firstname="Szanli" gender="M" lastname="Ulasz" nation="POL" license="502611200015" athleteid="10708">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:23)" eventid="1079" reactiontime="+67" status="DSQ" swimtime="00:00:36.08" resultid="10709" heatid="13906" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1681" points="180" reactiontime="+114" swimtime="00:00:46.77" resultid="10710" heatid="14091" lane="0" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="10705">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1222" points="188" reactiontime="+111" swimtime="00:04:02.65" resultid="10706" heatid="13960" lane="1" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.22" />
                    <SPLIT distance="100" swimtime="00:01:57.38" />
                    <SPLIT distance="150" swimtime="00:03:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="188" reactiontime="+105" swimtime="00:01:52.32" resultid="10707" heatid="14001" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-27" firstname="Danuta" gender="F" lastname="Skorupa" nation="POL" athleteid="10716">
              <RESULTS>
                <RESULT eventid="1187" points="78" reactiontime="+82" swimtime="00:01:03.16" resultid="10717" heatid="13944" lane="3" entrytime="00:00:59.65" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12000" name="Wks Śląsk Wrocław">
          <CONTACT email="murtacha68@gmail.com" name="Marta Frank" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="12244">
              <RESULTS>
                <RESULT eventid="1062" points="227" swimtime="00:00:38.90" resultid="12245" heatid="13899" lane="9" entrytime="00:00:37.10" />
                <RESULT eventid="1096" points="180" reactiontime="+87" swimtime="00:03:43.11" resultid="12246" heatid="13919" lane="4" entrytime="00:03:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.05" />
                    <SPLIT distance="100" swimtime="00:01:51.63" />
                    <SPLIT distance="150" swimtime="00:02:52.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="171" reactiontime="+84" swimtime="00:00:48.70" resultid="12247" heatid="13945" lane="5" entrytime="00:00:47.20" />
                <RESULT eventid="1256" points="231" reactiontime="+89" swimtime="00:01:24.79" resultid="12248" heatid="13972" lane="5" entrytime="00:01:30.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="210" reactiontime="+88" swimtime="00:01:48.20" resultid="12249" heatid="14002" lane="0" entrytime="00:01:46.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="180" reactiontime="+83" swimtime="00:03:20.07" resultid="12250" heatid="14040" lane="8" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:36.83" />
                    <SPLIT distance="150" swimtime="00:02:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="251" reactiontime="+86" swimtime="00:00:46.73" resultid="12251" heatid="14084" lane="5" entrytime="00:00:46.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-24" firstname="Tomasz" gender="M" lastname="Olas" nation="POL" athleteid="12271">
              <RESULTS>
                <RESULT eventid="1079" points="248" reactiontime="+78" swimtime="00:00:33.25" resultid="12272" heatid="13907" lane="6" entrytime="00:00:34.12" />
                <RESULT eventid="1273" points="212" reactiontime="+86" swimtime="00:01:18.63" resultid="12273" heatid="13981" lane="2" entrytime="00:01:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="231" reactiontime="+86" swimtime="00:00:36.54" resultid="12274" heatid="14020" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="12275" heatid="14048" lane="3" entrytime="00:02:42.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-13" firstname="Cezary" gender="M" lastname="Wereszczyński" nation="POL" athleteid="12276">
              <RESULTS>
                <RESULT eventid="1079" points="458" reactiontime="+75" swimtime="00:00:27.11" resultid="12277" heatid="13915" lane="7" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="345" reactiontime="+75" swimtime="00:01:06.88" resultid="12278" heatid="13986" lane="7" entrytime="00:01:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="371" reactiontime="+67" swimtime="00:00:31.20" resultid="12279" heatid="14023" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="12280" heatid="14053" lane="0" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-19" firstname="Kinga" gender="F" lastname="Murawska" nation="POL" athleteid="12252">
              <RESULTS>
                <RESULT eventid="1147" points="186" reactiontime="+95" swimtime="00:14:12.90" resultid="12253" heatid="13935" lane="3" entrytime="00:16:10.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:38.74" />
                    <SPLIT distance="150" swimtime="00:02:31.67" />
                    <SPLIT distance="200" swimtime="00:03:25.18" />
                    <SPLIT distance="250" swimtime="00:04:18.53" />
                    <SPLIT distance="300" swimtime="00:05:12.49" />
                    <SPLIT distance="350" swimtime="00:06:06.70" />
                    <SPLIT distance="400" swimtime="00:07:01.41" />
                    <SPLIT distance="450" swimtime="00:07:55.78" />
                    <SPLIT distance="500" swimtime="00:08:50.33" />
                    <SPLIT distance="550" swimtime="00:09:44.13" />
                    <SPLIT distance="600" swimtime="00:10:39.21" />
                    <SPLIT distance="650" swimtime="00:11:33.34" />
                    <SPLIT distance="700" swimtime="00:12:27.31" />
                    <SPLIT distance="750" swimtime="00:13:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="186" reactiontime="+97" swimtime="00:01:31.20" resultid="12254" heatid="13973" lane="1" entrytime="00:01:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="183" swimtime="00:01:42.37" resultid="12255" heatid="14029" lane="3" entrytime="00:01:45.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="180" swimtime="00:07:54.88" resultid="12256" heatid="14058" lane="9" entrytime="00:07:45.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                    <SPLIT distance="100" swimtime="00:01:56.78" />
                    <SPLIT distance="150" swimtime="00:02:57.60" />
                    <SPLIT distance="200" swimtime="00:03:54.56" />
                    <SPLIT distance="250" swimtime="00:04:59.83" />
                    <SPLIT distance="300" swimtime="00:06:05.76" />
                    <SPLIT distance="350" swimtime="00:07:01.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M11 - Brak dotknięcia sciany obydwoma rozłonczonymi dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 9:24)" eventid="1595" status="DSQ" swimtime="00:01:55.14" resultid="12257" heatid="14064" lane="9" entrytime="00:01:50.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="187" reactiontime="+94" swimtime="00:06:56.11" resultid="12258" heatid="14103" lane="7" entrytime="00:06:57.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                    <SPLIT distance="100" swimtime="00:01:39.63" />
                    <SPLIT distance="150" swimtime="00:02:31.92" />
                    <SPLIT distance="200" swimtime="00:03:24.70" />
                    <SPLIT distance="250" swimtime="00:04:17.88" />
                    <SPLIT distance="300" swimtime="00:05:11.77" />
                    <SPLIT distance="350" swimtime="00:06:04.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="12301">
              <RESULTS>
                <RESULT eventid="1205" points="509" reactiontime="+64" swimtime="00:00:30.09" resultid="12302" heatid="13958" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="1474" points="497" reactiontime="+65" swimtime="00:01:05.56" resultid="12303" heatid="14038" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="468" reactiontime="+64" swimtime="00:02:24.11" resultid="12304" heatid="14082" lane="6" entrytime="00:02:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:47.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-11" firstname="Głowiak" gender="F" lastname="Anna" nation="POL" athleteid="12230">
              <RESULTS>
                <RESULT eventid="1062" points="373" reactiontime="+82" swimtime="00:00:32.96" resultid="12231" heatid="13900" lane="2" entrytime="00:00:33.38" />
                <RESULT eventid="1187" points="284" reactiontime="+88" swimtime="00:00:41.12" resultid="12232" heatid="13946" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1256" points="348" reactiontime="+78" swimtime="00:01:13.97" resultid="12233" heatid="13974" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="260" reactiontime="+75" swimtime="00:01:40.81" resultid="12234" heatid="14002" lane="3" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="275" reactiontime="+95" swimtime="00:02:53.69" resultid="12235" heatid="14042" lane="1" entrytime="00:02:48.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:02:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="309" reactiontime="+78" swimtime="00:00:43.58" resultid="12236" heatid="14085" lane="7" entrytime="00:00:44.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-09-07" firstname="Radek" gender="M" lastname="Stefurak" nation="POL" athleteid="12259">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="12260" heatid="13968" lane="9" entrytime="00:03:05.00" />
                <RESULT eventid="1406" points="291" reactiontime="+85" swimtime="00:01:27.34" resultid="12261" heatid="14009" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="230" reactiontime="+77" swimtime="00:02:46.32" resultid="12262" heatid="14049" lane="8" entrytime="00:02:39.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="290" reactiontime="+85" swimtime="00:00:39.87" resultid="12263" heatid="14093" lane="5" entrytime="00:00:38.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Marta" gender="F" lastname="Frank" nation="POL" athleteid="12305">
              <RESULTS>
                <RESULT eventid="1187" points="365" reactiontime="+72" swimtime="00:00:37.84" resultid="12306" heatid="13948" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1457" points="267" reactiontime="+120" swimtime="00:01:30.24" resultid="12307" heatid="14031" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="257" reactiontime="+85" swimtime="00:01:27.44" resultid="12308" heatid="14064" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="298" reactiontime="+79" swimtime="00:03:05.72" resultid="12309" heatid="14075" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:19.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-13" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="12264">
              <RESULTS>
                <RESULT eventid="1113" points="273" reactiontime="+91" swimtime="00:02:55.63" resultid="12265" heatid="13926" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="330" reactiontime="+70" swimtime="00:00:34.76" resultid="12266" heatid="13956" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="12267" heatid="14021" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1474" points="285" reactiontime="+80" swimtime="00:01:18.87" resultid="12268" heatid="14036" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="255" reactiontime="+76" swimtime="00:02:56.35" resultid="12270" heatid="14080" lane="2" entrytime="00:02:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:02:12.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-11" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="12237">
              <RESULTS>
                <RESULT eventid="1062" points="329" reactiontime="+86" swimtime="00:00:34.35" resultid="12238" heatid="13899" lane="3" entrytime="00:00:35.20" />
                <RESULT eventid="1187" points="271" reactiontime="+110" swimtime="00:00:41.79" resultid="12239" heatid="13946" lane="0" entrytime="00:00:42.50" />
                <RESULT eventid="1256" points="285" reactiontime="+78" swimtime="00:01:19.11" resultid="12240" heatid="13973" lane="3" entrytime="00:01:20.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="252" reactiontime="+82" swimtime="00:01:41.82" resultid="12241" heatid="14002" lane="5" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="217" reactiontime="+86" swimtime="00:03:07.86" resultid="12242" heatid="14041" lane="6" entrytime="00:02:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:28.05" />
                    <SPLIT distance="150" swimtime="00:02:18.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="296" reactiontime="+77" swimtime="00:00:44.21" resultid="12243" heatid="14085" lane="2" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="370" reactiontime="+62" swimtime="00:02:10.11" resultid="12285" heatid="13998" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12301" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="12259" number="2" />
                    <RELAYPOSITION athleteid="12276" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="12264" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="371" reactiontime="+79" swimtime="00:01:58.07" resultid="12286" heatid="14056" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="100" swimtime="00:00:58.74" />
                    <SPLIT distance="150" swimtime="00:01:30.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12301" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="12264" number="2" />
                    <RELAYPOSITION athleteid="12271" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="12276" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="304" reactiontime="+72" swimtime="00:02:37.84" resultid="12287" heatid="13996" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:04.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12305" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="12244" number="2" />
                    <RELAYPOSITION athleteid="12237" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="12230" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="344" reactiontime="+80" swimtime="00:02:17.76" resultid="12288" heatid="14054" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:43.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12305" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="12230" number="2" />
                    <RELAYPOSITION athleteid="12244" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="12237" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="321" reactiontime="+79" swimtime="00:02:03.86" resultid="12281" heatid="13934" lane="1" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                    <SPLIT distance="100" swimtime="00:00:59.46" />
                    <SPLIT distance="150" swimtime="00:01:33.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12276" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="12230" number="2" />
                    <RELAYPOSITION athleteid="12237" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="12264" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="288" reactiontime="+75" swimtime="00:02:21.39" resultid="12282" heatid="14101" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:50.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12301" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="12230" number="2" />
                    <RELAYPOSITION athleteid="12305" number="3" />
                    <RELAYPOSITION athleteid="12264" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="12283" heatid="13934" lane="0" entrytime="00:02:07.11">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12237" number="1" />
                    <RELAYPOSITION athleteid="12259" number="2" />
                    <RELAYPOSITION athleteid="12244" number="3" />
                    <RELAYPOSITION athleteid="12276" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="244" swimtime="00:02:29.42" resultid="12284" heatid="14100" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:01:52.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12237" number="1" />
                    <RELAYPOSITION athleteid="12259" number="2" />
                    <RELAYPOSITION athleteid="12276" number="3" />
                    <RELAYPOSITION athleteid="12244" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WOPRWL" nation="POL" region="LBS" clubid="10831" name="WOPR Województwa Lubuskiego">
          <CONTACT city="Warszawa" email="kifertnat@gmail.com" name="Kifert Natalia" state="LUBUS" street="Lisowskiego 1" zip="65-072" />
          <ATHLETES>
            <ATHLETE birthdate="1975-04-11" firstname="Radomir" gender="M" lastname="Kifert" nation="POL" athleteid="11521">
              <RESULTS>
                <RESULT eventid="1079" points="398" reactiontime="+86" swimtime="00:00:28.41" resultid="11522" heatid="13909" lane="6" entrytime="00:00:31.22" />
                <RESULT eventid="1205" points="399" reactiontime="+77" swimtime="00:00:32.63" resultid="11523" heatid="13957" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1440" points="412" reactiontime="+93" swimtime="00:00:30.14" resultid="11524" heatid="14023" lane="0" entrytime="00:00:32.80" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="11525" heatid="14037" lane="8" entrytime="00:01:12.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-20" firstname="Kalina" gender="F" lastname="Chęcińska" nation="POL" athleteid="11513">
              <RESULTS>
                <RESULT eventid="1062" points="373" reactiontime="+86" swimtime="00:00:32.96" resultid="11514" heatid="13900" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1147" points="256" reactiontime="+99" swimtime="00:12:47.05" resultid="11515" heatid="13936" lane="0" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:14.97" />
                    <SPLIT distance="200" swimtime="00:03:03.39" />
                    <SPLIT distance="250" swimtime="00:03:52.13" />
                    <SPLIT distance="300" swimtime="00:04:41.06" />
                    <SPLIT distance="350" swimtime="00:05:29.73" />
                    <SPLIT distance="400" swimtime="00:06:18.96" />
                    <SPLIT distance="450" swimtime="00:07:07.59" />
                    <SPLIT distance="500" swimtime="00:07:57.25" />
                    <SPLIT distance="550" swimtime="00:08:46.08" />
                    <SPLIT distance="600" swimtime="00:09:35.44" />
                    <SPLIT distance="650" swimtime="00:10:24.38" />
                    <SPLIT distance="700" swimtime="00:11:13.29" />
                    <SPLIT distance="750" swimtime="00:12:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="383" reactiontime="+87" swimtime="00:01:11.70" resultid="11516" heatid="13974" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="268" reactiontime="+95" swimtime="00:00:37.86" resultid="11517" heatid="14016" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1491" points="314" reactiontime="+93" swimtime="00:02:46.19" resultid="11518" heatid="14041" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="242" reactiontime="+91" swimtime="00:01:29.22" resultid="11519" heatid="14064" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="274" reactiontime="+94" swimtime="00:06:06.98" resultid="11520" heatid="14104" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:02:12.94" />
                    <SPLIT distance="200" swimtime="00:03:00.73" />
                    <SPLIT distance="250" swimtime="00:03:48.51" />
                    <SPLIT distance="300" swimtime="00:04:35.84" />
                    <SPLIT distance="350" swimtime="00:05:22.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-25" firstname="Mieszko" gender="M" lastname="Bencych" nation="POL" athleteid="11526">
              <RESULTS>
                <RESULT eventid="1113" points="279" reactiontime="+94" swimtime="00:02:54.29" resultid="11527" heatid="13929" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:10.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="286" reactiontime="+87" swimtime="00:03:12.77" resultid="11528" heatid="13969" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                    <SPLIT distance="150" swimtime="00:02:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="11529" heatid="14010" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="1681" points="370" reactiontime="+85" swimtime="00:00:36.80" resultid="11530" heatid="14094" lane="8" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-20" firstname="Mateusz" gender="M" lastname="Chęciński" nation="POL" athleteid="11534">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1079" points="534" reactiontime="+78" swimtime="00:00:25.77" resultid="11535" heatid="13914" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1205" points="492" swimtime="00:00:30.45" resultid="11536" heatid="13958" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1273" points="518" reactiontime="+90" swimtime="00:00:58.38" resultid="11537" heatid="13987" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="492" reactiontime="+73" swimtime="00:01:05.78" resultid="11538" heatid="14038" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="11539" heatid="14082" lane="2" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-02" firstname="Natalia" gender="F" lastname="Kifert" nation="POL" athleteid="11531">
              <RESULTS>
                <RESULT eventid="1187" points="326" reactiontime="+67" swimtime="00:00:39.30" resultid="11532" heatid="13946" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="11533" heatid="14030" lane="4" entrytime="00:01:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="346" reactiontime="+77" swimtime="00:02:00.76" resultid="11540" heatid="13934" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="100" swimtime="00:00:58.42" />
                    <SPLIT distance="150" swimtime="00:01:32.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11534" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="11513" number="2" />
                    <RELAYPOSITION athleteid="11531" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="11521" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="299" reactiontime="+70" swimtime="00:02:19.70" resultid="11541" heatid="14101" lane="1" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11531" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="11526" number="2" />
                    <RELAYPOSITION athleteid="11513" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="11534" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9728" name="WSB Dąbrowa Górnicza">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="9729">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="9730" heatid="13915" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="9731" heatid="13928" lane="8" entrytime="00:02:45.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="9732" heatid="13957" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="9733" heatid="13967" lane="5" entrytime="00:03:05.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="9734" heatid="14009" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1474" points="272" reactiontime="+73" swimtime="00:01:20.11" resultid="9735" heatid="14035" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="9736" heatid="14080" lane="7" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9354" name="Zawodnicy Niezrzeszeni">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="10762">
              <RESULTS>
                <RESULT eventid="1096" points="200" reactiontime="+91" swimtime="00:03:35.37" resultid="10763" heatid="13919" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="247" swimtime="00:01:42.44" resultid="10764" heatid="14002" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="186" swimtime="00:00:42.76" resultid="10765" heatid="14015" lane="6" entrytime="00:00:44.00" />
                <RESULT eventid="1664" points="245" reactiontime="+92" swimtime="00:00:47.07" resultid="10766" heatid="14085" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-28" firstname="Rafał" gender="M" lastname="Wójcicki" nation="POL" athleteid="9425">
              <RESULTS>
                <RESULT eventid="1205" points="278" reactiontime="+75" swimtime="00:00:36.80" resultid="9426" heatid="13953" lane="2" entrytime="00:00:38.64" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-23" firstname="Marek" gender="M" lastname="Pisulak" nation="POL" athleteid="9934">
              <RESULTS>
                <RESULT eventid="1079" points="101" reactiontime="+106" swimtime="00:00:44.85" resultid="9935" heatid="13905" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="Zieleziński" nation="POL" athleteid="9936">
              <RESULTS>
                <RESULT eventid="1079" points="205" reactiontime="+115" swimtime="00:00:35.42" resultid="9937" heatid="13907" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1205" points="179" reactiontime="+79" swimtime="00:00:42.58" resultid="9939" heatid="13952" lane="6" entrytime="00:00:41.50" />
                <RESULT eventid="1273" points="176" reactiontime="+128" swimtime="00:01:23.61" resultid="9940" heatid="13980" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="142" reactiontime="+85" swimtime="00:01:39.44" resultid="9941" heatid="14032" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="9942" heatid="14046" lane="5" entrytime="00:03:03.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="9943" heatid="14078" lane="6" entrytime="00:03:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-07" firstname="Jerzy" gender="M" lastname="Demetraki-Paleolog" nation="POL" athleteid="9720">
              <RESULTS>
                <RESULT eventid="1113" points="193" reactiontime="+106" swimtime="00:03:17.09" resultid="9721" heatid="13924" lane="5" entrytime="00:03:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="9722" heatid="13965" lane="6" entrytime="00:03:45.10" />
                <RESULT eventid="1341" points="140" reactiontime="+109" swimtime="00:03:34.32" resultid="9723" heatid="13993" lane="3" entrytime="00:03:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                    <SPLIT distance="100" swimtime="00:01:43.71" />
                    <SPLIT distance="150" swimtime="00:02:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="209" reactiontime="+104" swimtime="00:02:51.65" resultid="9724" heatid="14046" lane="4" entrytime="00:03:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="150" swimtime="00:02:09.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="180" reactiontime="+114" swimtime="00:07:11.19" resultid="9725" heatid="14060" lane="7" entrytime="00:07:26.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.37" />
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                    <SPLIT distance="150" swimtime="00:02:43.01" />
                    <SPLIT distance="200" swimtime="00:03:38.41" />
                    <SPLIT distance="250" swimtime="00:04:38.41" />
                    <SPLIT distance="300" swimtime="00:05:39.37" />
                    <SPLIT distance="350" swimtime="00:06:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="164" reactiontime="+107" swimtime="00:01:30.93" resultid="9726" heatid="14068" lane="8" entrytime="00:01:29.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="210" reactiontime="+111" swimtime="00:06:09.96" resultid="9727" heatid="14109" lane="0" entrytime="00:06:17.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:18.52" />
                    <SPLIT distance="200" swimtime="00:03:07.92" />
                    <SPLIT distance="250" swimtime="00:03:54.59" />
                    <SPLIT distance="300" swimtime="00:04:41.94" />
                    <SPLIT distance="350" swimtime="00:05:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-03-29" firstname="Mateusz" gender="M" lastname="Burzawa" nation="POL" athleteid="12463">
              <RESULTS>
                <RESULT eventid="1079" points="500" reactiontime="+73" swimtime="00:00:26.34" resultid="12464" heatid="13914" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1113" points="468" reactiontime="+76" swimtime="00:02:26.79" resultid="12465" heatid="13930" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="442" reactiontime="+76" swimtime="00:00:31.54" resultid="12466" heatid="13956" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1239" points="441" reactiontime="+81" swimtime="00:02:46.84" resultid="12467" heatid="13970" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:02:03.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="457" reactiontime="+77" swimtime="00:01:15.16" resultid="12468" heatid="14012" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="520" reactiontime="+78" swimtime="00:02:06.79" resultid="12469" heatid="14052" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:01.65" />
                    <SPLIT distance="150" swimtime="00:01:34.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-08" firstname="Paweł" gender="M" lastname="Obrzut" nation="POL" athleteid="10759">
              <RESULTS>
                <RESULT eventid="1079" points="252" reactiontime="+77" swimtime="00:00:33.09" resultid="10760" heatid="13908" lane="6" entrytime="00:00:32.17" />
                <RESULT eventid="1273" points="236" reactiontime="+85" swimtime="00:01:15.86" resultid="10761" heatid="13981" lane="1" entrytime="00:01:12.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-02" firstname="Daniel" gender="M" lastname="Osik" nation="POL" athleteid="11081">
              <RESULTS>
                <RESULT eventid="1165" points="382" reactiontime="+90" swimtime="00:19:59.77" resultid="11082" heatid="13943" lane="7" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:46.19" />
                    <SPLIT distance="200" swimtime="00:02:24.40" />
                    <SPLIT distance="250" swimtime="00:03:03.17" />
                    <SPLIT distance="300" swimtime="00:03:42.89" />
                    <SPLIT distance="350" swimtime="00:04:22.67" />
                    <SPLIT distance="400" swimtime="00:05:03.19" />
                    <SPLIT distance="450" swimtime="00:05:43.04" />
                    <SPLIT distance="500" swimtime="00:06:24.34" />
                    <SPLIT distance="550" swimtime="00:11:08.63" />
                    <SPLIT distance="600" swimtime="00:07:45.06" />
                    <SPLIT distance="650" swimtime="00:13:53.66" />
                    <SPLIT distance="700" swimtime="00:09:06.29" />
                    <SPLIT distance="750" swimtime="00:15:15.67" />
                    <SPLIT distance="800" swimtime="00:10:27.86" />
                    <SPLIT distance="900" swimtime="00:11:50.16" />
                    <SPLIT distance="1000" swimtime="00:13:12.38" />
                    <SPLIT distance="1050" swimtime="00:16:39.80" />
                    <SPLIT distance="1100" swimtime="00:14:34.72" />
                    <SPLIT distance="1150" swimtime="00:18:01.87" />
                    <SPLIT distance="1200" swimtime="00:15:58.71" />
                    <SPLIT distance="1300" swimtime="00:17:20.75" />
                    <SPLIT distance="1400" swimtime="00:18:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="400" reactiontime="+75" swimtime="00:02:18.37" resultid="11083" heatid="14052" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="150" swimtime="00:01:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="373" reactiontime="+73" swimtime="00:02:35.46" resultid="11084" heatid="14082" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="417" swimtime="00:04:54.55" resultid="11168" heatid="14106" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="200" swimtime="00:02:25.98" />
                    <SPLIT distance="300" swimtime="00:03:40.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-04-25" firstname="Adriana" gender="F" lastname="Hofman" nation="POL" athleteid="9709">
              <RESULTS>
                <RESULT eventid="1388" points="516" reactiontime="+75" swimtime="00:01:20.21" resultid="9710" heatid="14003" lane="5" entrytime="00:01:30.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="533" reactiontime="+78" swimtime="00:00:36.34" resultid="9711" heatid="14087" lane="7" entrytime="00:00:38.46" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-04-09" firstname="Jerzy" gender="M" lastname="Zaklukiewicz" nation="POL" athleteid="10751">
              <RESULTS>
                <RESULT eventid="1079" points="142" reactiontime="+105" swimtime="00:00:40.03" resultid="10752" heatid="13903" lane="6" />
                <RESULT eventid="1239" points="145" reactiontime="+120" swimtime="00:04:01.49" resultid="10753" heatid="13963" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                    <SPLIT distance="100" swimtime="00:01:53.28" />
                    <SPLIT distance="150" swimtime="00:02:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="78" reactiontime="+106" swimtime="00:01:49.72" resultid="10754" heatid="13977" lane="0" />
                <RESULT eventid="1406" points="152" swimtime="00:01:48.40" resultid="10755" heatid="14005" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="76" reactiontime="+109" swimtime="00:00:52.86" resultid="10756" heatid="14018" lane="5" />
                <RESULT eventid="1681" points="165" reactiontime="+98" swimtime="00:00:48.11" resultid="10757" heatid="14088" lane="5" />
                <RESULT eventid="1744" points="52" reactiontime="+112" swimtime="00:09:46.42" resultid="10758" heatid="14106" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.59" />
                    <SPLIT distance="100" swimtime="00:02:11.62" />
                    <SPLIT distance="150" swimtime="00:03:25.57" />
                    <SPLIT distance="200" swimtime="00:04:44.90" />
                    <SPLIT distance="250" swimtime="00:06:02.67" />
                    <SPLIT distance="300" swimtime="00:07:22.21" />
                    <SPLIT distance="350" swimtime="00:08:37.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="12455">
              <RESULTS>
                <RESULT eventid="1079" points="252" swimtime="00:00:33.07" resultid="12456" heatid="13909" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1165" points="179" reactiontime="+114" swimtime="00:25:43.47" resultid="12457" heatid="13941" lane="0" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:31.08" />
                    <SPLIT distance="150" swimtime="00:05:51.81" />
                    <SPLIT distance="200" swimtime="00:03:14.55" />
                    <SPLIT distance="250" swimtime="00:09:20.25" />
                    <SPLIT distance="300" swimtime="00:04:58.96" />
                    <SPLIT distance="350" swimtime="00:11:05.58" />
                    <SPLIT distance="400" swimtime="00:08:28.35" />
                    <SPLIT distance="450" swimtime="00:12:52.01" />
                    <SPLIT distance="500" swimtime="00:11:57.62" />
                    <SPLIT distance="550" swimtime="00:14:35.80" />
                    <SPLIT distance="600" swimtime="00:13:43.25" />
                    <SPLIT distance="650" swimtime="00:16:23.46" />
                    <SPLIT distance="700" swimtime="00:15:30.12" />
                    <SPLIT distance="750" swimtime="00:18:09.11" />
                    <SPLIT distance="800" swimtime="00:17:16.86" />
                    <SPLIT distance="850" swimtime="00:19:54.63" />
                    <SPLIT distance="900" swimtime="00:19:02.42" />
                    <SPLIT distance="950" swimtime="00:21:37.01" />
                    <SPLIT distance="1000" swimtime="00:20:46.07" />
                    <SPLIT distance="1050" swimtime="00:23:19.63" />
                    <SPLIT distance="1100" swimtime="00:22:28.77" />
                    <SPLIT distance="1200" swimtime="00:24:10.85" />
                    <SPLIT distance="1450" swimtime="00:25:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="267" reactiontime="+96" swimtime="00:01:12.84" resultid="12458" heatid="13981" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="204" reactiontime="+102" swimtime="00:02:53.02" resultid="12459" heatid="14048" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:10.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="205" swimtime="00:06:12.63" resultid="12460" heatid="14109" lane="6" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:14.32" />
                    <SPLIT distance="200" swimtime="00:03:03.08" />
                    <SPLIT distance="250" swimtime="00:03:50.95" />
                    <SPLIT distance="300" swimtime="00:04:39.35" />
                    <SPLIT distance="350" swimtime="00:05:28.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" athleteid="10873">
              <RESULTS>
                <RESULT eventid="1079" points="471" reactiontime="+76" swimtime="00:00:26.87" resultid="10874" heatid="13916" lane="4" entrytime="00:00:25.80" entrycourse="LCM" />
                <RESULT eventid="1273" points="525" reactiontime="+87" swimtime="00:00:58.13" resultid="10875" heatid="13989" lane="1" entrytime="00:00:56.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="440" reactiontime="+76" swimtime="00:02:14.05" resultid="10876" heatid="14053" lane="7" entrytime="00:02:08.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.83" />
                    <SPLIT distance="150" swimtime="00:01:38.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-19" firstname="Marcin" gender="M" lastname="Patyk" nation="POL" athleteid="9857">
              <RESULTS>
                <RESULT eventid="1079" points="328" reactiontime="+92" swimtime="00:00:30.29" resultid="9858" heatid="13910" lane="5" entrytime="00:00:30.50" entrycourse="SCM" />
                <RESULT eventid="1273" points="273" reactiontime="+94" swimtime="00:01:12.30" resultid="9859" heatid="13980" lane="4" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="338" reactiontime="+97" swimtime="00:00:32.18" resultid="9860" heatid="14023" lane="7" entrytime="00:00:32.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-03" firstname="Patryk" gender="M" lastname="Dzwonek" nation="POL" athleteid="12754">
              <RESULTS>
                <RESULT eventid="1079" points="464" reactiontime="+105" swimtime="00:00:27.00" resultid="12755" heatid="13903" lane="7" />
                <RESULT eventid="1273" points="439" swimtime="00:01:01.72" resultid="12756" heatid="13977" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="12757" heatid="14032" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="9355">
              <RESULTS>
                <RESULT eventid="1165" points="112" reactiontime="+107" swimtime="00:30:04.90" resultid="9356" heatid="13939" lane="7" entrytime="00:33:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                    <SPLIT distance="100" swimtime="00:01:48.32" />
                    <SPLIT distance="150" swimtime="00:02:46.44" />
                    <SPLIT distance="200" swimtime="00:03:45.88" />
                    <SPLIT distance="250" swimtime="00:04:45.81" />
                    <SPLIT distance="300" swimtime="00:05:46.36" />
                    <SPLIT distance="350" swimtime="00:06:46.54" />
                    <SPLIT distance="400" swimtime="00:07:46.77" />
                    <SPLIT distance="450" swimtime="00:08:46.58" />
                    <SPLIT distance="500" swimtime="00:09:46.11" />
                    <SPLIT distance="550" swimtime="00:10:46.39" />
                    <SPLIT distance="600" swimtime="00:11:47.40" />
                    <SPLIT distance="650" swimtime="00:12:47.72" />
                    <SPLIT distance="700" swimtime="00:13:48.14" />
                    <SPLIT distance="750" swimtime="00:14:49.12" />
                    <SPLIT distance="800" swimtime="00:15:49.75" />
                    <SPLIT distance="850" swimtime="00:16:50.55" />
                    <SPLIT distance="900" swimtime="00:17:51.30" />
                    <SPLIT distance="950" swimtime="00:18:51.76" />
                    <SPLIT distance="1000" swimtime="00:19:53.28" />
                    <SPLIT distance="1050" swimtime="00:20:53.83" />
                    <SPLIT distance="1100" swimtime="00:21:55.78" />
                    <SPLIT distance="1150" swimtime="00:22:57.02" />
                    <SPLIT distance="1200" swimtime="00:24:00.18" />
                    <SPLIT distance="1250" swimtime="00:25:02.32" />
                    <SPLIT distance="1300" swimtime="00:26:05.74" />
                    <SPLIT distance="1350" swimtime="00:27:06.98" />
                    <SPLIT distance="1400" swimtime="00:28:09.70" />
                    <SPLIT distance="1450" swimtime="00:29:09.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="115" reactiontime="+104" swimtime="00:01:36.20" resultid="9357" heatid="13978" lane="4" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="106" reactiontime="+103" swimtime="00:03:35.48" resultid="9358" heatid="14046" lane="9" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:45.42" />
                    <SPLIT distance="150" swimtime="00:02:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="111" reactiontime="+126" swimtime="00:07:37.70" resultid="9359" heatid="14107" lane="2" entrytime="00:07:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                    <SPLIT distance="100" swimtime="00:01:48.38" />
                    <SPLIT distance="150" swimtime="00:02:47.04" />
                    <SPLIT distance="200" swimtime="00:03:46.12" />
                    <SPLIT distance="250" swimtime="00:04:44.92" />
                    <SPLIT distance="300" swimtime="00:05:43.55" />
                    <SPLIT distance="350" swimtime="00:06:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kaziemierz" gender="M" lastname="Sinicki" nation="POL" athleteid="9600">
              <RESULTS>
                <RESULT eventid="1079" points="326" reactiontime="+85" swimtime="00:00:30.37" resultid="9601" heatid="13910" lane="1" entrytime="00:00:30.65" />
                <RESULT eventid="1273" points="311" reactiontime="+89" swimtime="00:01:09.23" resultid="9602" heatid="13982" lane="2" entrytime="00:01:09.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="249" reactiontime="+85" swimtime="00:00:35.63" resultid="9603" heatid="14020" lane="1" entrytime="00:00:37.65" />
                <RESULT eventid="1508" points="260" reactiontime="+88" swimtime="00:02:39.72" resultid="9604" heatid="14049" lane="0" entrytime="00:02:39.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Aleksandra" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="11800">
              <RESULTS>
                <RESULT eventid="1187" points="553" reactiontime="+65" swimtime="00:00:32.96" resultid="11801" heatid="13948" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="1256" points="507" reactiontime="+69" swimtime="00:01:05.26" resultid="11802" heatid="13975" lane="4" entrytime="00:01:08.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="11803" heatid="14003" lane="9" entrytime="00:01:35.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="11804" heatid="14031" lane="7" entrytime="00:01:15.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-30" firstname="Patryk" gender="M" lastname="Suchodolski" nation="POL" athleteid="11636">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="11637" heatid="13928" lane="9" entrytime="00:02:45.00" />
                <RESULT eventid="1205" points="478" reactiontime="+64" swimtime="00:00:30.73" resultid="11638" heatid="13957" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1239" points="439" reactiontime="+75" swimtime="00:02:47.07" resultid="11639" heatid="13970" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:02:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="11640" heatid="14013" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="11641" heatid="14026" lane="5" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-02" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="10739">
              <RESULTS>
                <RESULT eventid="1113" points="229" reactiontime="+90" swimtime="00:03:06.09" resultid="10740" heatid="13925" lane="4" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:21.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="185" reactiontime="+102" swimtime="00:03:15.65" resultid="10741" heatid="13994" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:28.39" />
                    <SPLIT distance="150" swimtime="00:02:22.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="277" reactiontime="+89" swimtime="00:00:34.39" resultid="10742" heatid="14021" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1613" points="214" swimtime="00:01:23.21" resultid="10743" heatid="14069" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-21" firstname="Robert" gender="M" lastname="Maciejewski" nation="POL" athleteid="10744">
              <RESULTS>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="10745" heatid="14076" lane="5" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="10746" heatid="14088" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-09-10" firstname="Agnieszka" gender="F" lastname="Podstawska" nation="POL" athleteid="9983">
              <RESULTS>
                <RESULT eventid="1062" points="217" reactiontime="+96" swimtime="00:00:39.43" resultid="9984" heatid="13898" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1187" points="151" reactiontime="+80" swimtime="00:00:50.75" resultid="9985" heatid="13945" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="1256" points="198" reactiontime="+91" swimtime="00:01:29.22" resultid="9986" heatid="13972" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="185" reactiontime="+93" swimtime="00:03:17.97" resultid="9987" heatid="14040" lane="7" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="100" swimtime="00:01:34.52" />
                    <SPLIT distance="150" swimtime="00:02:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="135" reactiontime="+101" swimtime="00:00:57.36" resultid="9988" heatid="14083" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1721" points="174" swimtime="00:07:06.30" resultid="9989" heatid="14103" lane="0" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:37.03" />
                    <SPLIT distance="200" swimtime="00:03:25.64" />
                    <SPLIT distance="250" swimtime="00:04:22.02" />
                    <SPLIT distance="300" swimtime="00:05:18.12" />
                    <SPLIT distance="350" swimtime="00:06:14.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-02" firstname="Janusz" gender="M" lastname="Konstanty" nation="POL" athleteid="9769">
              <RESULTS>
                <RESULT eventid="1113" points="212" reactiontime="+104" swimtime="00:03:10.98" resultid="9770" heatid="13924" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="254" reactiontime="+83" swimtime="00:00:37.93" resultid="9771" heatid="13953" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1474" points="232" reactiontime="+80" swimtime="00:01:24.41" resultid="9772" heatid="14034" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="9773" heatid="14059" lane="4" entrytime="00:07:45.00" />
                <RESULT eventid="1647" points="217" reactiontime="+57" swimtime="00:03:06.02" resultid="9774" heatid="14079" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="150" swimtime="00:02:19.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-03-06" firstname="Andrzej" gender="M" lastname="Pawlak" nation="POL" athleteid="9647">
              <RESULTS>
                <RESULT eventid="1079" points="246" reactiontime="+113" swimtime="00:00:33.36" resultid="9648" heatid="13907" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1113" points="163" reactiontime="+110" swimtime="00:03:28.63" resultid="9649" heatid="13924" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:41.30" />
                    <SPLIT distance="150" swimtime="00:02:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="209" reactiontime="+74" swimtime="00:00:40.50" resultid="9650" heatid="13952" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="9651" heatid="14078" lane="3" entrytime="00:03:30.00" />
                <RESULT eventid="1744" points="130" reactiontime="+112" swimtime="00:07:13.69" resultid="9652" heatid="14108" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="150" swimtime="00:02:34.41" />
                    <SPLIT distance="200" swimtime="00:03:30.43" />
                    <SPLIT distance="250" swimtime="00:04:26.74" />
                    <SPLIT distance="300" swimtime="00:05:23.71" />
                    <SPLIT distance="350" swimtime="00:06:20.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" athleteid="9427">
              <RESULTS>
                <RESULT eventid="1165" points="448" reactiontime="+90" swimtime="00:18:58.15" resultid="9428" heatid="13943" lane="1" entrytime="00:19:28.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:45.92" />
                    <SPLIT distance="200" swimtime="00:02:23.44" />
                    <SPLIT distance="250" swimtime="00:03:00.60" />
                    <SPLIT distance="300" swimtime="00:04:54.08" />
                    <SPLIT distance="350" swimtime="00:04:16.13" />
                    <SPLIT distance="400" swimtime="00:06:10.43" />
                    <SPLIT distance="450" swimtime="00:05:32.14" />
                    <SPLIT distance="550" swimtime="00:06:48.47" />
                    <SPLIT distance="600" swimtime="00:07:26.96" />
                    <SPLIT distance="650" swimtime="00:08:05.26" />
                    <SPLIT distance="700" swimtime="00:08:43.54" />
                    <SPLIT distance="750" swimtime="00:09:21.74" />
                    <SPLIT distance="800" swimtime="00:10:00.57" />
                    <SPLIT distance="850" swimtime="00:10:38.79" />
                    <SPLIT distance="900" swimtime="00:11:17.33" />
                    <SPLIT distance="950" swimtime="00:11:55.97" />
                    <SPLIT distance="1000" swimtime="00:12:34.35" />
                    <SPLIT distance="1050" swimtime="00:13:12.79" />
                    <SPLIT distance="1100" swimtime="00:13:51.01" />
                    <SPLIT distance="1150" swimtime="00:14:29.48" />
                    <SPLIT distance="1200" swimtime="00:15:08.21" />
                    <SPLIT distance="1250" swimtime="00:15:46.54" />
                    <SPLIT distance="1300" swimtime="00:16:25.12" />
                    <SPLIT distance="1350" swimtime="00:17:03.73" />
                    <SPLIT distance="1400" swimtime="00:17:42.20" />
                    <SPLIT distance="1450" swimtime="00:18:20.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="361" reactiontime="+60" swimtime="00:01:12.93" resultid="9429" heatid="14036" lane="4" entrytime="00:01:14.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="438" reactiontime="+91" swimtime="00:02:14.25" resultid="9430" heatid="14052" lane="8" entrytime="00:02:14.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="405" reactiontime="+67" swimtime="00:02:31.23" resultid="9431" heatid="14081" lane="4" entrytime="00:02:34.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="464" reactiontime="+92" swimtime="00:04:44.06" resultid="9432" heatid="14113" lane="7" entrytime="00:04:54.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:41.29" />
                    <SPLIT distance="200" swimtime="00:02:17.80" />
                    <SPLIT distance="250" swimtime="00:02:54.15" />
                    <SPLIT distance="300" swimtime="00:03:31.37" />
                    <SPLIT distance="350" swimtime="00:04:07.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="9397">
              <RESULTS>
                <RESULT eventid="1079" points="132" reactiontime="+108" swimtime="00:00:41.01" resultid="9398" heatid="13906" lane="0" entrytime="00:00:39.50" />
                <RESULT eventid="1165" points="112" reactiontime="+129" swimtime="00:30:03.76" resultid="9399" heatid="13939" lane="3" entrytime="00:29:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                    <SPLIT distance="100" swimtime="00:01:50.38" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                    <SPLIT distance="200" swimtime="00:03:48.89" />
                    <SPLIT distance="250" swimtime="00:04:48.30" />
                    <SPLIT distance="300" swimtime="00:05:48.22" />
                    <SPLIT distance="350" swimtime="00:06:48.70" />
                    <SPLIT distance="400" swimtime="00:07:49.75" />
                    <SPLIT distance="450" swimtime="00:08:49.58" />
                    <SPLIT distance="500" swimtime="00:09:50.99" />
                    <SPLIT distance="550" swimtime="00:10:51.20" />
                    <SPLIT distance="600" swimtime="00:11:52.48" />
                    <SPLIT distance="650" swimtime="00:12:54.41" />
                    <SPLIT distance="700" swimtime="00:13:55.36" />
                    <SPLIT distance="750" swimtime="00:14:56.89" />
                    <SPLIT distance="800" swimtime="00:15:56.72" />
                    <SPLIT distance="850" swimtime="00:16:57.29" />
                    <SPLIT distance="900" swimtime="00:17:59.32" />
                    <SPLIT distance="950" swimtime="00:19:01.59" />
                    <SPLIT distance="1000" swimtime="00:20:02.36" />
                    <SPLIT distance="1050" swimtime="00:21:04.24" />
                    <SPLIT distance="1100" swimtime="00:22:05.15" />
                    <SPLIT distance="1150" swimtime="00:23:06.40" />
                    <SPLIT distance="1200" swimtime="00:24:05.51" />
                    <SPLIT distance="1250" swimtime="00:25:07.31" />
                    <SPLIT distance="1300" swimtime="00:26:08.03" />
                    <SPLIT distance="1350" swimtime="00:27:09.99" />
                    <SPLIT distance="1400" swimtime="00:28:10.75" />
                    <SPLIT distance="1450" swimtime="00:29:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="102" reactiontime="+116" swimtime="00:00:51.43" resultid="9400" heatid="13951" lane="3" entrytime="00:00:49.50" />
                <RESULT eventid="1273" points="116" reactiontime="+112" swimtime="00:01:35.93" resultid="9401" heatid="13979" lane="7" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="122" reactiontime="+119" swimtime="00:00:45.17" resultid="9402" heatid="14019" lane="2" entrytime="00:00:43.50" />
                <RESULT eventid="1474" points="80" reactiontime="+100" swimtime="00:02:00.17" resultid="9403" heatid="14033" lane="5" entrytime="00:01:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="78" reactiontime="+100" swimtime="00:04:21.62" resultid="9404" heatid="14077" lane="4" entrytime="00:04:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.08" />
                    <SPLIT distance="100" swimtime="00:02:10.80" />
                    <SPLIT distance="150" swimtime="00:03:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="117" reactiontime="+112" swimtime="00:07:29.14" resultid="9405" heatid="14107" lane="3" entrytime="00:07:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                    <SPLIT distance="100" swimtime="00:01:46.46" />
                    <SPLIT distance="150" swimtime="00:02:45.45" />
                    <SPLIT distance="200" swimtime="00:03:43.21" />
                    <SPLIT distance="250" swimtime="00:04:42.85" />
                    <SPLIT distance="300" swimtime="00:05:39.39" />
                    <SPLIT distance="350" swimtime="00:06:37.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="9712">
              <RESULTS>
                <RESULT eventid="1079" points="386" reactiontime="+78" swimtime="00:00:28.70" resultid="9713" heatid="13912" lane="7" entrytime="00:00:28.75" />
                <RESULT eventid="1113" points="338" reactiontime="+82" swimtime="00:02:43.56" resultid="9714" heatid="13928" lane="3" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:02:04.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="388" reactiontime="+83" swimtime="00:01:04.30" resultid="9715" heatid="13985" lane="2" entrytime="00:01:02.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="387" reactiontime="+84" swimtime="00:00:30.76" resultid="9716" heatid="14025" lane="0" entrytime="00:00:30.75" />
                <RESULT eventid="1508" points="322" reactiontime="+88" swimtime="00:02:28.79" resultid="9717" heatid="14050" lane="2" entrytime="00:02:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="328" reactiontime="+82" swimtime="00:01:12.23" resultid="9718" heatid="14070" lane="7" entrytime="00:01:10.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="334" swimtime="00:00:38.05" resultid="9719" heatid="14093" lane="6" entrytime="00:00:38.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Weronika" gender="F" lastname="Kabut" nation="POL" athleteid="11085">
              <RESULTS>
                <RESULT eventid="1062" points="485" reactiontime="+74" swimtime="00:00:30.19" resultid="11086" heatid="13901" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1096" points="388" reactiontime="+71" swimtime="00:02:52.79" resultid="11087" heatid="13920" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="336" reactiontime="+79" swimtime="00:00:38.91" resultid="11088" heatid="13947" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1256" points="470" reactiontime="+75" swimtime="00:01:06.93" resultid="11089" heatid="13975" lane="3" entrytime="00:01:09.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="358" reactiontime="+78" swimtime="00:00:34.39" resultid="11090" heatid="14016" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1491" points="411" reactiontime="+78" swimtime="00:02:31.90" resultid="11091" heatid="14042" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="300" reactiontime="+81" swimtime="00:01:23.10" resultid="11092" heatid="14065" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="354" reactiontime="+81" swimtime="00:05:36.93" resultid="11093" heatid="14104" lane="2" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="150" swimtime="00:02:00.50" />
                    <SPLIT distance="200" swimtime="00:02:44.35" />
                    <SPLIT distance="250" swimtime="00:03:28.26" />
                    <SPLIT distance="300" swimtime="00:04:12.81" />
                    <SPLIT distance="350" swimtime="00:04:56.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="11542">
              <RESULTS>
                <RESULT eventid="1079" points="156" reactiontime="+130" swimtime="00:00:38.82" resultid="11543" heatid="13906" lane="1" entrytime="00:00:38.22" />
                <RESULT eventid="1681" points="144" swimtime="00:00:50.38" resultid="11544" heatid="14090" lane="6" entrytime="00:00:49.76" />
                <RESULT eventid="1744" points="122" reactiontime="+113" swimtime="00:07:22.52" resultid="11545" heatid="14108" lane="7" entrytime="00:06:43.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                    <SPLIT distance="100" swimtime="00:01:41.30" />
                    <SPLIT distance="150" swimtime="00:02:38.41" />
                    <SPLIT distance="200" swimtime="00:03:36.03" />
                    <SPLIT distance="250" swimtime="00:04:32.73" />
                    <SPLIT distance="300" swimtime="00:05:31.12" />
                    <SPLIT distance="350" swimtime="00:06:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-24" firstname="Igor" gender="M" lastname="Okarmus" nation="POL" athleteid="9645">
              <RESULTS>
                <RESULT eventid="1744" points="303" reactiontime="+97" swimtime="00:05:27.35" resultid="9646" heatid="14113" lane="0" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:33.99" />
                    <SPLIT distance="250" swimtime="00:03:17.02" />
                    <SPLIT distance="300" swimtime="00:04:01.30" />
                    <SPLIT distance="350" swimtime="00:04:44.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="9421">
              <RESULTS>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="9423" heatid="14045" lane="8" />
                <RESULT eventid="1744" points="138" reactiontime="+110" swimtime="00:07:05.80" resultid="9424" heatid="14106" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:33.20" />
                    <SPLIT distance="150" swimtime="00:02:29.42" />
                    <SPLIT distance="200" swimtime="00:03:25.08" />
                    <SPLIT distance="250" swimtime="00:04:22.12" />
                    <SPLIT distance="300" swimtime="00:05:18.81" />
                    <SPLIT distance="350" swimtime="00:06:14.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZKS DRZONK" nation="POL" region="LBS" clubid="9738" name="ZKS Drzonków">
          <CONTACT city="łężyca/Zielona Góra" email="llfpiotr@gmail.com" name="Barta" phone="602347348" state="LUBUS" street="Odrzańska" zip="66-016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="Piotr" gender="M" lastname="Barta" nameprefix="Mr." nation="POL" athleteid="9739">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1239" points="509" reactiontime="+82" swimtime="00:02:38.99" resultid="9740" heatid="13970" lane="2" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="494" reactiontime="+77" swimtime="00:01:13.26" resultid="9741" heatid="14013" lane="1" entrytime="00:01:13.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="1578" points="411" reactiontime="+82" swimtime="00:05:27.77" resultid="9742" heatid="14062" lane="7" entrytime="00:05:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                    <SPLIT distance="200" swimtime="00:02:43.26" />
                    <SPLIT distance="250" swimtime="00:03:27.28" />
                    <SPLIT distance="300" swimtime="00:04:12.32" />
                    <SPLIT distance="350" swimtime="00:04:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="9743" heatid="14097" lane="5" entrytime="00:00:33.13" entrycourse="LCM" />
                <RESULT eventid="1744" points="450" reactiontime="+80" swimtime="00:04:47.07" resultid="9744" heatid="14113" lane="4" entrytime="00:04:44.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:47.09" />
                    <SPLIT distance="200" swimtime="00:02:23.57" />
                    <SPLIT distance="250" swimtime="00:02:59.31" />
                    <SPLIT distance="300" swimtime="00:03:35.26" />
                    <SPLIT distance="350" swimtime="00:04:11.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

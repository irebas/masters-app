<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KS Warszawianka" version="11.71436">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Warszawa" name="XXVI WARSAW OPEN MISTRZOSTWA WARSZAWY MASTERS W PŁYWANIU" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-12-04" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Warszawa" nation="POL" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <QUALIFY from="2020-01-01" until="2021-12-03" />
      <SESSIONS>
        <SESSION date="2021-12-04" daytime="16:30" endtime="19:13" name="I BLOK" number="1" warmupfrom="15:30" warmupuntil="16:15">
          <EVENTS>
            <EVENT eventid="1058" daytime="16:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1102" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3361" />
                    <RANKING order="2" place="2" resultid="3735" />
                    <RANKING order="3" place="3" resultid="3505" />
                    <RANKING order="4" place="4" resultid="3256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3763" />
                    <RANKING order="2" place="2" resultid="3275" />
                    <RANKING order="3" place="3" resultid="3502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3388" />
                    <RANKING order="2" place="2" resultid="3598" />
                    <RANKING order="3" place="3" resultid="3493" />
                    <RANKING order="4" place="4" resultid="3771" />
                    <RANKING order="5" place="5" resultid="3792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3695" />
                    <RANKING order="2" place="2" resultid="3290" />
                    <RANKING order="3" place="3" resultid="3343" />
                    <RANKING order="4" place="4" resultid="3465" />
                    <RANKING order="5" place="5" resultid="3341" />
                    <RANKING order="6" place="-1" resultid="3363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3583" />
                    <RANKING order="2" place="2" resultid="3412" />
                    <RANKING order="3" place="3" resultid="3808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3441" />
                    <RANKING order="2" place="2" resultid="3810" />
                    <RANKING order="3" place="3" resultid="3628" />
                    <RANKING order="4" place="4" resultid="3569" />
                    <RANKING order="5" place="5" resultid="3744" />
                    <RANKING order="6" place="6" resultid="3270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1095" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1096" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1097" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1099" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1100" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1101" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3932" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3933" daytime="16:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3934" daytime="16:33" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="16:35" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3741" />
                    <RANKING order="2" place="2" resultid="3604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3224" />
                    <RANKING order="2" place="2" resultid="3618" />
                    <RANKING order="3" place="3" resultid="3400" />
                    <RANKING order="4" place="4" resultid="3680" />
                    <RANKING order="5" place="5" resultid="3683" />
                    <RANKING order="6" place="6" resultid="3373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                    <RANKING order="2" place="2" resultid="3471" />
                    <RANKING order="3" place="3" resultid="3444" />
                    <RANKING order="4" place="-1" resultid="3349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3586" />
                    <RANKING order="2" place="2" resultid="3300" />
                    <RANKING order="3" place="3" resultid="3382" />
                    <RANKING order="4" place="4" resultid="3576" />
                    <RANKING order="5" place="5" resultid="3760" />
                    <RANKING order="6" place="6" resultid="3287" />
                    <RANKING order="7" place="7" resultid="3533" />
                    <RANKING order="8" place="8" resultid="3520" />
                    <RANKING order="9" place="9" resultid="3247" />
                    <RANKING order="10" place="10" resultid="3798" />
                    <RANKING order="11" place="11" resultid="3755" />
                    <RANKING order="12" place="-1" resultid="3786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3571" />
                    <RANKING order="2" place="2" resultid="3462" />
                    <RANKING order="3" place="3" resultid="3397" />
                    <RANKING order="4" place="4" resultid="3558" />
                    <RANKING order="5" place="5" resultid="3718" />
                    <RANKING order="6" place="6" resultid="3631" />
                    <RANKING order="7" place="7" resultid="3804" />
                    <RANKING order="8" place="8" resultid="3647" />
                    <RANKING order="9" place="9" resultid="3447" />
                    <RANKING order="10" place="10" resultid="3459" />
                    <RANKING order="11" place="11" resultid="3738" />
                    <RANKING order="12" place="12" resultid="3496" />
                    <RANKING order="13" place="13" resultid="3757" />
                    <RANKING order="14" place="14" resultid="3439" />
                    <RANKING order="15" place="15" resultid="3357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3601" />
                    <RANKING order="2" place="2" resultid="3221" />
                    <RANKING order="3" place="3" resultid="3483" />
                    <RANKING order="4" place="4" resultid="3726" />
                    <RANKING order="5" place="5" resultid="3214" />
                    <RANKING order="6" place="6" resultid="3335" />
                    <RANKING order="7" place="-1" resultid="3701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3514" />
                    <RANKING order="2" place="2" resultid="3250" />
                    <RANKING order="3" place="3" resultid="3231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3766" />
                    <RANKING order="2" place="2" resultid="3774" />
                    <RANKING order="3" place="3" resultid="3474" />
                    <RANKING order="4" place="4" resultid="3235" />
                    <RANKING order="5" place="5" resultid="3297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3477" />
                    <RANKING order="2" place="2" resultid="3715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3330" />
                    <RANKING order="2" place="2" resultid="3421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1116" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1117" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1118" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3935" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3936" daytime="16:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3937" daytime="16:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3938" daytime="16:39" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3939" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3940" daytime="16:42" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="16:44" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1120" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1121" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3732" />
                    <RANKING order="2" place="2" resultid="3309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1124" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3584" />
                    <RANKING order="2" place="2" resultid="3698" />
                    <RANKING order="3" place="3" resultid="3809" />
                    <RANKING order="4" place="4" resultid="3753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3811" />
                    <RANKING order="2" place="2" resultid="3427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1128" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1129" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1130" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1131" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1132" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1133" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1134" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3941" daytime="16:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="16:45" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1136" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3225" />
                    <RANKING order="2" place="2" resultid="3621" />
                    <RANKING order="3" place="3" resultid="3777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1140" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3281" />
                    <RANKING order="2" place="2" resultid="3460" />
                    <RANKING order="3" place="3" resultid="3634" />
                    <RANKING order="4" place="-1" resultid="3278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3594" />
                    <RANKING order="2" place="2" resultid="3272" />
                    <RANKING order="3" place="-1" resultid="3541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3538" />
                    <RANKING order="2" place="2" resultid="3515" />
                    <RANKING order="3" place="3" resultid="3232" />
                    <RANKING order="4" place="4" resultid="3267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3650" />
                    <RANKING order="2" place="2" resultid="3298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3724" />
                    <RANKING order="2" place="2" resultid="3712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1148" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1149" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1150" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3942" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3943" daytime="16:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3944" daytime="16:49" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="16:51" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3506" />
                    <RANKING order="2" place="2" resultid="3736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3764" />
                    <RANKING order="2" place="2" resultid="3550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3437" />
                    <RANKING order="2" place="2" resultid="3703" />
                    <RANKING order="3" place="3" resultid="3772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3344" />
                    <RANKING order="2" place="2" resultid="3931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                    <RANKING order="2" place="2" resultid="3508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1160" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1161" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1162" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1163" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1164" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1165" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1166" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3945" daytime="16:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3946" daytime="16:53" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="16:55" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1168" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1169" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3306" />
                    <RANKING order="2" place="2" resultid="3684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3761" />
                    <RANKING order="2" place="-1" resultid="3787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3653" />
                    <RANKING order="2" place="2" resultid="3463" />
                    <RANKING order="3" place="3" resultid="3317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1174" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3370" />
                    <RANKING order="2" place="2" resultid="3561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1180" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1181" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1182" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3947" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3948" daytime="16:57" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="16:59" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1185" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3733" />
                    <RANKING order="2" place="2" resultid="3310" />
                    <RANKING order="3" place="3" resultid="3276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3456" />
                    <RANKING order="2" place="2" resultid="3291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1189" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1190" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1193" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1194" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1195" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1196" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1197" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1198" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3949" daytime="16:59" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="17:01" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3619" />
                    <RANKING order="2" place="2" resultid="3401" />
                    <RANKING order="3" place="3" resultid="3929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3780" />
                    <RANKING order="2" place="2" resultid="3391" />
                    <RANKING order="3" place="-1" resultid="3624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3359" />
                    <RANKING order="2" place="2" resultid="3430" />
                    <RANKING order="3" place="3" resultid="3729" />
                    <RANKING order="4" place="4" resultid="3383" />
                    <RANKING order="5" place="5" resultid="3577" />
                    <RANKING order="6" place="6" resultid="3521" />
                    <RANKING order="7" place="7" resultid="3801" />
                    <RANKING order="8" place="8" resultid="3241" />
                    <RANKING order="9" place="9" resultid="3346" />
                    <RANKING order="10" place="-1" resultid="3799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3654" />
                    <RANKING order="2" place="2" resultid="3398" />
                    <RANKING order="3" place="3" resultid="3632" />
                    <RANKING order="4" place="4" resultid="3805" />
                    <RANKING order="5" place="5" resultid="3573" />
                    <RANKING order="6" place="-1" resultid="3480" />
                    <RANKING order="7" place="-1" resultid="3279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3727" />
                    <RANKING order="2" place="2" resultid="3273" />
                    <RANKING order="3" place="-1" resultid="3336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3579" />
                    <RANKING order="2" place="2" resultid="3637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3544" />
                    <RANKING order="2" place="2" resultid="3475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1210" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1212" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1213" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1214" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3950" daytime="17:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3951" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3952" daytime="17:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3953" daytime="17:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1215" daytime="17:08" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1216" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1217" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1219" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1220" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3565" />
                    <RANKING order="2" place="2" resultid="3413" />
                    <RANKING order="3" place="3" resultid="3263" />
                    <RANKING order="4" place="4" resultid="3323" />
                    <RANKING order="5" place="-1" resultid="3403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3207" />
                    <RANKING order="2" place="2" resultid="3320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1224" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1226" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1227" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1228" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1229" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1230" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3954" daytime="17:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1231" daytime="17:13" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1232" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1236" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3203" />
                    <RANKING order="2" place="2" resultid="3662" />
                    <RANKING order="3" place="3" resultid="3739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3394" />
                    <RANKING order="2" place="2" resultid="3659" />
                    <RANKING order="3" place="3" resultid="3614" />
                    <RANKING order="4" place="4" resultid="3326" />
                    <RANKING order="5" place="5" resultid="3376" />
                    <RANKING order="6" place="6" resultid="3217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1243" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1244" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1245" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1246" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3955" daytime="17:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3956" daytime="17:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1247" daytime="17:24" gender="F" number="11" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3145" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3146" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3201" />
                    <RANKING order="2" place="2" resultid="3747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3147" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3677" />
                    <RANKING order="2" place="-1" resultid="3793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3148" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3466" />
                    <RANKING order="2" place="2" resultid="3259" />
                    <RANKING order="3" place="-1" resultid="3364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3149" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="3150" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3629" />
                    <RANKING order="2" place="2" resultid="3415" />
                    <RANKING order="3" place="3" resultid="3745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3151" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3152" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3153" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="3154" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="3155" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3156" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3157" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3158" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3159" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3957" daytime="17:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3958" daytime="17:27" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1295" daytime="17:29" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1296" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1297" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3681" />
                    <RANKING order="2" place="2" resultid="3750" />
                    <RANKING order="3" place="3" resultid="3930" />
                    <RANKING order="4" place="4" resultid="3374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3783" />
                    <RANKING order="2" place="2" resultid="3304" />
                    <RANKING order="3" place="3" resultid="3472" />
                    <RANKING order="4" place="4" resultid="3445" />
                    <RANKING order="5" place="5" resultid="3517" />
                    <RANKING order="6" place="6" resultid="3284" />
                    <RANKING order="7" place="-1" resultid="3625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3587" />
                    <RANKING order="2" place="2" resultid="3730" />
                    <RANKING order="3" place="3" resultid="3301" />
                    <RANKING order="4" place="4" resultid="3288" />
                    <RANKING order="5" place="5" resultid="3802" />
                    <RANKING order="6" place="6" resultid="3248" />
                    <RANKING order="7" place="7" resultid="3610" />
                    <RANKING order="8" place="8" resultid="3347" />
                    <RANKING order="9" place="9" resultid="3689" />
                    <RANKING order="10" place="10" resultid="3692" />
                    <RANKING order="11" place="11" resultid="3242" />
                    <RANKING order="12" place="-1" resultid="3709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                    <RANKING order="2" place="2" resultid="3448" />
                    <RANKING order="3" place="3" resultid="3648" />
                    <RANKING order="4" place="4" resultid="3481" />
                    <RANKING order="5" place="5" resultid="3758" />
                    <RANKING order="6" place="6" resultid="3253" />
                    <RANKING order="7" place="7" resultid="3318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3595" />
                    <RANKING order="2" place="2" resultid="3602" />
                    <RANKING order="3" place="3" resultid="3643" />
                    <RANKING order="4" place="4" resultid="3484" />
                    <RANKING order="5" place="5" resultid="3215" />
                    <RANKING order="6" place="-1" resultid="3542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="2" resultid="3640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3434" />
                    <RANKING order="2" place="-1" resultid="3789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1308" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1309" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1310" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3959" daytime="17:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3960" daytime="17:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3961" daytime="17:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3962" daytime="17:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3963" daytime="17:38" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1311" daytime="17:41" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1312" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1313" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="1314" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1315" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1316" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1317" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1318" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1320" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1321" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1322" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1323" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1324" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1325" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1326" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3964" daytime="17:41" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3044" daytime="17:44" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3045" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3046" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3047" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3673" />
                    <RANKING order="2" place="2" resultid="3285" />
                    <RANKING order="3" place="3" resultid="3518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3048" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3049" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3282" />
                    <RANKING order="2" place="2" resultid="3379" />
                    <RANKING order="3" place="3" resultid="3354" />
                    <RANKING order="4" place="4" resultid="3635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3050" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3051" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3539" />
                    <RANKING order="2" place="2" resultid="3251" />
                    <RANKING order="3" place="3" resultid="3268" />
                    <RANKING order="4" place="-1" resultid="3245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3052" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="3053" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3054" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3469" />
                    <RANKING order="2" place="2" resultid="3668" />
                    <RANKING order="3" place="-1" resultid="3716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3055" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3056" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3057" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3058" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3059" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3965" daytime="17:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3966" daytime="17:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3060" daytime="17:49" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3061" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3062" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3063" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3064" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="3065" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="3066" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="3067" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="3068" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="3069" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="3070" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="3071" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3072" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3073" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3074" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3075" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3967" daytime="17:49" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3076" daytime="17:52" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3077" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3078" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3079" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3080" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="3081" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3082" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3083" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3084" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3591" />
                    <RANKING order="2" place="2" resultid="3491" />
                    <RANKING order="3" place="3" resultid="3236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3085" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3086" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3087" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3088" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3089" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3090" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3091" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3968" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3969" daytime="17:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3092" daytime="17:58" gender="F" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3093" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3094" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="3095" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="3096" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3097" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="3098" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3099" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="3100" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="3101" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3102" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="3103" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3104" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3105" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3106" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3107" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3970" daytime="17:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3108" daytime="18:01" gender="M" number="18" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3109" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3110" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3111" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3112" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="3113" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3114" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3115" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3638" />
                    <RANKING order="2" place="2" resultid="3687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3116" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3117" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="3118" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3119" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3120" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3121" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3122" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3123" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3971" daytime="18:01" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3124" daytime="18:04" number="19" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3125" agemax="119" agemin="100" />
                <AGEGROUP agegroupid="3144" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3525" />
                    <RANKING order="2" place="2" resultid="3927" />
                    <RANKING order="3" place="3" resultid="3311" />
                    <RANKING order="4" place="4" resultid="3523" />
                    <RANKING order="5" place="5" resultid="3312" />
                    <RANKING order="6" place="6" resultid="3524" />
                    <RANKING order="7" place="-1" resultid="3528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3143" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3527" />
                    <RANKING order="2" place="2" resultid="3546" />
                    <RANKING order="3" place="3" resultid="3526" />
                    <RANKING order="4" place="4" resultid="3313" />
                    <RANKING order="5" place="5" resultid="3928" />
                    <RANKING order="6" place="6" resultid="3332" />
                    <RANKING order="7" place="7" resultid="3314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3142" agemax="239" agemin="200" />
                <AGEGROUP agegroupid="3141" agemax="279" agemin="240" />
                <AGEGROUP agegroupid="3140" agemax="-1" agemin="280" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3972" daytime="18:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3973" daytime="18:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3160" daytime="18:13" gender="F" number="20" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3167" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3168" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3748" />
                    <RANKING order="2" place="2" resultid="3503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3169" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3678" />
                    <RANKING order="2" place="2" resultid="3494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3170" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3457" />
                    <RANKING order="2" place="2" resultid="3696" />
                    <RANKING order="3" place="3" resultid="3260" />
                    <RANKING order="4" place="4" resultid="3721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3171" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3566" />
                    <RANKING order="2" place="2" resultid="3264" />
                    <RANKING order="3" place="3" resultid="3324" />
                    <RANKING order="4" place="4" resultid="3675" />
                    <RANKING order="5" place="-1" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3172" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3509" />
                    <RANKING order="2" place="2" resultid="3428" />
                    <RANKING order="3" place="3" resultid="3416" />
                    <RANKING order="4" place="4" resultid="3321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3173" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3174" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="3175" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="3176" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="3177" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3178" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3179" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3180" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3181" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3976" daytime="18:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3977" daytime="18:21" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3182" daytime="18:31" gender="M" number="21" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3183" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="3184" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3751" />
                    <RANKING order="2" place="2" resultid="3352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3185" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3666" />
                    <RANKING order="2" place="2" resultid="3784" />
                    <RANKING order="3" place="3" resultid="3392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3186" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3431" />
                    <RANKING order="2" place="2" resultid="3693" />
                    <RANKING order="3" place="3" resultid="3690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3187" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3204" />
                    <RANKING order="2" place="2" resultid="3425" />
                    <RANKING order="3" place="3" resultid="3380" />
                    <RANKING order="4" place="4" resultid="3355" />
                    <RANKING order="5" place="5" resultid="3254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3188" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3395" />
                    <RANKING order="2" place="2" resultid="3211" />
                    <RANKING order="3" place="3" resultid="3327" />
                    <RANKING order="4" place="4" resultid="3644" />
                    <RANKING order="5" place="5" resultid="3377" />
                    <RANKING order="6" place="6" resultid="3218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3189" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3580" />
                    <RANKING order="2" place="2" resultid="3371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3190" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3775" />
                    <RANKING order="2" place="2" resultid="3486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3191" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3641" />
                    <RANKING order="2" place="2" resultid="3512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3192" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3193" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="3194" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="3195" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="3196" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="3197" agemax="94" agemin="90" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3978" daytime="18:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3979" daytime="18:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3980" daytime="18:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="3261" name="Masters Łódź">
          <ATHLETES>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="503605600029" swrid="5464091" athleteid="3262">
              <RESULTS>
                <RESULT eventid="1215" points="167" swimtime="00:03:48.92" resultid="3263" heatid="3954" lane="8" entrytime="00:03:47.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:53.85" />
                    <SPLIT distance="150" swimtime="00:02:55.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="175" swimtime="00:07:01.96" resultid="3264" heatid="3977" lane="3" entrytime="00:07:17.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:36.86" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                    <SPLIT distance="200" swimtime="00:03:26.27" />
                    <SPLIT distance="250" swimtime="00:04:21.55" />
                    <SPLIT distance="300" swimtime="00:05:16.70" />
                    <SPLIT distance="350" swimtime="00:06:11.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3333" name="5 Styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Łatkowska" birthdate="1965-10-06" gender="F" nation="POL" athleteid="3337">
              <RESULTS>
                <RESULT eventid="1183" points="105" swimtime="00:00:51.67" resultid="3338" heatid="3949" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1247" points="148" swimtime="00:01:37.56" resultid="3339" heatid="3957" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Usielska" birthdate="1985-12-09" gender="F" nation="POL" athleteid="3362">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3363" heatid="3933" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1247" status="DNS" swimtime="00:00:00.00" resultid="3364" heatid="3957" lane="8" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Broniszewski" birthdate="1980-09-26" gender="M" nation="POL" athleteid="3356">
              <RESULTS>
                <RESULT eventid="1103" points="150" swimtime="00:00:39.35" resultid="3357" heatid="3939" lane="0" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Tomaszewski" birthdate="1976-01-26" gender="M" nation="POL" athleteid="3334">
              <RESULTS>
                <RESULT eventid="1103" points="154" swimtime="00:00:38.97" resultid="3335" heatid="3939" lane="8" entrytime="00:00:45.00" />
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1199" status="DSQ" swimtime="00:00:00.00" resultid="3336" heatid="3952" lane="6" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Pilarska" birthdate="1997-02-16" gender="F" nation="POL" swrid="4282150" athleteid="3360">
              <RESULTS>
                <RESULT eventid="1058" points="536" swimtime="00:00:29.13" resultid="3361" heatid="3932" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Dzikiewicz" birthdate="1990-10-27" gender="M" nation="POL" athleteid="3348">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="3349" heatid="3938" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Kamiński" birthdate="1986-11-02" gender="M" nation="POL" athleteid="3345">
              <RESULTS>
                <RESULT eventid="1199" points="140" swimtime="00:00:42.82" resultid="3346" heatid="3952" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1295" points="212" swimtime="00:01:18.60" resultid="3347" heatid="3961" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-04-02" gender="M" nation="POL" swrid="4273597" athleteid="3365">
              <RESULTS>
                <RESULT eventid="3108" points="338" swimtime="00:01:11.02" resultid="3367" heatid="3971" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="378" swimtime="00:00:30.80" resultid="3929" heatid="3951" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Korzeniowski" birthdate="1985-07-09" gender="M" nation="POL" swrid="4042751" athleteid="3358">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters" eventid="1199" points="725" swimtime="00:00:24.78" resultid="3359" heatid="3950" lane="4" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Iwanowski" birthdate="1980-03-30" gender="M" nation="POL" athleteid="3353">
              <RESULTS>
                <RESULT eventid="3044" points="276" swimtime="00:01:27.29" resultid="3354" heatid="3965" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="172" swimtime="00:06:35.32" resultid="3355" heatid="3979" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:02:19.25" />
                    <SPLIT distance="200" swimtime="00:03:09.60" />
                    <SPLIT distance="250" swimtime="00:04:01.32" />
                    <SPLIT distance="300" swimtime="00:04:53.49" />
                    <SPLIT distance="350" swimtime="00:05:45.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Błażkiewicz" birthdate="1986-06-11" gender="F" nation="POL" athleteid="3342">
              <RESULTS>
                <RESULT eventid="1058" points="264" swimtime="00:00:36.87" resultid="3343" heatid="3933" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1151" points="214" swimtime="00:00:45.05" resultid="3344" heatid="3945" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Miśkiewicz" birthdate="1985-12-03" gender="F" nation="POL" athleteid="3340">
              <RESULTS>
                <RESULT eventid="1058" points="127" swimtime="00:00:47.05" resultid="3341" heatid="3934" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="1151" points="100" swimtime="00:00:57.96" resultid="3931" heatid="3945" lane="0" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="3350">
              <RESULTS>
                <RESULT eventid="3182" points="318" swimtime="00:05:22.37" resultid="3352" heatid="3978" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:55.71" />
                    <SPLIT distance="200" swimtime="00:02:36.87" />
                    <SPLIT distance="250" swimtime="00:03:17.76" />
                    <SPLIT distance="300" swimtime="00:03:59.96" />
                    <SPLIT distance="350" swimtime="00:04:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="336" swimtime="00:01:07.43" resultid="3930" heatid="3959" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="3124" points="396" swimtime="00:02:14.52" resultid="3927" heatid="3973" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:01:44.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3342" number="1" />
                    <RELAYPOSITION athleteid="3365" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3358" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3360" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="3124" points="157" swimtime="00:03:03.01" resultid="3928" heatid="3973" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:42.02" />
                    <SPLIT distance="150" swimtime="00:02:23.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3337" number="1" />
                    <RELAYPOSITION athleteid="3340" number="2" />
                    <RELAYPOSITION athleteid="3345" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3334" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" clubid="3219" name="Uks Delfin Legionowo">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Perl" birthdate="1996-06-07" gender="M" nation="POL" license="101414700068" swrid="4282344" athleteid="3223">
              <RESULTS>
                <RESULT eventid="1103" points="603" swimtime="00:00:24.75" resultid="3224" heatid="3935" lane="4" entrytime="00:00:23.00" />
                <RESULT eventid="1135" points="561" swimtime="00:00:31.46" resultid="3225" heatid="3942" lane="4" entrytime="00:00:28.96" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andzrej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" license="101414700141" athleteid="3220">
              <RESULTS>
                <RESULT eventid="1103" points="288" swimtime="00:00:31.66" resultid="3221" heatid="3937" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="3076" points="221" swimtime="00:01:25.75" resultid="3222" heatid="3968" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="3574" name="Stowarzyszenie Pływackie MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" athleteid="3578">
              <RESULTS>
                <RESULT eventid="1199" points="173" swimtime="00:00:39.95" resultid="3579" heatid="3953" lane="5" />
                <RESULT eventid="3182" points="175" swimtime="00:06:32.90" resultid="3580" heatid="3980" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:32.77" />
                    <SPLIT distance="150" swimtime="00:02:23.16" />
                    <SPLIT distance="200" swimtime="00:03:14.16" />
                    <SPLIT distance="250" swimtime="00:04:04.44" />
                    <SPLIT distance="300" swimtime="00:04:55.52" />
                    <SPLIT distance="350" swimtime="00:05:47.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-03-13" gender="M" nation="POL" license="103503700029" athleteid="3575">
              <RESULTS>
                <RESULT eventid="1103" points="379" swimtime="00:00:28.88" resultid="3576" heatid="3940" lane="8" />
                <RESULT eventid="1199" points="287" swimtime="00:00:33.73" resultid="3577" heatid="3952" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="09514" nation="POL" region="14" clubid="3592" name="UKP ,,Polonia Warszawa&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Rybiński" birthdate="1975-06-10" gender="M" nation="POL" license="509514700463" swrid="5240950" athleteid="3593">
              <RESULTS>
                <RESULT eventid="1135" points="269" swimtime="00:00:40.15" resultid="3594" heatid="3944" lane="4" />
                <RESULT eventid="1295" points="297" swimtime="00:01:10.27" resultid="3595" heatid="3962" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" clubid="3209" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Kowalczyk" birthdate="1974-10-02" gender="M" nation="POL" swrid="4992788" athleteid="3210">
              <RESULTS>
                <RESULT eventid="3182" points="382" swimtime="00:05:03.06" resultid="3211" heatid="3978" lane="6" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                    <SPLIT distance="200" swimtime="00:02:30.22" />
                    <SPLIT distance="250" swimtime="00:03:08.95" />
                    <SPLIT distance="300" swimtime="00:03:48.06" />
                    <SPLIT distance="350" swimtime="00:04:27.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3265" name="Niezrzeszeni KU AZS Politechnika Gdańska">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Nadolski" birthdate="1977-10-10" gender="M" nation="POL" athleteid="3280">
              <RESULTS>
                <RESULT eventid="1135" points="350" swimtime="00:00:36.81" resultid="3281" heatid="3942" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="3044" points="310" swimtime="00:01:24.03" resultid="3282" heatid="3965" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Rudzki" birthdate="1983-06-13" gender="M" nation="POL" athleteid="3292" />
            <ATHLETE firstname="Szymon" lastname="Kowalski" birthdate="1995-08-30" gender="M" nation="POL" swrid="4104892" athleteid="3305">
              <RESULTS>
                <RESULT eventid="1167" points="464" swimtime="00:00:31.00" resultid="3306" heatid="3947" lane="5" entrytime="00:00:29.88" />
                <RESULT eventid="3076" points="373" swimtime="00:01:11.97" resultid="3307" heatid="3968" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Miszewska" birthdate="1986-07-12" gender="F" nation="POL" athleteid="3289">
              <RESULTS>
                <RESULT eventid="1058" points="292" swimtime="00:00:35.67" resultid="3290" heatid="3933" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1183" points="265" swimtime="00:00:38.02" resultid="3291" heatid="3949" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Stankiewicz" birthdate="1969-03-01" gender="F" nation="POL" athleteid="3293">
              <RESULTS>
                <RESULT eventid="1247" points="189" swimtime="00:01:30.07" resultid="3294" heatid="3958" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="162" swimtime="00:07:13.23" resultid="3295" heatid="3977" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="100" swimtime="00:01:34.96" />
                    <SPLIT distance="150" swimtime="00:02:29.99" />
                    <SPLIT distance="200" swimtime="00:03:26.92" />
                    <SPLIT distance="250" swimtime="00:04:23.57" />
                    <SPLIT distance="300" swimtime="00:05:21.05" />
                    <SPLIT distance="350" swimtime="00:06:19.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Węckowicz" birthdate="1983-05-24" gender="M" nation="POL" athleteid="3299">
              <RESULTS>
                <RESULT eventid="1103" points="404" swimtime="00:00:28.28" resultid="3300" heatid="3936" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1295" points="384" swimtime="00:01:04.52" resultid="3301" heatid="3959" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Jakóbczyk" birthdate="1993-04-13" gender="F" nation="POL" swrid="4086939" athleteid="3274">
              <RESULTS>
                <RESULT eventid="1058" points="499" swimtime="00:00:29.84" resultid="3275" heatid="3932" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1183" points="402" swimtime="00:00:33.08" resultid="3276" heatid="3949" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Remizowicz" birthdate="1984-09-23" gender="M" nation="POL" athleteid="3286">
              <RESULTS>
                <RESULT eventid="1103" points="336" swimtime="00:00:30.07" resultid="3287" heatid="3937" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1295" points="328" swimtime="00:01:08.02" resultid="3288" heatid="3959" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wawrzyniec" lastname="Rawicz-Zegrzda" birthdate="1987-02-28" gender="M" nation="POL" athleteid="3283">
              <RESULTS>
                <RESULT eventid="1295" points="171" swimtime="00:01:24.46" resultid="3284" heatid="3962" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3044" points="190" swimtime="00:01:38.87" resultid="3285" heatid="3966" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Gawarkiewicz" birthdate="1973-06-03" gender="M" nation="POL" athleteid="3271">
              <RESULTS>
                <RESULT eventid="1135" points="238" swimtime="00:00:41.86" resultid="3272" heatid="3943" lane="7" />
                <RESULT eventid="1199" points="128" swimtime="00:00:44.17" resultid="3273" heatid="3952" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Abramski" birthdate="1971-07-10" gender="M" nation="POL" athleteid="3266">
              <RESULTS>
                <RESULT eventid="1135" points="102" swimtime="00:00:55.52" resultid="3267" heatid="3943" lane="1" />
                <RESULT eventid="3044" points="92" swimtime="00:02:05.58" resultid="3268" heatid="3966" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Janowicz" birthdate="1977-04-12" gender="M" nation="POL" athleteid="3277">
              <RESULTS>
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="3278" heatid="3943" lane="5" />
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="3279" heatid="3953" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Maciesza" birthdate="1996-03-20" gender="F" nation="POL" swrid="4157882" athleteid="3308">
              <RESULTS>
                <RESULT eventid="1119" points="365" swimtime="00:00:41.13" resultid="3309" heatid="3941" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1183" points="429" swimtime="00:00:32.38" resultid="3310" heatid="3949" lane="4" entrytime="00:00:31.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Żylewicz" birthdate="1989-11-26" gender="M" nation="POL" athleteid="3302">
              <RESULTS>
                <RESULT eventid="1103" points="337" swimtime="00:00:30.03" resultid="3303" heatid="3937" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1295" points="311" swimtime="00:01:09.23" resultid="3304" heatid="3960" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Wasilczuk" birthdate="1962-05-10" gender="M" nation="POL" athleteid="3296">
              <RESULTS>
                <RESULT eventid="1103" points="100" swimtime="00:00:44.99" resultid="3297" heatid="3940" lane="1" />
                <RESULT eventid="1135" points="95" swimtime="00:00:56.79" resultid="3298" heatid="3943" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Borucka" birthdate="1975-10-07" gender="F" nation="POL" athleteid="3269">
              <RESULTS>
                <RESULT eventid="1058" points="53" swimtime="00:01:02.93" resultid="3270" heatid="3934" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="3124" points="379" swimtime="00:02:16.47" resultid="3311" heatid="3972" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:45.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3274" number="1" />
                    <RELAYPOSITION athleteid="3280" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3299" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3302" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="3124" points="267" swimtime="00:02:33.41" resultid="3312" heatid="3972" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:18.88" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3286" number="1" />
                    <RELAYPOSITION athleteid="3283" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3308" number="3" />
                    <RELAYPOSITION athleteid="3292" number="4" reactiontime="+99" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="3124" points="167" swimtime="00:02:59.37" resultid="3313" heatid="3972" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:21.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3289" number="1" />
                    <RELAYPOSITION athleteid="3296" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3271" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3293" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="3124" points="131" swimtime="00:03:14.18" resultid="3314" heatid="3973" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                    <SPLIT distance="150" swimtime="00:02:09.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3305" number="1" />
                    <RELAYPOSITION athleteid="3266" number="2" />
                    <RELAYPOSITION athleteid="3277" number="3" />
                    <RELAYPOSITION athleteid="3269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3233" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" athleteid="3234">
              <RESULTS>
                <RESULT eventid="1103" points="128" swimtime="00:00:41.44" resultid="3235" heatid="3939" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="3076" points="103" swimtime="00:01:50.57" resultid="3236" heatid="3968" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Romiszowski" birthdate="1983-02-14" gender="M" nation="POL" athleteid="3246">
              <RESULTS>
                <RESULT eventid="1103" points="266" swimtime="00:00:32.51" resultid="3247" heatid="3936" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1295" points="233" swimtime="00:01:16.14" resultid="3248" heatid="3960" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Buczyńska" birthdate="2001-02-15" gender="F" nation="POL" athleteid="3255">
              <RESULTS>
                <RESULT eventid="1058" points="278" swimtime="00:00:36.24" resultid="3256" heatid="3933" lane="6" entrytime="00:00:37.42" />
                <RESULT eventid="1247" points="248" swimtime="00:01:22.21" resultid="3257" heatid="3957" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Ostapczuk" birthdate="1970-07-13" gender="M" nation="POL" athleteid="3243">
              <RESULTS>
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3244" heatid="3961" lane="7" entrytime="00:01:29.00" />
                <RESULT eventid="3044" status="DNS" swimtime="00:00:00.00" resultid="3245" heatid="3965" lane="7" entrytime="00:01:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="3543">
              <RESULTS>
                <RESULT eventid="1199" points="160" swimtime="00:00:40.98" resultid="3544" heatid="3953" lane="3" />
                <RESULT eventid="3108" points="110" swimtime="00:01:43.18" resultid="3545" heatid="3971" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kosiela" birthdate="1985-02-03" gender="M" nation="POL" athleteid="3240">
              <RESULTS>
                <RESULT eventid="1199" points="145" swimtime="00:00:42.30" resultid="3241" heatid="3951" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1295" points="156" swimtime="00:01:26.97" resultid="3242" heatid="3960" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Prugar-Fukowska" birthdate="1983-05-28" gender="F" nation="POL" athleteid="3258">
              <RESULTS>
                <RESULT eventid="1247" points="185" swimtime="00:01:30.62" resultid="3259" heatid="3957" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="211" swimtime="00:06:37.07" resultid="3260" heatid="3977" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                    <SPLIT distance="100" swimtime="00:01:34.00" />
                    <SPLIT distance="150" swimtime="00:02:25.31" />
                    <SPLIT distance="200" swimtime="00:03:15.94" />
                    <SPLIT distance="250" swimtime="00:04:06.30" />
                    <SPLIT distance="300" swimtime="00:04:56.83" />
                    <SPLIT distance="350" swimtime="00:05:46.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Siergiej" lastname="Kulinicz" birthdate="1986-05-08" gender="M" nation="POL" license="510414700071" swrid="5471787" athleteid="3532">
              <RESULTS>
                <RESULT eventid="1103" points="335" swimtime="00:00:30.08" resultid="3533" heatid="3936" lane="8" entrytime="00:00:29.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="510414600003" swrid="5240601" athleteid="3534">
              <RESULTS>
                <RESULT eventid="1119" points="432" swimtime="00:00:38.88" resultid="3535" heatid="3941" lane="3" entrytime="00:00:39.14" entrycourse="LCM" />
                <RESULT eventid="1311" points="377" swimtime="00:01:28.72" resultid="3536" heatid="3964" lane="4" entrytime="00:01:31.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Januszewski" birthdate="1970-08-05" gender="M" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1103" points="137" swimtime="00:00:40.56" resultid="3250" heatid="3939" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="3044" points="130" swimtime="00:01:52.28" resultid="3251" heatid="3965" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Cybulski" birthdate="1972-08-08" gender="M" nation="POL" license="510414700015" athleteid="3540">
              <RESULTS>
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="3541" heatid="3943" lane="3" />
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3542" heatid="3963" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Olesiński" birthdate="1980-11-25" gender="M" nation="POL" athleteid="3252">
              <RESULTS>
                <RESULT eventid="1295" points="146" swimtime="00:01:29.01" resultid="3253" heatid="3961" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="114" swimtime="00:07:32.81" resultid="3254" heatid="3979" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:38.33" />
                    <SPLIT distance="200" swimtime="00:03:34.71" />
                    <SPLIT distance="250" swimtime="00:04:33.90" />
                    <SPLIT distance="300" swimtime="00:05:32.64" />
                    <SPLIT distance="350" swimtime="00:06:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="3537">
              <RESULTS>
                <RESULT eventid="1135" points="195" swimtime="00:00:44.74" resultid="3538" heatid="3942" lane="8" entrytime="00:00:45.48" entrycourse="LCM" />
                <RESULT eventid="3044" points="157" swimtime="00:01:45.33" resultid="3539" heatid="3965" lane="8" entrytime="00:01:45.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="3124" points="218" swimtime="00:02:44.08" resultid="3546" heatid="3973" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3246" number="1" />
                    <RELAYPOSITION athleteid="3534" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="3240" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="3258" number="4" reactiontime="+96" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06414" nation="POL" region="14" clubid="3567" name="MKS Piaseczno">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Susabowski" birthdate="1981-05-02" gender="M" nation="POL" license="506414700267" athleteid="3572">
              <RESULTS>
                <RESULT eventid="1199" points="218" swimtime="00:00:36.95" resultid="3573" heatid="3952" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Turczyński" birthdate="1979-02-21" gender="M" nation="POL" license="300714700065" athleteid="3570">
              <RESULTS>
                <RESULT eventid="1103" points="543" swimtime="00:00:25.63" resultid="3571" heatid="3935" lane="5" entrytime="00:00:25.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Szpala" birthdate="1975-11-23" gender="F" nation="POL" license="506414600256" athleteid="3568">
              <RESULTS>
                <RESULT eventid="1058" points="94" swimtime="00:00:51.92" resultid="3569" heatid="3934" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="14" clubid="3556" name="Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Wilczęga" birthdate="1981-10-24" gender="M" nation="POL" license="106614700042" swrid="4992879" athleteid="3557">
              <RESULTS>
                <RESULT eventid="1103" points="455" swimtime="00:00:27.18" resultid="3558" heatid="3935" lane="1" entrytime="00:00:26.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASBYD" nation="POL" region="02" clubid="3914" name=" Astoria Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Michałowska" gender="F" nation="POL" athleteid="3913">
              <RESULTS>
                <RESULT eventid="1247" points="412" swimtime="00:01:09.46" resultid="3915" heatid="3958" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="337" swimtime="00:01:22.72" resultid="3924" heatid="3967" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="3612" name="UKS ,,Trójka&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="3613">
              <RESULTS>
                <RESULT eventid="1231" points="333" swimtime="00:02:44.46" resultid="3614" heatid="3956" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:02:06.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3044" status="DNS" swimtime="00:00:00.00" resultid="3615" heatid="3966" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00306" nation="POL" region="06" clubid="3552" name="KS Korona Kraków">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" license="500306600160" swrid="4992827" athleteid="3553">
              <RESULTS>
                <RESULT eventid="1215" points="257" swimtime="00:03:18.28" resultid="3554" heatid="3954" lane="6" entrytime="00:03:18.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:34.65" />
                    <SPLIT distance="150" swimtime="00:02:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3092" points="217" swimtime="00:01:32.29" resultid="3555" heatid="3970" lane="5" entrytime="00:01:32.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03114" nation="POL" region="14" clubid="3596" name="Uks ,,Pingwiny&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Karol" lastname="Perl" birthdate="1976-11-03" gender="M" nation="POL" license="103114700212" swrid="5120236" athleteid="3600">
              <RESULTS>
                <RESULT eventid="1103" points="313" swimtime="00:00:30.79" resultid="3601" heatid="3940" lane="3" />
                <RESULT eventid="1295" points="294" swimtime="00:01:10.52" resultid="3602" heatid="3962" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Kostanowicz" birthdate="1998-04-03" gender="M" nation="POL" license="103114700307" swrid="4363163" athleteid="3606">
              <RESULTS>
                <RESULT eventid="1231" points="361" swimtime="00:02:40.08" resultid="3607" heatid="3956" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:02:02.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3076" points="464" swimtime="00:01:06.96" resultid="3608" heatid="3968" lane="4" entrytime="00:01:00.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Bocianiak" birthdate="1988-04-22" gender="F" nation="POL" license="503114600308" athleteid="3597">
              <RESULTS>
                <RESULT eventid="1058" points="332" swimtime="00:00:34.18" resultid="3598" heatid="3934" lane="8" />
                <RESULT eventid="1183" points="256" swimtime="00:00:38.43" resultid="3599" heatid="3949" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Żarłok" birthdate="1983-09-26" gender="M" nation="POL" license="103114700213" athleteid="3609">
              <RESULTS>
                <RESULT eventid="1295" points="217" swimtime="00:01:18.04" resultid="3610" heatid="3962" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3044" points="175" swimtime="00:01:41.56" resultid="3611" heatid="3966" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Pawlak" birthdate="2001-04-17" gender="M" nation="POL" license="503114700309" swrid="4580147" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1103" points="392" swimtime="00:00:28.56" resultid="3604" heatid="3940" lane="7" />
                <RESULT eventid="1135" points="274" swimtime="00:00:39.92" resultid="3605" heatid="3943" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="3563" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-07-14" gender="F" nation="POL" license="500309600228" swrid="4595750" athleteid="3564">
              <RESULTS>
                <RESULT eventid="1215" points="389" swimtime="00:02:52.63" resultid="3565" heatid="3954" lane="5" entrytime="00:02:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:12.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="432" swimtime="00:05:12.64" resultid="3566" heatid="3976" lane="5" entrytime="00:05:23.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:52.21" />
                    <SPLIT distance="200" swimtime="00:02:32.39" />
                    <SPLIT distance="250" swimtime="00:03:13.20" />
                    <SPLIT distance="300" swimtime="00:03:53.80" />
                    <SPLIT distance="350" swimtime="00:04:34.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11514" nation="POL" region="14" clubid="3581" name="Stowarzyszenie Pływackie Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Łukasiuk" birthdate="1980-01-02" gender="F" nation="POL" license="511514600187" athleteid="3582">
              <RESULTS>
                <RESULT eventid="1058" points="394" swimtime="00:00:32.27" resultid="3583" heatid="3934" lane="0" />
                <RESULT eventid="1119" points="349" swimtime="00:00:41.73" resultid="3584" heatid="3941" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Fuliński" birthdate="1982-06-03" gender="M" nation="POL" license="111514700186" swrid="4992686" athleteid="3585">
              <RESULTS>
                <RESULT eventid="1103" points="480" swimtime="00:00:26.70" resultid="3586" heatid="3940" lane="2" />
                <RESULT eventid="1295" points="502" swimtime="00:00:58.99" resultid="3587" heatid="3962" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="3645" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" swrid="5416809" athleteid="3646">
              <RESULTS>
                <RESULT eventid="1103" points="304" swimtime="00:00:31.08" resultid="3647" heatid="3937" lane="0" entrytime="00:00:31.48" entrycourse="LCM" />
                <RESULT eventid="1295" points="302" swimtime="00:01:09.88" resultid="3648" heatid="3960" lane="2" entrytime="00:01:12.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="3649">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski Masters" eventid="1135" points="421" swimtime="00:00:34.62" resultid="3650" heatid="3944" lane="3" />
                <RESULT eventid="1295" points="344" swimtime="00:01:06.93" resultid="3651" heatid="3962" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" swrid="5471789" athleteid="3658">
              <RESULTS>
                <RESULT eventid="1231" points="355" swimtime="00:02:40.97" resultid="3659" heatid="3956" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3108" points="363" swimtime="00:01:09.35" resultid="3660" heatid="3971" lane="4" entrytime="00:01:08.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" swrid="4043251" athleteid="3652">
              <RESULTS>
                <RESULT eventid="1167" points="613" swimtime="00:00:28.25" resultid="3653" heatid="3948" lane="3" />
                <RESULT eventid="1199" points="554" swimtime="00:00:27.11" resultid="3654" heatid="3952" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="3655">
              <RESULTS>
                <RESULT eventid="1167" points="152" swimtime="00:00:44.95" resultid="3656" heatid="3948" lane="6" />
                <RESULT eventid="3076" points="147" swimtime="00:01:38.09" resultid="3657" heatid="3968" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Miński" birthdate="1956-01-14" gender="M" nation="POL" license="512914700021" swrid="4754653" athleteid="3667">
              <RESULTS>
                <RESULT eventid="3044" points="80" swimtime="00:02:11.61" resultid="3668" heatid="3966" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kotlarski" birthdate="1989-05-02" gender="M" nation="POL" license="512914700025" swrid="4071566" athleteid="3664">
              <RESULTS>
                <RESULT eventid="1231" points="401" swimtime="00:02:34.53" resultid="3665" heatid="3956" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:59.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="398" swimtime="00:04:59.10" resultid="3666" heatid="3980" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:10.25" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                    <SPLIT distance="200" swimtime="00:02:27.42" />
                    <SPLIT distance="250" swimtime="00:03:05.68" />
                    <SPLIT distance="300" swimtime="00:03:45.00" />
                    <SPLIT distance="350" swimtime="00:04:23.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" swrid="5312396" athleteid="3661">
              <RESULTS>
                <RESULT eventid="1231" points="324" swimtime="00:02:45.85" resultid="3662" heatid="3956" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:17.37" />
                    <SPLIT distance="150" swimtime="00:02:07.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3076" points="324" swimtime="00:01:15.44" resultid="3663" heatid="3968" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PASPO" nation="POL" region="14" clubid="3907" name="Parasportowi">
          <ATHLETES>
            <ATHLETE firstname="Oliwia" lastname="Szadkowska" gender="F" nation="POL" athleteid="3918">
              <RESULTS>
                <RESULT eventid="1247" points="104" swimtime="00:01:49.88" resultid="3919" heatid="3958" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="80" swimtime="00:02:13.51" resultid="3926" heatid="3967" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Perkowski" gender="F" nation="POL" athleteid="3909">
              <RESULTS>
                <RESULT eventid="1247" points="188" swimtime="00:01:30.22" resultid="3910" heatid="3958" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="146" swimtime="00:01:49.26" resultid="3922" heatid="3967" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Mroziński" gender="F" nation="POL" athleteid="3906">
              <RESULTS>
                <RESULT eventid="1247" points="89" swimtime="00:01:55.78" resultid="3908" heatid="3958" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="97" swimtime="00:02:05.02" resultid="3921" heatid="3967" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Urbański" gender="F" nation="POL" athleteid="3911">
              <RESULTS>
                <RESULT eventid="1247" points="374" swimtime="00:01:11.75" resultid="3912" heatid="3958" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="220" swimtime="00:01:35.26" resultid="3923" heatid="3967" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natasza" lastname="Jaworska " gender="F" nation="POL" athleteid="3916">
              <RESULTS>
                <RESULT eventid="1247" points="76" swimtime="00:02:01.73" resultid="3917" heatid="3958" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3060" points="72" swimtime="00:02:18.09" resultid="3925" heatid="3967" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03508" nation="POL" region="08" clubid="3548" name="Ks &quot;Prestige&quot;">
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Rupa" birthdate="1996-01-11" gender="F" nation="POL" license="103508600006" swrid="4108567" athleteid="3549">
              <RESULTS>
                <RESULT eventid="1151" points="493" swimtime="00:00:34.13" resultid="3550" heatid="3945" lane="5" entrytime="00:00:34.24" entrycourse="LCM" />
                <RESULT eventid="3060" points="473" swimtime="00:01:13.84" resultid="3551" heatid="3967" lane="4" entrytime="00:01:15.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="11" clubid="3616" name="UKS Trójka">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" swrid="4762175" athleteid="3617">
              <RESULTS>
                <RESULT eventid="1103" points="559" swimtime="00:00:25.38" resultid="3618" heatid="3935" lane="3" entrytime="00:00:25.35" entrycourse="LCM" />
                <RESULT eventid="1199" points="569" swimtime="00:00:26.86" resultid="3619" heatid="3950" lane="5" entrytime="00:00:27.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kozioł" birthdate="1990-08-26" gender="M" nation="POL" license="100111700090" swrid="4112682" athleteid="3623">
              <RESULTS>
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="3624" heatid="3950" lane="7" entrytime="00:00:30.29" entrycourse="SCM" />
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3625" heatid="3963" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Chowaniec" birthdate="1995-06-07" gender="M" nation="POL" license="100111700079" swrid="5265087" athleteid="3620">
              <RESULTS>
                <RESULT eventid="1135" points="520" swimtime="00:00:32.26" resultid="3621" heatid="3942" lane="5" entrytime="00:00:31.57" entrycourse="LCM" />
                <RESULT eventid="1231" points="460" swimtime="00:02:27.66" resultid="3622" heatid="3955" lane="5" entrytime="00:02:30.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:52.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="102705" nation="POL" clubid="3315" name="Olimpijczy Tomaszów Maz.">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Bucholz" birthdate="1972-01-26" gender="M" nation="POL" swrid="4754642" athleteid="3325">
              <RESULTS>
                <RESULT eventid="1231" points="216" swimtime="00:03:09.80" resultid="3326" heatid="3955" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                    <SPLIT distance="150" swimtime="00:02:23.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="251" swimtime="00:05:48.68" resultid="3327" heatid="3978" lane="9" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:02.29" />
                    <SPLIT distance="200" swimtime="00:02:47.60" />
                    <SPLIT distance="250" swimtime="00:03:33.28" />
                    <SPLIT distance="300" swimtime="00:04:18.59" />
                    <SPLIT distance="350" swimtime="00:05:05.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bucholz" birthdate="1973-12-01" gender="F" nation="POL" license="502705600074" swrid="4919376" athleteid="3319">
              <RESULTS>
                <RESULT eventid="1215" points="86" swimtime="00:04:45.12" resultid="3320" heatid="3954" lane="9" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.29" />
                    <SPLIT distance="100" swimtime="00:02:21.41" />
                    <SPLIT distance="150" swimtime="00:03:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="100" swimtime="00:08:28.93" resultid="3321" heatid="3977" lane="7" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.07" />
                    <SPLIT distance="100" swimtime="00:01:54.02" />
                    <SPLIT distance="150" swimtime="00:02:58.59" />
                    <SPLIT distance="200" swimtime="00:04:05.27" />
                    <SPLIT distance="250" swimtime="00:05:11.78" />
                    <SPLIT distance="300" swimtime="00:06:19.16" />
                    <SPLIT distance="350" swimtime="00:07:25.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Kozłowska" birthdate="1979-03-01" gender="F" nation="POL" license="502705600074" swrid="4992866" athleteid="3322">
              <RESULTS>
                <RESULT eventid="1215" points="160" swimtime="00:03:52.28" resultid="3323" heatid="3954" lane="1" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:52.81" />
                    <SPLIT distance="150" swimtime="00:02:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="156" swimtime="00:07:18.96" resultid="3324" heatid="3977" lane="6" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:35.24" />
                    <SPLIT distance="150" swimtime="00:02:31.27" />
                    <SPLIT distance="200" swimtime="00:03:30.43" />
                    <SPLIT distance="250" swimtime="00:04:30.06" />
                    <SPLIT distance="300" swimtime="00:05:29.85" />
                    <SPLIT distance="350" swimtime="00:06:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartek" lastname="Masłocha" birthdate="1979-01-23" gender="M" nation="POL" license="502705700076" athleteid="3316">
              <RESULTS>
                <RESULT eventid="1167" points="135" swimtime="00:00:46.71" resultid="3317" heatid="3948" lane="5" entrytime="00:01:09.00" />
                <RESULT eventid="1295" points="128" swimtime="00:01:32.88" resultid="3318" heatid="3962" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="3124" points="155" swimtime="00:03:03.61" resultid="3332" heatid="3973" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:48.00" />
                    <SPLIT distance="150" swimtime="00:02:24.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3316" number="1" />
                    <RELAYPOSITION athleteid="3319" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3325" number="3" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3322" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TK" nation="POL" clubid="3212" name="Team Karaś">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" athleteid="3216">
              <RESULTS>
                <RESULT eventid="1231" points="92" swimtime="00:04:12.02" resultid="3217" heatid="3955" lane="9" entrytime="00:04:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.73" />
                    <SPLIT distance="100" swimtime="00:02:07.46" />
                    <SPLIT distance="150" swimtime="00:03:20.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="114" swimtime="00:07:33.10" resultid="3218" heatid="3979" lane="0" entrytime="00:07:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:38.10" />
                    <SPLIT distance="150" swimtime="00:02:35.26" />
                    <SPLIT distance="200" swimtime="00:03:34.00" />
                    <SPLIT distance="250" swimtime="00:04:35.39" />
                    <SPLIT distance="300" swimtime="00:05:35.97" />
                    <SPLIT distance="350" swimtime="00:06:36.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" athleteid="3213">
              <RESULTS>
                <RESULT eventid="1103" points="195" swimtime="00:00:36.02" resultid="3214" heatid="3938" lane="9" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1295" points="182" swimtime="00:01:22.65" resultid="3215" heatid="3960" lane="3" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3670" name="Zawodnicy niezrzeszeni">
          <ATHLETES>
            <ATHLETE firstname="Sławek" lastname="Kacprowicz" birthdate="1958-06-15" gender="M" nation="POL" athleteid="3711">
              <RESULTS>
                <RESULT eventid="1135" points="39" swimtime="00:01:16.42" resultid="3712" heatid="3943" lane="4" entrytime="00:01:15.00" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="3044" status="DSQ" swimtime="00:03:11.57" resultid="3713" heatid="3966" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Baltaza" birthdate="1999-04-13" gender="M" nation="POL" swrid="4418613" athleteid="3740">
              <RESULTS>
                <RESULT eventid="1103" points="555" swimtime="00:00:25.44" resultid="3741" heatid="3937" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="3742" heatid="3950" lane="9" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Malczewska" birthdate="2000-06-26" gender="F" nation="POL" swrid="4585023" athleteid="3734">
              <RESULTS>
                <RESULT eventid="1058" points="488" swimtime="00:00:30.06" resultid="3735" heatid="3932" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1151" points="453" swimtime="00:00:35.11" resultid="3736" heatid="3945" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Fojudzki" birthdate="1982-05-31" gender="M" nation="POL" athleteid="3708">
              <RESULTS>
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3709" heatid="3960" lane="6" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Swianiewicz" birthdate="1985-06-28" gender="M" nation="POL" athleteid="3691">
              <RESULTS>
                <RESULT eventid="1295" points="183" swimtime="00:01:22.51" resultid="3692" heatid="3960" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="185" swimtime="00:06:25.85" resultid="3693" heatid="3979" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:16.59" />
                    <SPLIT distance="200" swimtime="00:03:06.82" />
                    <SPLIT distance="250" swimtime="00:03:57.34" />
                    <SPLIT distance="300" swimtime="00:04:47.49" />
                    <SPLIT distance="350" swimtime="00:05:37.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Wasiuk" birthdate="1953-09-27" gender="M" nation="POL" swrid="4313185" athleteid="3705">
              <RESULTS>
                <RESULT eventid="1231" points="74" swimtime="00:04:30.86" resultid="3706" heatid="3956" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:02:16.58" />
                    <SPLIT distance="150" swimtime="00:03:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3108" points="53" swimtime="00:02:11.58" resultid="3707" heatid="3971" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Stachera" birthdate="1995-07-11" gender="M" nation="POL" athleteid="3682">
              <RESULTS>
                <RESULT eventid="1103" points="412" swimtime="00:00:28.08" resultid="3683" heatid="3935" lane="0" entrytime="00:00:28.50" />
                <RESULT eventid="1167" points="316" swimtime="00:00:35.21" resultid="3684" heatid="3947" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jędrzej" lastname="Sanok" birthdate="1989-02-24" gender="M" nation="POL" athleteid="3779">
              <RESULTS>
                <RESULT eventid="1199" points="332" swimtime="00:00:32.15" resultid="3780" heatid="3951" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="3108" points="226" swimtime="00:01:21.15" resultid="3781" heatid="3971" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Mazur" birthdate="1958-12-23" gender="M" nation="POL" athleteid="3722">
              <RESULTS>
                <RESULT eventid="1103" points="98" swimtime="00:00:45.29" resultid="3723" heatid="3939" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1135" points="104" swimtime="00:00:55.03" resultid="3724" heatid="3942" lane="9" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Łasica" birthdate="1990-09-06" gender="F" nation="POL" athleteid="3770">
              <RESULTS>
                <RESULT eventid="1058" points="116" swimtime="00:00:48.47" resultid="3771" heatid="3934" lane="7" />
                <RESULT eventid="1151" points="114" swimtime="00:00:55.56" resultid="3772" heatid="3946" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Kukułka" birthdate="1978-12-05" gender="M" nation="POL" athleteid="3737">
              <RESULTS>
                <RESULT eventid="1103" points="279" swimtime="00:00:31.98" resultid="3738" heatid="3937" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1231" points="163" swimtime="00:03:28.61" resultid="3739" heatid="3955" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:43.01" />
                    <SPLIT distance="150" swimtime="00:02:42.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Rybicki" birthdate="1963-05-11" gender="M" nation="POL" swrid="4340488" athleteid="3765">
              <RESULTS>
                <RESULT eventid="1103" points="288" swimtime="00:00:31.64" resultid="3766" heatid="3937" lane="8" entrytime="00:00:31.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Cieślak" birthdate="1961-12-21" gender="M" nation="POL" athleteid="3794">
              <RESULTS>
                <RESULT eventid="1199" points="69" swimtime="00:00:54.07" resultid="3795" heatid="3952" lane="7" entrytime="00:01:00.00" />
                <RESULT eventid="1231" points="65" swimtime="00:04:42.90" resultid="3796" heatid="3955" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                    <SPLIT distance="100" swimtime="00:02:19.95" />
                    <SPLIT distance="150" swimtime="00:03:41.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Walerzak" birthdate="1978-09-23" gender="F" nation="POL" athleteid="3697">
              <RESULTS>
                <RESULT eventid="1119" points="190" swimtime="00:00:51.12" resultid="3698" heatid="3941" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1151" points="78" swimtime="00:01:03.08" resultid="3699" heatid="3945" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Janicka" birthdate="1984-04-18" gender="F" nation="POL" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1058" points="443" swimtime="00:00:31.05" resultid="3695" heatid="3932" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="3160" points="265" swimtime="00:06:07.82" resultid="3696" heatid="3976" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:02:10.27" />
                    <SPLIT distance="200" swimtime="00:02:57.85" />
                    <SPLIT distance="250" swimtime="00:03:45.89" />
                    <SPLIT distance="300" swimtime="00:04:35.03" />
                    <SPLIT distance="350" swimtime="00:05:23.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sabadasz" birthdate="1975-11-04" gender="M" nation="POL" athleteid="3725">
              <RESULTS>
                <RESULT eventid="1103" points="240" swimtime="00:00:33.64" resultid="3726" heatid="3938" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1199" points="181" swimtime="00:00:39.32" resultid="3727" heatid="3951" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Kotowska" birthdate="1980-12-11" gender="F" nation="POL" athleteid="3752">
              <RESULTS>
                <RESULT eventid="1119" points="178" swimtime="00:00:52.17" resultid="3753" heatid="3941" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Ogłoblin" birthdate="1992-02-27" gender="M" nation="POL" swrid="4806326" athleteid="3749">
              <RESULTS>
                <RESULT eventid="1295" points="430" swimtime="00:01:02.14" resultid="3750" heatid="3959" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="325" swimtime="00:05:19.98" resultid="3751" heatid="3978" lane="1" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:01:54.24" />
                    <SPLIT distance="200" swimtime="00:02:35.67" />
                    <SPLIT distance="250" swimtime="00:03:17.65" />
                    <SPLIT distance="300" swimtime="00:03:59.52" />
                    <SPLIT distance="350" swimtime="00:04:41.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Białek" birthdate="1989-08-25" gender="F" nation="POL" athleteid="3702">
              <RESULTS>
                <RESULT eventid="1151" points="147" swimtime="00:00:51.04" resultid="3703" heatid="3946" lane="3" />
                <RESULT eventid="3060" points="127" swimtime="00:01:54.27" resultid="3704" heatid="3967" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Zieliński" birthdate="1954-09-17" gender="M" nation="POL" athleteid="3788">
              <RESULTS>
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3789" heatid="3962" lane="5" entrytime="00:01:45.00" />
                <RESULT eventid="3076" status="DNS" swimtime="00:00:00.00" resultid="3790" heatid="3969" lane="4" entrytime="00:02:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kotowski" birthdate="1978-04-13" gender="M" nation="POL" athleteid="3756">
              <RESULTS>
                <RESULT eventid="1103" points="246" swimtime="00:00:33.37" resultid="3757" heatid="3938" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1295" points="245" swimtime="00:01:14.96" resultid="3758" heatid="3961" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jędrzej" lastname="Wengerski" birthdate="1992-07-25" gender="M" nation="POL" swrid="4112868" athleteid="3679">
              <RESULTS>
                <RESULT eventid="1103" points="513" swimtime="00:00:26.11" resultid="3680" heatid="3935" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1295" points="515" swimtime="00:00:58.52" resultid="3681" heatid="3959" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" swrid="4282341" athleteid="3731">
              <RESULTS>
                <RESULT eventid="1119" points="546" swimtime="00:00:35.97" resultid="3732" heatid="3941" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1183" points="442" swimtime="00:00:32.05" resultid="3733" heatid="3949" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Maścianica" birthdate="1985-04-17" gender="M" nation="POL" athleteid="3759">
              <RESULTS>
                <RESULT eventid="1103" points="357" swimtime="00:00:29.47" resultid="3760" heatid="3937" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1167" points="307" swimtime="00:00:35.57" resultid="3761" heatid="3947" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vasyl" lastname="Rybalka" birthdate="1985-09-25" gender="M" nation="POL" athleteid="3728">
              <RESULTS>
                <RESULT eventid="1199" points="435" swimtime="00:00:29.39" resultid="3729" heatid="3950" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1295" points="427" swimtime="00:01:02.27" resultid="3730" heatid="3959" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Kacprowicz" birthdate="1955-04-14" gender="M" nation="POL" athleteid="3714">
              <RESULTS>
                <RESULT eventid="1103" points="48" swimtime="00:00:57.18" resultid="3715" heatid="3939" lane="9" entrytime="00:00:58.00" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="3044" status="DSQ" swimtime="00:02:33.39" resultid="3716" heatid="3966" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Kaczmarek" birthdate="1976-11-27" gender="F" nation="POL" athleteid="3743">
              <RESULTS>
                <RESULT eventid="1058" points="77" swimtime="00:00:55.47" resultid="3744" heatid="3934" lane="3" />
                <RESULT eventid="1247" points="58" swimtime="00:02:13.28" resultid="3745" heatid="3958" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Osmola" birthdate="1991-02-21" gender="F" nation="POL" swrid="4124814" athleteid="3676">
              <RESULTS>
                <RESULT eventid="1247" points="373" swimtime="00:01:11.81" resultid="3677" heatid="3957" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="279" swimtime="00:06:01.56" resultid="3678" heatid="3976" lane="4" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:20.66" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                    <SPLIT distance="200" swimtime="00:02:48.86" />
                    <SPLIT distance="250" swimtime="00:03:35.53" />
                    <SPLIT distance="300" swimtime="00:04:23.75" />
                    <SPLIT distance="350" swimtime="00:05:12.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Wawrzyniak" birthdate="1986-11-27" gender="M" nation="POL" athleteid="3800">
              <RESULTS>
                <RESULT eventid="1199" points="202" swimtime="00:00:37.90" resultid="3801" heatid="3951" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1295" points="267" swimtime="00:01:12.77" resultid="3802" heatid="3959" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Zieliński" birthdate="1989-04-27" gender="M" nation="POL" swrid="4071551" athleteid="3671">
              <RESULTS>
                <RESULT eventid="1135" points="467" swimtime="00:00:33.43" resultid="3672" heatid="3942" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="3044" points="441" swimtime="00:01:14.70" resultid="3673" heatid="3965" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Konecki" birthdate="1982-02-22" gender="M" nation="POL" athleteid="3785">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="3786" heatid="3936" lane="1" entrytime="00:00:29.74" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="3787" heatid="3947" lane="7" entrytime="00:00:34.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Kuratczyk" birthdate="1979-06-27" gender="M" nation="POL" athleteid="3717">
              <RESULTS>
                <RESULT eventid="1103" points="394" swimtime="00:00:28.52" resultid="3718" heatid="3936" lane="0" entrytime="00:00:29.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Łopuszański" birthdate="1969-11-10" gender="M" nation="POL" athleteid="3685">
              <RESULTS>
                <RESULT eventid="1231" points="105" swimtime="00:04:01.57" resultid="3686" heatid="3955" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:57.03" />
                    <SPLIT distance="150" swimtime="00:03:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3108" points="94" swimtime="00:01:48.55" resultid="3687" heatid="3971" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Woźniak" birthdate="1986-08-22" gender="M" nation="POL" athleteid="3754">
              <RESULTS>
                <RESULT eventid="1103" points="141" swimtime="00:00:40.08" resultid="3755" heatid="3939" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Cylwik-Rokicka" birthdate="1970-05-12" gender="F" nation="POL" athleteid="3767">
              <RESULTS>
                <RESULT eventid="1151" points="117" swimtime="00:00:55.15" resultid="3768" heatid="3945" lane="9" />
                <RESULT eventid="1183" points="95" swimtime="00:00:53.47" resultid="3769" heatid="3949" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Szot" birthdate="1995-01-14" gender="M" nation="POL" swrid="4196783" athleteid="3776">
              <RESULTS>
                <RESULT eventid="1135" points="498" swimtime="00:00:32.73" resultid="3777" heatid="3942" lane="3" entrytime="00:00:32.55" />
                <RESULT eventid="3044" points="470" swimtime="00:01:13.15" resultid="3778" heatid="3965" lane="5" entrytime="00:01:11.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabella" lastname="Sylwestrzak" birthdate="1996-01-12" gender="F" nation="POL" swrid="4800790" athleteid="3746">
              <RESULTS>
                <RESULT eventid="1247" points="377" swimtime="00:01:11.57" resultid="3747" heatid="3957" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="297" swimtime="00:05:54.21" resultid="3748" heatid="3976" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:19.88" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                    <SPLIT distance="200" swimtime="00:02:50.99" />
                    <SPLIT distance="250" swimtime="00:03:37.50" />
                    <SPLIT distance="300" swimtime="00:04:24.09" />
                    <SPLIT distance="350" swimtime="00:05:09.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Hydrow" birthdate="1985-05-10" gender="M" nation="POL" athleteid="3797">
              <RESULTS>
                <RESULT eventid="1103" points="190" swimtime="00:00:36.32" resultid="3798" heatid="3940" lane="9" entrytime="00:00:29.00" />
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1199" status="DSQ" swimtime="00:00:00.00" resultid="3799" heatid="3951" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Kukla" birthdate="1990-12-20" gender="F" nation="POL" athleteid="3791">
              <RESULTS>
                <RESULT eventid="1058" points="91" swimtime="00:00:52.58" resultid="3792" heatid="3932" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1247" status="DNS" swimtime="00:00:00.00" resultid="3793" heatid="3957" lane="4" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Fijałkowski" birthdate="1972-01-27" gender="M" nation="POL" athleteid="3700">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="3701" heatid="3940" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kamut" birthdate="1977-12-29" gender="F" nation="POL" athleteid="3674">
              <RESULTS>
                <RESULT eventid="3160" points="118" swimtime="00:08:01.75" resultid="3675" heatid="3976" lane="8" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:47.28" />
                    <SPLIT distance="150" swimtime="00:02:50.19" />
                    <SPLIT distance="200" swimtime="00:03:52.77" />
                    <SPLIT distance="250" swimtime="00:04:56.64" />
                    <SPLIT distance="300" swimtime="00:06:00.28" />
                    <SPLIT distance="350" swimtime="00:07:03.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Szyszka" birthdate="1990-07-19" gender="M" nation="POL" athleteid="3782">
              <RESULTS>
                <RESULT eventid="1295" points="367" swimtime="00:01:05.50" resultid="3783" heatid="3960" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="350" swimtime="00:05:12.10" resultid="3784" heatid="3978" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:50.64" />
                    <SPLIT distance="200" swimtime="00:02:31.18" />
                    <SPLIT distance="250" swimtime="00:03:11.89" />
                    <SPLIT distance="300" swimtime="00:03:52.76" />
                    <SPLIT distance="350" swimtime="00:04:33.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Senger" birthdate="1982-03-27" gender="M" nation="POL" athleteid="3688">
              <RESULTS>
                <RESULT eventid="1295" points="192" swimtime="00:01:21.19" resultid="3689" heatid="3961" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="160" swimtime="00:06:45.08" resultid="3690" heatid="3979" lane="1" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:34.14" />
                    <SPLIT distance="150" swimtime="00:02:26.23" />
                    <SPLIT distance="200" swimtime="00:03:18.86" />
                    <SPLIT distance="250" swimtime="00:04:11.81" />
                    <SPLIT distance="300" swimtime="00:05:04.19" />
                    <SPLIT distance="350" swimtime="00:05:56.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Dębski" birthdate="1978-02-01" gender="M" nation="POL" athleteid="3803">
              <RESULTS>
                <RESULT eventid="1103" points="360" swimtime="00:00:29.37" resultid="3804" heatid="3937" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1199" points="284" swimtime="00:00:33.87" resultid="3805" heatid="3951" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamila" lastname="Patejko" birthdate="1984-05-17" gender="F" nation="POL" athleteid="3719">
              <RESULTS>
                <RESULT eventid="3092" points="120" swimtime="00:01:52.44" resultid="3720" heatid="3970" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="198" swimtime="00:06:45.40" resultid="3721" heatid="3976" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:36.94" />
                    <SPLIT distance="150" swimtime="00:02:27.87" />
                    <SPLIT distance="200" swimtime="00:03:19.27" />
                    <SPLIT distance="250" swimtime="00:04:10.98" />
                    <SPLIT distance="300" swimtime="00:05:03.35" />
                    <SPLIT distance="350" swimtime="00:05:55.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Petryszyn" birthdate="1994-07-31" gender="F" nation="POL" swrid="4369524" athleteid="3762">
              <RESULTS>
                <RESULT eventid="1058" points="508" swimtime="00:00:29.65" resultid="3763" heatid="3932" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1151" points="525" swimtime="00:00:33.43" resultid="3764" heatid="3945" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="3368" name="Warsaw Masters Team ">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Szymański" birthdate="1981-11-04" gender="M" nation="POL" license="504214700060" swrid="4542568" athleteid="3630">
              <RESULTS>
                <RESULT eventid="1103" points="375" swimtime="00:00:28.98" resultid="3631" heatid="3936" lane="4" entrytime="00:00:28.95" entrycourse="LCM" />
                <RESULT eventid="1199" points="329" swimtime="00:00:32.23" resultid="3632" heatid="3950" lane="8" entrytime="00:00:31.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Barcicka" birthdate="1993-09-28" gender="F" nation="POL" athleteid="3501">
              <RESULTS>
                <RESULT eventid="1058" points="249" swimtime="00:00:37.62" resultid="3502" heatid="3933" lane="3" entrytime="00:00:36.92" />
                <RESULT eventid="3160" points="177" swimtime="00:07:00.89" resultid="3503" heatid="3977" lane="4" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:35.34" />
                    <SPLIT distance="150" swimtime="00:02:26.57" />
                    <SPLIT distance="200" swimtime="00:03:19.20" />
                    <SPLIT distance="250" swimtime="00:04:12.83" />
                    <SPLIT distance="300" swimtime="00:05:08.41" />
                    <SPLIT distance="350" swimtime="00:06:05.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" athleteid="3396">
              <RESULTS>
                <RESULT eventid="1103" points="465" swimtime="00:00:26.98" resultid="3397" heatid="3935" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="1199" points="406" swimtime="00:00:30.07" resultid="3398" heatid="3950" lane="0" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Mostowska" birthdate="1977-06-20" gender="F" nation="POL" athleteid="3402">
              <RESULTS>
                <RESULT comment="GR 5.1, GR 5.2, GR 5.3" eventid="1215" status="DSQ" swimtime="00:00:00.00" resultid="3403" heatid="3954" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                    <SPLIT distance="100" swimtime="00:01:45.10" />
                    <SPLIT distance="150" swimtime="00:02:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="GR 5.1, GR 5.2, GR 5.3" eventid="3160" status="DSQ" swimtime="00:06:11.61" resultid="3404" heatid="3976" lane="7" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                    <SPLIT distance="150" swimtime="00:02:14.04" />
                    <SPLIT distance="200" swimtime="00:03:01.28" />
                    <SPLIT distance="250" swimtime="00:03:48.96" />
                    <SPLIT distance="300" swimtime="00:04:36.51" />
                    <SPLIT distance="350" swimtime="00:05:24.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Church" birthdate="1973-01-04" gender="F" nation="POL" athleteid="3414">
              <RESULTS>
                <RESULT eventid="1247" points="106" swimtime="00:01:49.02" resultid="3415" heatid="3957" lane="9" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3160" points="115" swimtime="00:08:06.08" resultid="3416" heatid="3977" lane="2" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:01:55.21" />
                    <SPLIT distance="150" swimtime="00:02:57.29" />
                    <SPLIT distance="200" swimtime="00:03:59.25" />
                    <SPLIT distance="250" swimtime="00:05:02.20" />
                    <SPLIT distance="300" swimtime="00:06:04.76" />
                    <SPLIT distance="350" swimtime="00:07:07.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Ostrzycki" birthdate="1949-04-10" gender="M" nation="POL" athleteid="3417">
              <RESULTS>
                <RESULT eventid="1135" points="157" swimtime="00:00:48.08" resultid="3418" heatid="3942" lane="0" entrytime="00:00:49.70" />
                <RESULT eventid="1295" status="DNS" swimtime="00:00:00.00" resultid="3419" heatid="3963" lane="4" entrytime="00:01:52.80" />
                <RESULT eventid="3044" points="141" swimtime="00:01:49.21" resultid="3975" heatid="3966" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Nowicki" birthdate="1963-02-18" gender="M" nation="POL" swrid="4754751" athleteid="3485">
              <RESULTS>
                <RESULT eventid="3182" points="93" swimtime="00:08:04.69" resultid="3486" heatid="3980" lane="4" entrytime="00:07:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.29" />
                    <SPLIT distance="100" swimtime="00:01:48.38" />
                    <SPLIT distance="150" swimtime="00:02:49.89" />
                    <SPLIT distance="200" swimtime="00:03:53.52" />
                    <SPLIT distance="250" swimtime="00:04:57.14" />
                    <SPLIT distance="300" swimtime="00:06:00.98" />
                    <SPLIT distance="350" swimtime="00:07:04.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kochanowski" birthdate="1981-11-11" gender="M" nation="POL" license="104214700135" athleteid="3633">
              <RESULTS>
                <RESULT eventid="1135" points="151" swimtime="00:00:48.71" resultid="3634" heatid="3943" lane="8" />
                <RESULT eventid="3044" points="146" swimtime="00:01:47.93" resultid="3635" heatid="3966" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlena" lastname="Dobrasiewicz" birthdate="1988-05-24" gender="F" nation="POL" athleteid="3488" />
            <ATHLETE firstname="Michał" lastname="Jabłoński" birthdate="1980-09-13" gender="M" nation="POL" swrid="5471784" athleteid="3446">
              <RESULTS>
                <RESULT eventid="1103" points="299" swimtime="00:00:31.25" resultid="3447" heatid="3936" lane="7" entrytime="00:00:29.70" />
                <RESULT eventid="1295" points="313" swimtime="00:01:09.05" resultid="3448" heatid="3959" lane="1" entrytime="00:01:07.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Guimard" birthdate="1970-01-09" gender="M" nation="POL" athleteid="3513">
              <RESULTS>
                <RESULT eventid="1103" points="199" swimtime="00:00:35.76" resultid="3514" heatid="3940" lane="6" />
                <RESULT eventid="1135" points="191" swimtime="00:00:45.04" resultid="3515" heatid="3943" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Wojciechowski" birthdate="1968-03-16" gender="M" nation="POL" athleteid="3369">
              <RESULTS>
                <RESULT eventid="1167" points="119" swimtime="00:00:48.79" resultid="3370" heatid="3947" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="3182" points="67" swimtime="00:08:59.50" resultid="3371" heatid="3980" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="100" swimtime="00:02:02.71" />
                    <SPLIT distance="150" swimtime="00:03:12.40" />
                    <SPLIT distance="200" swimtime="00:04:22.10" />
                    <SPLIT distance="250" swimtime="00:05:32.93" />
                    <SPLIT distance="300" swimtime="00:06:42.30" />
                    <SPLIT distance="350" swimtime="00:07:52.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kozysa" birthdate="1981-05-07" gender="M" nation="POL" athleteid="3435" />
            <ATHLETE firstname="Wojciech" lastname="Kałużyński" birthdate="1980-05-14" gender="M" nation="POL" swrid="4992656" athleteid="3479">
              <RESULTS>
                <RESULT comment="M4 - Pływak wykonał nierównoczesne ruchy ramion." eventid="1199" status="DSQ" swimtime="00:00:00.00" resultid="3480" heatid="3952" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1295" points="260" swimtime="00:01:13.42" resultid="3481" heatid="3960" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" athleteid="3381">
              <RESULTS>
                <RESULT eventid="1103" points="394" swimtime="00:00:28.51" resultid="3382" heatid="3935" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="1199" points="384" swimtime="00:00:30.63" resultid="3383" heatid="3950" lane="1" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Derezińska" birthdate="1974-03-27" gender="F" nation="POL" athleteid="3426">
              <RESULTS>
                <RESULT eventid="1119" points="211" swimtime="00:00:49.31" resultid="3427" heatid="3941" lane="8" entrytime="00:00:47.62" />
                <RESULT eventid="3160" points="161" swimtime="00:07:14.60" resultid="3428" heatid="3976" lane="0" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:42.87" />
                    <SPLIT distance="150" swimtime="00:02:36.85" />
                    <SPLIT distance="200" swimtime="00:03:32.71" />
                    <SPLIT distance="250" swimtime="00:04:27.50" />
                    <SPLIT distance="300" swimtime="00:05:24.45" />
                    <SPLIT distance="350" swimtime="00:06:19.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Wierciński" birthdate="1988-04-04" gender="M" nation="POL" athleteid="3516">
              <RESULTS>
                <RESULT eventid="1295" points="177" swimtime="00:01:23.44" resultid="3517" heatid="3961" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3044" points="165" swimtime="00:01:43.62" resultid="3518" heatid="3965" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Galica" birthdate="1985-11-26" gender="F" nation="POL" athleteid="3455">
              <RESULTS>
                <RESULT eventid="1183" points="303" swimtime="00:00:36.35" resultid="3456" heatid="3949" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="3160" points="316" swimtime="00:05:47.15" resultid="3457" heatid="3976" lane="3" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="150" swimtime="00:02:00.07" />
                    <SPLIT distance="200" swimtime="00:02:45.03" />
                    <SPLIT distance="250" swimtime="00:03:31.14" />
                    <SPLIT distance="300" swimtime="00:04:17.53" />
                    <SPLIT distance="350" swimtime="00:05:04.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Chrostowski" birthdate="1989-01-11" gender="M" nation="POL" swrid="5471781" athleteid="3443">
              <RESULTS>
                <RESULT eventid="1103" points="228" swimtime="00:00:34.19" resultid="3444" heatid="3939" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1295" points="191" swimtime="00:01:21.35" resultid="3445" heatid="3961" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Giejsztowt" birthdate="1978-06-13" gender="M" nation="POL" swrid="5241012" athleteid="3423">
              <RESULTS>
                <RESULT eventid="1295" points="431" swimtime="00:01:02.06" resultid="3424" heatid="3959" lane="6" entrytime="00:01:02.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="376" swimtime="00:05:04.66" resultid="3425" heatid="3978" lane="3" entrytime="00:05:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:51.60" />
                    <SPLIT distance="200" swimtime="00:02:31.55" />
                    <SPLIT distance="250" swimtime="00:03:09.64" />
                    <SPLIT distance="300" swimtime="00:03:47.21" />
                    <SPLIT distance="350" swimtime="00:04:26.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Prasał" birthdate="1977-05-29" gender="M" nation="POL" athleteid="3438">
              <RESULTS>
                <RESULT eventid="1103" points="236" swimtime="00:00:33.83" resultid="3439" heatid="3938" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Suchecka" birthdate="1999-09-09" gender="F" nation="POL" swrid="4493009" athleteid="3504">
              <RESULTS>
                <RESULT eventid="1058" points="443" swimtime="00:00:31.03" resultid="3505" heatid="3932" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1151" points="510" swimtime="00:00:33.75" resultid="3506" heatid="3945" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Sutowski" birthdate="1959-12-03" gender="M" nation="POL" license="104214700079" swrid="4992657" athleteid="3639">
              <RESULTS>
                <RESULT eventid="1295" points="144" swimtime="00:01:29.31" resultid="3640" heatid="3962" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="158" swimtime="00:06:46.91" resultid="3641" heatid="3980" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                    <SPLIT distance="100" swimtime="00:01:36.54" />
                    <SPLIT distance="150" swimtime="00:02:29.06" />
                    <SPLIT distance="200" swimtime="00:03:22.34" />
                    <SPLIT distance="250" swimtime="00:04:16.52" />
                    <SPLIT distance="300" swimtime="00:05:08.13" />
                    <SPLIT distance="350" swimtime="00:05:59.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Sołtan" birthdate="1975-12-02" gender="M" nation="POL" swrid="4384324" athleteid="3393">
              <RESULTS>
                <RESULT eventid="1231" points="365" swimtime="00:02:39.47" resultid="3394" heatid="3955" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:02:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="396" swimtime="00:04:59.61" resultid="3395" heatid="3978" lane="2" entrytime="00:05:12.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:51.98" />
                    <SPLIT distance="200" swimtime="00:02:31.00" />
                    <SPLIT distance="250" swimtime="00:03:08.42" />
                    <SPLIT distance="300" swimtime="00:03:45.49" />
                    <SPLIT distance="350" swimtime="00:04:22.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Dargas-Miszczak" birthdate="1981-09-06" gender="F" nation="POL" swrid="5486407" athleteid="3411">
              <RESULTS>
                <RESULT eventid="1058" points="285" swimtime="00:00:35.96" resultid="3412" heatid="3933" lane="5" entrytime="00:00:36.25" />
                <RESULT eventid="1215" points="238" swimtime="00:03:23.28" resultid="3413" heatid="3954" lane="2" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:40.48" />
                    <SPLIT distance="150" swimtime="00:02:35.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Saienko" birthdate="1994-08-03" gender="M" nation="UKR" athleteid="3399">
              <RESULTS>
                <RESULT eventid="1103" points="521" swimtime="00:00:25.98" resultid="3400" heatid="3935" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1199" points="489" swimtime="00:00:28.26" resultid="3401" heatid="3950" lane="3" entrytime="00:00:27.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magda" lastname="Mazurkiewicz" birthdate="1976-03-14" gender="F" nation="POL" athleteid="3507">
              <RESULTS>
                <RESULT eventid="1151" points="193" swimtime="00:00:46.62" resultid="3508" heatid="3946" lane="5" />
                <RESULT eventid="3160" points="164" swimtime="00:07:11.30" resultid="3509" heatid="3977" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:36.11" />
                    <SPLIT distance="150" swimtime="00:02:30.79" />
                    <SPLIT distance="200" swimtime="00:03:26.26" />
                    <SPLIT distance="250" swimtime="00:04:23.91" />
                    <SPLIT distance="300" swimtime="00:05:20.18" />
                    <SPLIT distance="350" swimtime="00:06:16.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Kuc" birthdate="1976-03-16" gender="F" nation="POL" license="504214600040" athleteid="3627">
              <RESULTS>
                <RESULT eventid="1058" points="145" swimtime="00:00:44.96" resultid="3628" heatid="3934" lane="6" />
                <RESULT eventid="1247" points="139" swimtime="00:01:39.75" resultid="3629" heatid="3958" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zenon" lastname="Kuliś" birthdate="1954-06-04" gender="M" nation="POL" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1167" points="95" swimtime="00:00:52.42" resultid="3433" heatid="3947" lane="9" entrytime="00:00:54.50" />
                <RESULT eventid="1295" points="118" swimtime="00:01:35.57" resultid="3434" heatid="3961" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Budek" birthdate="1974-10-20" gender="M" nation="POL" swrid="4992736" athleteid="3482">
              <RESULTS>
                <RESULT eventid="1103" points="254" swimtime="00:00:33.00" resultid="3483" heatid="3939" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1295" points="207" swimtime="00:01:19.27" resultid="3484" heatid="3961" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Wnuk" birthdate="1968-04-25" gender="F" nation="POL" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1058" points="119" swimtime="00:00:48.05" resultid="3406" heatid="3933" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1215" points="89" swimtime="00:04:42.45" resultid="3407" heatid="3954" lane="0" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.24" />
                    <SPLIT distance="100" swimtime="00:02:20.27" />
                    <SPLIT distance="150" swimtime="00:03:35.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" athleteid="3378">
              <RESULTS>
                <RESULT eventid="3044" points="293" swimtime="00:01:25.57" resultid="3379" heatid="3965" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="224" swimtime="00:06:02.05" resultid="3380" heatid="3979" lane="3" entrytime="00:06:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="150" swimtime="00:02:09.14" />
                    <SPLIT distance="200" swimtime="00:02:55.72" />
                    <SPLIT distance="250" swimtime="00:03:43.18" />
                    <SPLIT distance="300" swimtime="00:04:30.74" />
                    <SPLIT distance="350" swimtime="00:05:18.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" swrid="4183802" athleteid="3489">
              <RESULTS>
                <RESULT eventid="1231" points="381" swimtime="00:02:37.18" resultid="3490" heatid="3955" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:02:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3076" points="366" swimtime="00:01:12.44" resultid="3491" heatid="3968" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Olszewski" birthdate="1989-07-28" gender="M" nation="POL" swrid="4112408" athleteid="3449">
              <RESULTS>
                <RESULT eventid="1167" points="419" swimtime="00:00:32.06" resultid="3450" heatid="3947" lane="3" entrytime="00:00:32.41" />
                <RESULT eventid="3076" points="363" swimtime="00:01:12.65" resultid="3451" heatid="3968" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Białorucki" birthdate="1983-08-17" gender="M" nation="POL" athleteid="3519">
              <RESULTS>
                <RESULT eventid="1103" points="301" swimtime="00:00:31.20" resultid="3520" heatid="3938" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="1199" points="215" swimtime="00:00:37.14" resultid="3521" heatid="3951" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Sutowski" birthdate="1993-02-18" gender="M" nation="POL" swrid="4073514" athleteid="3372">
              <RESULTS>
                <RESULT eventid="1103" points="350" swimtime="00:00:29.67" resultid="3373" heatid="3936" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1295" points="312" swimtime="00:01:09.16" resultid="3374" heatid="3959" lane="0" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Maliszewski" birthdate="1974-03-01" gender="M" nation="POL" license="504214700126" athleteid="3642">
              <RESULTS>
                <RESULT eventid="1295" points="213" swimtime="00:01:18.43" resultid="3643" heatid="3962" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="172" swimtime="00:06:35.11" resultid="3644" heatid="3980" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:22.64" />
                    <SPLIT distance="200" swimtime="00:03:13.81" />
                    <SPLIT distance="250" swimtime="00:04:05.67" />
                    <SPLIT distance="300" swimtime="00:04:57.37" />
                    <SPLIT distance="350" swimtime="00:05:47.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Warakomski" birthdate="1981-04-17" gender="M" nation="POL" athleteid="3495">
              <RESULTS>
                <RESULT eventid="1103" points="271" swimtime="00:00:32.28" resultid="3496" heatid="3938" lane="4" entrytime="00:00:32.20" />
                <RESULT eventid="3108" points="182" swimtime="00:01:27.21" resultid="3497" heatid="3971" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szymański" birthdate="1980-10-04" gender="M" nation="POL" swrid="4542528" athleteid="3461">
              <RESULTS>
                <RESULT eventid="1103" points="522" swimtime="00:00:25.96" resultid="3462" heatid="3935" lane="6" entrytime="00:00:25.50" />
                <RESULT eventid="1167" points="514" swimtime="00:00:29.96" resultid="3463" heatid="3947" lane="4" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Pfitzner" birthdate="1986-05-24" gender="M" nation="POL" swrid="4992671" athleteid="3429">
              <RESULTS>
                <RESULT eventid="1199" points="436" swimtime="00:00:29.36" resultid="3430" heatid="3950" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="3182" points="383" swimtime="00:05:02.99" resultid="3431" heatid="3978" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:28.48" />
                    <SPLIT distance="250" swimtime="00:03:06.62" />
                    <SPLIT distance="300" swimtime="00:03:45.84" />
                    <SPLIT distance="350" swimtime="00:04:25.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Tomaszewski" birthdate="1950-06-24" gender="M" nation="POL" athleteid="3420">
              <RESULTS>
                <RESULT eventid="1103" points="42" swimtime="00:00:59.69" resultid="3421" heatid="3940" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="1167" points="43" swimtime="00:01:08.14" resultid="3422" heatid="3948" lane="4" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Kowalska" birthdate="1989-09-09" gender="F" nation="POL" athleteid="3492">
              <RESULTS>
                <RESULT eventid="1058" points="270" swimtime="00:00:36.61" resultid="3493" heatid="3933" lane="1" entrytime="00:00:38.20" />
                <RESULT eventid="3160" points="204" swimtime="00:06:41.14" resultid="3494" heatid="3976" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:33.24" />
                    <SPLIT distance="150" swimtime="00:02:23.61" />
                    <SPLIT distance="200" swimtime="00:03:14.79" />
                    <SPLIT distance="250" swimtime="00:04:06.68" />
                    <SPLIT distance="300" swimtime="00:04:58.46" />
                    <SPLIT distance="350" swimtime="00:05:51.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Grochowski" birthdate="1991-08-29" gender="M" nation="POL" swrid="5464090" athleteid="3390">
              <RESULTS>
                <RESULT eventid="1199" points="252" swimtime="00:00:35.25" resultid="3391" heatid="3951" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="3182" points="301" swimtime="00:05:28.26" resultid="3392" heatid="3978" lane="7" entrytime="00:05:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                    <SPLIT distance="200" swimtime="00:02:32.97" />
                    <SPLIT distance="250" swimtime="00:03:15.06" />
                    <SPLIT distance="300" swimtime="00:03:57.75" />
                    <SPLIT distance="350" swimtime="00:04:42.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Nowak" birthdate="1952-12-17" gender="M" nation="POL" swrid="4302652" athleteid="3467">
              <RESULTS>
                <RESULT eventid="1135" points="287" swimtime="00:00:39.34" resultid="3468" heatid="3942" lane="7" entrytime="00:00:37.90" />
                <RESULT eventid="3044" points="216" swimtime="00:01:34.71" resultid="3469" heatid="3965" lane="2" entrytime="00:01:38.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Szymańska" birthdate="1985-05-31" gender="F" nation="POL" swrid="5312493" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1058" points="244" swimtime="00:00:37.87" resultid="3465" heatid="3933" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1247" points="212" swimtime="00:01:26.67" resultid="3466" heatid="3957" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Mazurkiewicz" birthdate="1974-05-09" gender="M" nation="POL" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1231" points="128" swimtime="00:03:45.78" resultid="3376" heatid="3955" lane="1" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:53.80" />
                    <SPLIT distance="150" swimtime="00:02:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="163" swimtime="00:06:42.15" resultid="3377" heatid="3979" lane="2" entrytime="00:06:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:19.30" />
                    <SPLIT distance="200" swimtime="00:03:11.24" />
                    <SPLIT distance="250" swimtime="00:04:04.60" />
                    <SPLIT distance="300" swimtime="00:04:57.82" />
                    <SPLIT distance="350" swimtime="00:05:51.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Burdelak" birthdate="1991-07-06" gender="F" nation="POL" swrid="4072596" athleteid="3387">
              <RESULTS>
                <RESULT eventid="1058" points="521" swimtime="00:00:29.40" resultid="3388" heatid="3932" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1119" points="496" swimtime="00:00:37.14" resultid="3389" heatid="3941" lane="4" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kielczyk" birthdate="1974-10-22" gender="F" nation="POL" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1058" points="402" swimtime="00:00:32.05" resultid="3441" heatid="3932" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1151" points="404" swimtime="00:00:36.48" resultid="3442" heatid="3945" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Czupryn" birthdate="1958-06-02" gender="M" nation="POL" swrid="4992673" athleteid="3510">
              <RESULTS>
                <RESULT eventid="1295" points="145" swimtime="00:01:29.19" resultid="3511" heatid="3961" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="130" swimtime="00:07:13.39" resultid="3512" heatid="3979" lane="7" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:39.52" />
                    <SPLIT distance="150" swimtime="00:02:35.51" />
                    <SPLIT distance="200" swimtime="00:03:31.28" />
                    <SPLIT distance="250" swimtime="00:04:26.95" />
                    <SPLIT distance="300" swimtime="00:05:23.04" />
                    <SPLIT distance="350" swimtime="00:06:19.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Mukułowski" birthdate="1987-05-18" gender="M" nation="POL" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1103" points="294" swimtime="00:00:31.42" resultid="3471" heatid="3938" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1295" points="275" swimtime="00:01:12.09" resultid="3472" heatid="3960" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Skorykow" birthdate="1969-04-17" gender="M" nation="POL" athleteid="3487" />
            <ATHLETE firstname="Monika" lastname="Jarecka-Skorykow" birthdate="1974-01-30" gender="F" nation="POL" swrid="4992672" athleteid="3408">
              <RESULTS>
                <RESULT eventid="1058" points="384" swimtime="00:00:32.54" resultid="3810" heatid="3932" lane="0" entrytime="00:00:34.90" />
                <RESULT eventid="1119" points="314" swimtime="00:00:43.22" resultid="3811" heatid="3941" lane="1" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Rąpała" birthdate="1962-12-05" gender="M" nation="POL" athleteid="3473">
              <RESULTS>
                <RESULT eventid="1103" points="155" swimtime="00:00:38.92" resultid="3474" heatid="3938" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1199" points="79" swimtime="00:00:51.79" resultid="3475" heatid="3952" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Kubiszewski- Jakubiak" birthdate="1979-02-18" gender="M" nation="POL" athleteid="3458">
              <RESULTS>
                <RESULT eventid="1103" points="298" swimtime="00:00:31.29" resultid="3459" heatid="3937" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1135" points="253" swimtime="00:00:40.99" resultid="3460" heatid="3942" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" swrid="4302692" athleteid="3384">
              <RESULTS>
                <RESULT eventid="1058" points="71" swimtime="00:00:56.93" resultid="3385" heatid="3934" lane="4" entrytime="00:00:59.07" />
                <RESULT eventid="3160" points="73" swimtime="00:09:25.48" resultid="3386" heatid="3977" lane="1" entrytime="00:09:38.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.47" />
                    <SPLIT distance="100" swimtime="00:02:16.62" />
                    <SPLIT distance="150" swimtime="00:03:29.37" />
                    <SPLIT distance="200" swimtime="00:04:41.42" />
                    <SPLIT distance="250" swimtime="00:05:53.37" />
                    <SPLIT distance="300" swimtime="00:07:05.14" />
                    <SPLIT distance="350" swimtime="00:08:16.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Paluszak" birthdate="1967-02-17" gender="M" nation="POL" license="504214700102" swrid="5471792" athleteid="3636">
              <RESULTS>
                <RESULT eventid="1199" points="127" swimtime="00:00:44.25" resultid="3637" heatid="3952" lane="4" entrytime="00:00:43.35" entrycourse="LCM" />
                <RESULT eventid="3108" points="99" swimtime="00:01:46.91" resultid="3638" heatid="3971" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" swrid="4222718" athleteid="3476">
              <RESULTS>
                <RESULT eventid="1103" points="298" swimtime="00:00:31.29" resultid="3477" heatid="3936" lane="2" entrytime="00:00:29.65" />
                <RESULT eventid="3182" points="259" swimtime="00:05:44.85" resultid="3478" heatid="3979" lane="4" entrytime="00:05:46.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:03.73" />
                    <SPLIT distance="200" swimtime="00:02:48.14" />
                    <SPLIT distance="250" swimtime="00:03:32.60" />
                    <SPLIT distance="300" swimtime="00:04:17.57" />
                    <SPLIT distance="350" swimtime="00:05:02.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Worsztynowicz" birthdate="1987-06-14" gender="F" nation="POL" athleteid="3436">
              <RESULTS>
                <RESULT eventid="1151" points="207" swimtime="00:00:45.57" resultid="3437" heatid="3945" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 1" number="1">
              <RESULTS>
                <RESULT eventid="3124" points="491" swimtime="00:02:05.25" resultid="3525" heatid="3972" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="150" swimtime="00:01:33.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3461" number="1" />
                    <RELAYPOSITION athleteid="3387" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3399" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3440" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 2" number="2">
              <RESULTS>
                <RESULT eventid="3124" points="288" swimtime="00:02:29.58" resultid="3523" heatid="3972" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3390" number="1" />
                    <RELAYPOSITION athleteid="3464" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3381" number="3" />
                    <RELAYPOSITION athleteid="3455" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 4" number="4">
              <RESULTS>
                <RESULT eventid="3124" points="217" swimtime="00:02:44.34" resultid="3524" heatid="3972" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="100" swimtime="00:01:31.10" />
                    <SPLIT distance="150" swimtime="00:02:12.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3436" number="1" />
                    <RELAYPOSITION athleteid="3438" number="2" />
                    <RELAYPOSITION athleteid="3411" number="3" />
                    <RELAYPOSITION athleteid="3435" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 5" number="5">
              <RESULTS>
                <RESULT eventid="3124" points="170" swimtime="00:02:58.18" resultid="3526" heatid="3972" lane="2" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.36" />
                    <SPLIT distance="100" swimtime="00:01:42.90" />
                    <SPLIT distance="150" swimtime="00:01:20.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3375" number="1" />
                    <RELAYPOSITION athleteid="3426" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3495" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="3492" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 6" number="6">
              <RESULTS>
                <RESULT comment="K10 - Pływak przeniósł dłonie poza linię bioder (z wyjątkiem pierwszego ruchu ramion po starcie i nawrotach)." eventid="3124" status="DSQ" swimtime="00:03:03.26" resultid="3528" heatid="3972" lane="0" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:43.55" />
                    <SPLIT distance="150" swimtime="00:02:26.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3369" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3507" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3443" number="3" reactiontime="+60" status="DSQ" />
                    <RELAYPOSITION athleteid="3501" number="4" reactiontime="+37" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="WMT 7" number="7">
              <RESULTS>
                <RESULT eventid="3124" points="364" swimtime="00:02:18.28" resultid="3527" heatid="3972" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:47.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3487" number="1" />
                    <RELAYPOSITION athleteid="3408" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3396" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3488" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NEOSTR" nation="POL" clubid="3806" name="UKS NEPTUN Ostrów Mazowiecka">
          <ATHLETES>
            <ATHLETE firstname="Ewelina" lastname="Budek" birthdate="1979-01-16" gender="F" nation="POL" athleteid="3807">
              <RESULTS>
                <RESULT eventid="1058" points="168" swimtime="00:00:42.86" resultid="3808" heatid="3933" lane="7" entrytime="00:00:38.07" entrycourse="LCM" />
                <RESULT eventid="1119" points="182" swimtime="00:00:51.84" resultid="3809" heatid="3941" lane="6" entrytime="00:00:41.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3328" name="Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Boboli" birthdate="1948-01-01" gender="M" nation="POL" athleteid="3329">
              <RESULTS>
                <RESULT eventid="1103" points="149" swimtime="00:00:39.43" resultid="3330" heatid="3939" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1199" points="70" swimtime="00:00:53.95" resultid="3331" heatid="3951" lane="9" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3205" name="Masters Zdzieszowice">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" swrid="4992846" athleteid="3206">
              <RESULTS>
                <RESULT eventid="1215" points="267" swimtime="00:03:15.83" resultid="3207" heatid="3954" lane="3" entrytime="00:02:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="150" swimtime="00:02:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3092" points="259" swimtime="00:01:27.03" resultid="3208" heatid="3970" lane="4" entrytime="00:01:27.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" clubid="3226" name="Korona Kraków Masters">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Kaczmarczyk" birthdate="1968-01-02" gender="M" nation="POL" swrid="4992805" athleteid="3230">
              <RESULTS>
                <RESULT eventid="1103" points="77" swimtime="00:00:49.15" resultid="3231" heatid="3940" lane="0" />
                <RESULT eventid="1135" points="118" swimtime="00:00:52.86" resultid="3232" heatid="3944" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="3588" name="Towarzystwo Pływackie ,,Masters&apos;&apos; Opole">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" license="100607700003" swrid="4843497" athleteid="3589">
              <RESULTS>
                <RESULT eventid="1167" points="410" swimtime="00:00:32.28" resultid="3590" heatid="3947" lane="6" entrytime="00:00:32.47" entrycourse="LCM" />
                <RESULT eventid="3076" points="390" swimtime="00:01:10.92" resultid="3591" heatid="3968" lane="3" entrytime="00:01:10.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEOST" nation="POL" region="14" clubid="3974" name="Niezrzeszony Ostrołeka UŚKS">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Ambroziak" birthdate="1964-03-09" gender="M" nation="POL" athleteid="3773">
              <RESULTS>
                <RESULT eventid="1103" points="234" swimtime="00:00:33.90" resultid="3774" heatid="3938" lane="3" entrytime="00:00:33.30" />
                <RESULT eventid="3182" points="140" swimtime="00:07:03.81" resultid="3775" heatid="3979" lane="8" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:35.60" />
                    <SPLIT distance="100" swimtime="00:03:31.34" />
                    <SPLIT distance="150" swimtime="00:04:25.89" />
                    <SPLIT distance="200" swimtime="00:05:20.41" />
                    <SPLIT distance="300" swimtime="00:07:03.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" clubid="3198" name="Landsberg Crew Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Kaczmarek" birthdate="1992-08-23" gender="F" nation="POL" license="501304600002" athleteid="3199">
              <RESULTS>
                <RESULT eventid="1215" points="524" swimtime="00:02:36.41" resultid="3200" heatid="3954" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:59.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="507" swimtime="00:01:04.82" resultid="3201" heatid="3957" lane="5" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" license="501304700001" swrid="4432188" athleteid="3202">
              <RESULTS>
                <RESULT eventid="1231" points="470" swimtime="00:02:26.58" resultid="3203" heatid="3955" lane="4" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="150" swimtime="00:01:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3182" points="464" swimtime="00:04:44.16" resultid="3204" heatid="3978" lane="4" entrytime="00:04:28.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:47.01" />
                    <SPLIT distance="200" swimtime="00:02:23.97" />
                    <SPLIT distance="250" swimtime="00:03:00.37" />
                    <SPLIT distance="300" swimtime="00:03:36.42" />
                    <SPLIT distance="350" swimtime="00:04:11.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="3559" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="3560">
              <RESULTS>
                <RESULT eventid="1167" points="98" swimtime="00:00:51.89" resultid="3561" heatid="3947" lane="0" entrytime="00:00:53.36" entrycourse="SCM" />
                <RESULT eventid="3076" points="91" swimtime="00:01:55.01" resultid="3562" heatid="3968" lane="8" entrytime="00:01:55.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="MKS ZNICZ Koszalin" version="11.54147">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="Letnie Otwarte Mistrzostwa Polski w Pływaniu w Kategoriach MASTERS POZNAŃ 2018 PUCHAR MASTERS 2018" course="LCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2018-06-24" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Poznań" nation="POL" />
      <POINTTABLE pointtableid="3011" name="FINA Point Scoring" version="2018" />
      <SESSIONS>
        <SESSION date="2018-06-22" daytime="14:00" endtime="20:49" number="1">
          <EVENTS>
            <EVENT eventid="1229" daytime="14:52" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9655" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8887" />
                    <RANKING order="2" place="2" resultid="7702" />
                    <RANKING order="3" place="3" resultid="8858" />
                    <RANKING order="4" place="4" resultid="5751" />
                    <RANKING order="5" place="5" resultid="5675" />
                    <RANKING order="6" place="6" resultid="8311" />
                    <RANKING order="7" place="7" resultid="5735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9656" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7563" />
                    <RANKING order="2" place="2" resultid="5855" />
                    <RANKING order="3" place="3" resultid="6709" />
                    <RANKING order="4" place="4" resultid="8959" />
                    <RANKING order="5" place="5" resultid="8714" />
                    <RANKING order="6" place="6" resultid="7316" />
                    <RANKING order="7" place="-1" resultid="7103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9657" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7923" />
                    <RANKING order="2" place="2" resultid="7198" />
                    <RANKING order="3" place="3" resultid="8361" />
                    <RANKING order="4" place="4" resultid="8799" />
                    <RANKING order="5" place="-1" resultid="8339" />
                    <RANKING order="6" place="-1" resultid="8329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9658" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8849" />
                    <RANKING order="2" place="2" resultid="6244" />
                    <RANKING order="3" place="3" resultid="7362" />
                    <RANKING order="4" place="4" resultid="7298" />
                    <RANKING order="5" place="5" resultid="6679" />
                    <RANKING order="6" place="6" resultid="5969" />
                    <RANKING order="7" place="-1" resultid="7468" />
                    <RANKING order="8" place="-1" resultid="8366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9659" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8773" />
                    <RANKING order="2" place="2" resultid="8924" />
                    <RANKING order="3" place="3" resultid="7423" />
                    <RANKING order="4" place="4" resultid="7412" />
                    <RANKING order="5" place="5" resultid="7759" />
                    <RANKING order="6" place="6" resultid="7747" />
                    <RANKING order="7" place="7" resultid="7814" />
                    <RANKING order="8" place="8" resultid="8575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9660" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6534" />
                    <RANKING order="2" place="2" resultid="7694" />
                    <RANKING order="3" place="3" resultid="5744" />
                    <RANKING order="4" place="4" resultid="6556" />
                    <RANKING order="5" place="5" resultid="6427" />
                    <RANKING order="6" place="6" resultid="6370" />
                    <RANKING order="7" place="7" resultid="7239" />
                    <RANKING order="8" place="8" resultid="8275" />
                    <RANKING order="9" place="9" resultid="8781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9661" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6061" />
                    <RANKING order="2" place="2" resultid="7492" />
                    <RANKING order="3" place="3" resultid="7503" />
                    <RANKING order="4" place="4" resultid="5986" />
                    <RANKING order="5" place="5" resultid="7667" />
                    <RANKING order="6" place="-1" resultid="6646" />
                    <RANKING order="7" place="-1" resultid="7381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9662" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6085" />
                    <RANKING order="2" place="2" resultid="6120" />
                    <RANKING order="3" place="3" resultid="6608" />
                    <RANKING order="4" place="-1" resultid="6821" />
                    <RANKING order="5" place="-1" resultid="8297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9663" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6212" />
                    <RANKING order="2" place="2" resultid="7178" />
                    <RANKING order="3" place="3" resultid="6736" />
                    <RANKING order="4" place="4" resultid="8260" />
                    <RANKING order="5" place="5" resultid="7053" />
                    <RANKING order="6" place="6" resultid="8963" />
                    <RANKING order="7" place="7" resultid="6204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9664" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7738" />
                    <RANKING order="2" place="2" resultid="7349" />
                    <RANKING order="3" place="3" resultid="6809" />
                    <RANKING order="4" place="4" resultid="5795" />
                    <RANKING order="5" place="5" resultid="8613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9665" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6075" />
                    <RANKING order="2" place="2" resultid="6409" />
                    <RANKING order="3" place="3" resultid="5682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9666" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7150" />
                    <RANKING order="2" place="2" resultid="5779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9667" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9668" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9669" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9670" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9342" daytime="14:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9343" daytime="14:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9344" daytime="15:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9345" daytime="15:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9346" daytime="15:12" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9347" daytime="15:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9348" daytime="15:18" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9349" daytime="15:22" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1133" daytime="14:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6570" />
                    <RANKING order="2" place="2" resultid="6561" />
                    <RANKING order="3" place="3" resultid="8969" />
                    <RANKING order="4" place="4" resultid="6718" />
                    <RANKING order="5" place="5" resultid="8989" />
                    <RANKING order="6" place="6" resultid="8304" />
                    <RANKING order="7" place="7" resultid="8805" />
                    <RANKING order="8" place="8" resultid="7573" />
                    <RANKING order="9" place="9" resultid="7553" />
                    <RANKING order="10" place="10" resultid="9307" />
                    <RANKING order="11" place="-1" resultid="5824" />
                    <RANKING order="12" place="-1" resultid="7113" />
                    <RANKING order="13" place="-1" resultid="7649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7916" />
                    <RANKING order="2" place="2" resultid="7579" />
                    <RANKING order="3" place="3" resultid="6252" />
                    <RANKING order="4" place="4" resultid="5924" />
                    <RANKING order="5" place="5" resultid="7061" />
                    <RANKING order="6" place="6" resultid="8535" />
                    <RANKING order="7" place="7" resultid="7557" />
                    <RANKING order="8" place="8" resultid="6158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6352" />
                    <RANKING order="2" place="2" resultid="8678" />
                    <RANKING order="3" place="3" resultid="5849" />
                    <RANKING order="4" place="4" resultid="7304" />
                    <RANKING order="5" place="5" resultid="7187" />
                    <RANKING order="6" place="6" resultid="7935" />
                    <RANKING order="7" place="7" resultid="6024" />
                    <RANKING order="8" place="8" resultid="6760" />
                    <RANKING order="9" place="9" resultid="6640" />
                    <RANKING order="10" place="10" resultid="6749" />
                    <RANKING order="11" place="-1" resultid="8374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6577" />
                    <RANKING order="2" place="2" resultid="7968" />
                    <RANKING order="3" place="3" resultid="8766" />
                    <RANKING order="4" place="4" resultid="7485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7227" />
                    <RANKING order="2" place="2" resultid="7271" />
                    <RANKING order="3" place="3" resultid="7807" />
                    <RANKING order="4" place="4" resultid="7841" />
                    <RANKING order="5" place="5" resultid="8786" />
                    <RANKING order="6" place="6" resultid="7570" />
                    <RANKING order="7" place="7" resultid="8982" />
                    <RANKING order="8" place="8" resultid="8837" />
                    <RANKING order="9" place="-1" resultid="7639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6435" />
                    <RANKING order="2" place="2" resultid="7209" />
                    <RANKING order="3" place="3" resultid="6491" />
                    <RANKING order="4" place="4" resultid="6017" />
                    <RANKING order="5" place="-1" resultid="5919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6419" />
                    <RANKING order="2" place="2" resultid="6730" />
                    <RANKING order="3" place="3" resultid="8722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6270" />
                    <RANKING order="2" place="2" resultid="6219" />
                    <RANKING order="3" place="3" resultid="6448" />
                    <RANKING order="4" place="4" resultid="7627" />
                    <RANKING order="5" place="5" resultid="6315" />
                    <RANKING order="6" place="6" resultid="5951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8832" />
                    <RANKING order="2" place="2" resultid="6500" />
                    <RANKING order="3" place="3" resultid="5960" />
                    <RANKING order="4" place="4" resultid="5910" />
                    <RANKING order="5" place="5" resultid="8672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8283" />
                    <RANKING order="2" place="2" resultid="6901" />
                    <RANKING order="3" place="3" resultid="7158" />
                    <RANKING order="4" place="4" resultid="8880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6889" />
                    <RANKING order="2" place="2" resultid="6466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="1175" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="1194" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="1176" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9308" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9309" daytime="14:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9310" daytime="14:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9311" daytime="14:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9312" daytime="14:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9313" daytime="14:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9314" daytime="14:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9315" daytime="14:10" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1297" daytime="17:36" gender="F" number="8" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9703" agemax="24" agemin="20" name="Kat. 0" />
                <AGEGROUP agegroupid="9704" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="9705" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="9706" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="9707" agemax="44" agemin="40" name="Kat. D" />
                <AGEGROUP agegroupid="9708" agemax="49" agemin="45" name="Kat. E" />
                <AGEGROUP agegroupid="9709" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9710" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6336" />
                    <RANKING order="2" place="2" resultid="7847" />
                    <RANKING order="3" place="3" resultid="5952" />
                    <RANKING order="4" place="4" resultid="6633" />
                    <RANKING order="5" place="5" resultid="9436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9711" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="9712" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8284" />
                    <RANKING order="2" place="2" resultid="7397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9713" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="9714" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9715" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9716" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9717" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9718" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9364" daytime="17:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1263" daytime="15:32" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9671" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9672" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7057" />
                    <RANKING order="2" place="2" resultid="8976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9673" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7408" />
                    <RANKING order="2" place="2" resultid="9034" />
                    <RANKING order="3" place="-1" resultid="6641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9674" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6311" />
                    <RANKING order="2" place="2" resultid="8565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9675" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6169" />
                    <RANKING order="2" place="2" resultid="7219" />
                    <RANKING order="3" place="3" resultid="7616" />
                    <RANKING order="4" place="4" resultid="6383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9676" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6926" />
                    <RANKING order="2" place="2" resultid="7210" />
                    <RANKING order="3" place="3" resultid="7292" />
                    <RANKING order="4" place="4" resultid="8666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9677" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6844" />
                    <RANKING order="2" place="2" resultid="8861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9678" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6449" />
                    <RANKING order="2" place="2" resultid="6476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9679" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6501" />
                    <RANKING order="2" place="2" resultid="5883" />
                    <RANKING order="3" place="3" resultid="5911" />
                    <RANKING order="4" place="4" resultid="8909" />
                    <RANKING order="5" place="-1" resultid="5961" />
                    <RANKING order="6" place="-1" resultid="7074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9680" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9681" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="9682" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9683" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9684" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9685" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9686" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9355" daytime="15:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9356" daytime="15:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9357" daytime="16:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1246" daytime="15:24" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5255" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8999" />
                    <RANKING order="2" place="2" resultid="7603" />
                    <RANKING order="3" place="-1" resultid="7598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5256" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7976" />
                    <RANKING order="2" place="2" resultid="7596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5257" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7866" />
                    <RANKING order="2" place="-1" resultid="8388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5258" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6276" />
                    <RANKING order="2" place="2" resultid="7279" />
                    <RANKING order="3" place="3" resultid="7440" />
                    <RANKING order="4" place="4" resultid="6784" />
                    <RANKING order="5" place="-1" resultid="7867" />
                    <RANKING order="6" place="-1" resultid="7511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5259" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6524" />
                    <RANKING order="2" place="2" resultid="9000" />
                    <RANKING order="3" place="3" resultid="8698" />
                    <RANKING order="4" place="-1" resultid="5979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5260" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5261" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6937" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9353" daytime="15:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9354" daytime="15:28" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="14:12" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9623" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6618" />
                    <RANKING order="2" place="2" resultid="5835" />
                    <RANKING order="3" place="3" resultid="8886" />
                    <RANKING order="4" place="4" resultid="7546" />
                    <RANKING order="5" place="5" resultid="7959" />
                    <RANKING order="6" place="6" resultid="7701" />
                    <RANKING order="7" place="7" resultid="6365" />
                    <RANKING order="8" place="8" resultid="5842" />
                    <RANKING order="9" place="9" resultid="5674" />
                    <RANKING order="10" place="10" resultid="6038" />
                    <RANKING order="11" place="11" resultid="5750" />
                    <RANKING order="12" place="12" resultid="6854" />
                    <RANKING order="13" place="13" resultid="8310" />
                    <RANKING order="14" place="14" resultid="8654" />
                    <RANKING order="15" place="15" resultid="8316" />
                    <RANKING order="16" place="16" resultid="5734" />
                    <RANKING order="17" place="17" resultid="7577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9624" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7588" />
                    <RANKING order="2" place="2" resultid="6094" />
                    <RANKING order="3" place="3" resultid="6708" />
                    <RANKING order="4" place="4" resultid="8743" />
                    <RANKING order="5" place="5" resultid="7953" />
                    <RANKING order="6" place="6" resultid="8937" />
                    <RANKING order="7" place="7" resultid="6359" />
                    <RANKING order="8" place="8" resultid="8958" />
                    <RANKING order="9" place="9" resultid="6699" />
                    <RANKING order="10" place="10" resultid="7367" />
                    <RANKING order="11" place="11" resultid="7542" />
                    <RANKING order="12" place="12" resultid="7315" />
                    <RANKING order="13" place="13" resultid="7480" />
                    <RANKING order="14" place="14" resultid="7938" />
                    <RANKING order="15" place="15" resultid="8380" />
                    <RANKING order="16" place="-1" resultid="7102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9625" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6030" />
                    <RANKING order="2" place="2" resultid="7931" />
                    <RANKING order="3" place="3" resultid="6146" />
                    <RANKING order="4" place="4" resultid="7892" />
                    <RANKING order="5" place="5" resultid="7205" />
                    <RANKING order="6" place="6" resultid="7197" />
                    <RANKING order="7" place="7" resultid="7533" />
                    <RANKING order="8" place="8" resultid="7462" />
                    <RANKING order="9" place="9" resultid="7922" />
                    <RANKING order="10" place="10" resultid="6774" />
                    <RANKING order="11" place="11" resultid="7537" />
                    <RANKING order="12" place="12" resultid="8540" />
                    <RANKING order="13" place="13" resultid="7973" />
                    <RANKING order="14" place="14" resultid="8338" />
                    <RANKING order="15" place="15" resultid="7475" />
                    <RANKING order="16" place="16" resultid="8597" />
                    <RANKING order="17" place="17" resultid="7728" />
                    <RANKING order="18" place="18" resultid="8582" />
                    <RANKING order="19" place="-1" resultid="8384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9626" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6243" />
                    <RANKING order="2" place="2" resultid="7401" />
                    <RANKING order="3" place="3" resultid="8546" />
                    <RANKING order="4" place="4" resultid="8917" />
                    <RANKING order="5" place="5" resultid="7361" />
                    <RANKING order="6" place="6" resultid="7069" />
                    <RANKING order="7" place="7" resultid="6678" />
                    <RANKING order="8" place="8" resultid="7829" />
                    <RANKING order="9" place="9" resultid="7948" />
                    <RANKING order="10" place="10" resultid="5766" />
                    <RANKING order="11" place="11" resultid="7467" />
                    <RANKING order="12" place="12" resultid="7927" />
                    <RANKING order="13" place="13" resultid="8646" />
                    <RANKING order="14" place="14" resultid="6256" />
                    <RANKING order="15" place="15" resultid="6755" />
                    <RANKING order="16" place="-1" resultid="7320" />
                    <RANKING order="17" place="-1" resultid="8365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9627" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8944" />
                    <RANKING order="2" place="2" resultid="8923" />
                    <RANKING order="3" place="3" resultid="7435" />
                    <RANKING order="4" place="4" resultid="7943" />
                    <RANKING order="5" place="5" resultid="7855" />
                    <RANKING order="6" place="6" resultid="7822" />
                    <RANKING order="7" place="7" resultid="7456" />
                    <RANKING order="8" place="8" resultid="7773" />
                    <RANKING order="9" place="9" resultid="5774" />
                    <RANKING order="10" place="10" resultid="7247" />
                    <RANKING order="11" place="11" resultid="8759" />
                    <RANKING order="12" place="12" resultid="6068" />
                    <RANKING order="13" place="13" resultid="5762" />
                    <RANKING order="14" place="14" resultid="7255" />
                    <RANKING order="15" place="15" resultid="8574" />
                    <RANKING order="16" place="16" resultid="8750" />
                    <RANKING order="17" place="17" resultid="7910" />
                    <RANKING order="18" place="-1" resultid="7235" />
                    <RANKING order="19" place="-1" resultid="5804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9628" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6550" />
                    <RANKING order="2" place="2" resultid="5743" />
                    <RANKING order="3" place="3" resultid="6098" />
                    <RANKING order="4" place="4" resultid="8274" />
                    <RANKING order="5" place="5" resultid="6400" />
                    <RANKING order="6" place="6" resultid="7837" />
                    <RANKING order="7" place="7" resultid="6542" />
                    <RANKING order="8" place="8" resultid="6426" />
                    <RANKING order="9" place="9" resultid="5725" />
                    <RANKING order="10" place="10" resultid="7341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9629" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7491" />
                    <RANKING order="2" place="2" resultid="8012" />
                    <RANKING order="3" place="3" resultid="6198" />
                    <RANKING order="4" place="4" resultid="6345" />
                    <RANKING order="5" place="5" resultid="6602" />
                    <RANKING order="6" place="6" resultid="7861" />
                    <RANKING order="7" place="-1" resultid="7380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9630" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6153" />
                    <RANKING order="2" place="2" resultid="6084" />
                    <RANKING order="3" place="3" resultid="8869" />
                    <RANKING order="4" place="4" resultid="6863" />
                    <RANKING order="5" place="5" resultid="7663" />
                    <RANKING order="6" place="6" resultid="7768" />
                    <RANKING order="7" place="7" resultid="6484" />
                    <RANKING order="8" place="8" resultid="8026" />
                    <RANKING order="9" place="9" resultid="6830" />
                    <RANKING order="10" place="10" resultid="6402" />
                    <RANKING order="11" place="11" resultid="6004" />
                    <RANKING order="12" place="12" resultid="7168" />
                    <RANKING order="13" place="13" resultid="7389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9631" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8730" />
                    <RANKING order="2" place="2" resultid="8021" />
                    <RANKING order="3" place="3" resultid="5717" />
                    <RANKING order="4" place="4" resultid="6735" />
                    <RANKING order="5" place="5" resultid="6175" />
                    <RANKING order="6" place="6" resultid="6011" />
                    <RANKING order="7" place="7" resultid="6592" />
                    <RANKING order="8" place="8" resultid="6203" />
                    <RANKING order="9" place="-1" resultid="8706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9632" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7329" />
                    <RANKING order="2" place="2" resultid="8687" />
                    <RANKING order="3" place="3" resultid="6962" />
                    <RANKING order="4" place="4" resultid="8612" />
                    <RANKING order="5" place="-1" resultid="6110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9633" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6074" />
                    <RANKING order="2" place="2" resultid="6457" />
                    <RANKING order="3" place="3" resultid="5696" />
                    <RANKING order="4" place="4" resultid="6053" />
                    <RANKING order="5" place="5" resultid="7143" />
                    <RANKING order="6" place="6" resultid="8792" />
                    <RANKING order="7" place="7" resultid="6958" />
                    <RANKING order="8" place="-1" resultid="6236" />
                    <RANKING order="9" place="-1" resultid="8632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9634" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6916" />
                    <RANKING order="2" place="2" resultid="5975" />
                    <RANKING order="3" place="3" resultid="7123" />
                    <RANKING order="4" place="4" resultid="7149" />
                    <RANKING order="5" place="5" resultid="8621" />
                    <RANKING order="6" place="6" resultid="5778" />
                    <RANKING order="7" place="7" resultid="5787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9635" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6138" />
                    <RANKING order="2" place="2" resultid="8246" />
                    <RANKING order="3" place="3" resultid="8628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9636" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5902" />
                    <RANKING order="2" place="2" resultid="5934" />
                    <RANKING order="3" place="3" resultid="8428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9637" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9638" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9317" daytime="14:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9318" daytime="14:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9319" daytime="14:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9320" daytime="14:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9321" daytime="14:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9322" daytime="14:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9323" daytime="14:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9324" daytime="14:22" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9325" daytime="14:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9326" daytime="14:24" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9327" daytime="14:24" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9328" daytime="14:26" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9329" daytime="14:28" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="9330" daytime="14:28" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="9331" daytime="14:30" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="9332" daytime="14:30" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="14:32" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9639" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8895" />
                    <RANKING order="2" place="2" resultid="8990" />
                    <RANKING order="3" place="3" resultid="6562" />
                    <RANKING order="4" place="4" resultid="6719" />
                    <RANKING order="5" place="5" resultid="8806" />
                    <RANKING order="6" place="-1" resultid="7114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9640" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7580" />
                    <RANKING order="2" place="2" resultid="5925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9641" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8679" />
                    <RANKING order="2" place="2" resultid="7800" />
                    <RANKING order="3" place="3" resultid="7407" />
                    <RANKING order="4" place="-1" resultid="6353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9642" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6578" />
                    <RANKING order="2" place="2" resultid="8564" />
                    <RANKING order="3" place="3" resultid="8767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9643" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6382" />
                    <RANKING order="2" place="2" resultid="7272" />
                    <RANKING order="3" place="3" resultid="7887" />
                    <RANKING order="4" place="4" resultid="8291" />
                    <RANKING order="5" place="5" resultid="6509" />
                    <RANKING order="6" place="-1" resultid="6703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9644" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6229" />
                    <RANKING order="2" place="2" resultid="7291" />
                    <RANKING order="3" place="3" resultid="6492" />
                    <RANKING order="4" place="4" resultid="6018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9645" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6164" />
                    <RANKING order="2" place="2" resultid="6515" />
                    <RANKING order="3" place="3" resultid="7633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9646" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6335" />
                    <RANKING order="2" place="2" resultid="8900" />
                    <RANKING order="3" place="3" resultid="6632" />
                    <RANKING order="4" place="4" resultid="6475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9647" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7722" />
                    <RANKING order="2" place="2" resultid="5882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9648" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="9649" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9650" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9651" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9652" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9653" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9654" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9337" daytime="14:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9338" daytime="14:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9339" daytime="14:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9340" daytime="14:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1314" daytime="18:12" gender="M" number="9" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9719" agemax="24" agemin="20" name="Kat. 0" />
                <AGEGROUP agegroupid="9720" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7564" />
                    <RANKING order="2" place="-1" resultid="7047" />
                    <RANKING order="3" place="-1" resultid="7264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9721" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5859" />
                    <RANKING order="2" place="2" resultid="5819" />
                    <RANKING order="3" place="-1" resultid="8583" />
                    <RANKING order="4" place="-1" resultid="7729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9722" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9723" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9439" />
                    <RANKING order="2" place="2" resultid="8812" />
                    <RANKING order="3" place="3" resultid="5993" />
                    <RANKING order="4" place="4" resultid="6801" />
                    <RANKING order="5" place="5" resultid="7424" />
                    <RANKING order="6" place="6" resultid="7815" />
                    <RANKING order="7" place="7" resultid="7256" />
                    <RANKING order="8" place="-1" resultid="7748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9724" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6870" />
                    <RANKING order="2" place="2" resultid="7171" />
                    <RANKING order="3" place="3" resultid="9438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9725" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9726" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6831" />
                    <RANKING order="2" place="2" resultid="6121" />
                    <RANKING order="3" place="3" resultid="5998" />
                    <RANKING order="4" place="-1" resultid="8874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9727" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7054" />
                    <RANKING order="2" place="2" resultid="8707" />
                    <RANKING order="3" place="3" resultid="5944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9728" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7739" />
                    <RANKING order="2" place="2" resultid="5796" />
                    <RANKING order="3" place="-1" resultid="6584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9729" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9730" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9731" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9732" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9733" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9734" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9365" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9366" daytime="18:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9367" daytime="18:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9368" daytime="19:44" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1280" daytime="16:20" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9687" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6855" />
                    <RANKING order="2" place="2" resultid="9437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9688" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8639" />
                    <RANKING order="2" place="2" resultid="8713" />
                    <RANKING order="3" place="-1" resultid="5865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9689" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7893" />
                    <RANKING order="2" place="2" resultid="8659" />
                    <RANKING order="3" place="3" resultid="8598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9690" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8850" />
                    <RANKING order="2" place="2" resultid="7299" />
                    <RANKING order="3" place="3" resultid="8931" />
                    <RANKING order="4" place="4" resultid="7949" />
                    <RANKING order="5" place="-1" resultid="8647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9691" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8774" />
                    <RANKING order="2" place="2" resultid="7436" />
                    <RANKING order="3" place="3" resultid="7856" />
                    <RANKING order="4" place="4" resultid="7133" />
                    <RANKING order="5" place="5" resultid="8751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9692" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9435" />
                    <RANKING order="2" place="2" resultid="6099" />
                    <RANKING order="3" place="3" resultid="7240" />
                    <RANKING order="4" place="-1" resultid="6850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9693" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8842" />
                    <RANKING order="2" place="2" resultid="8013" />
                    <RANKING order="3" place="3" resultid="6346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9694" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6005" />
                    <RANKING order="2" place="2" resultid="6822" />
                    <RANKING order="3" place="3" resultid="7390" />
                    <RANKING order="4" place="4" resultid="8825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9695" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8731" />
                    <RANKING order="2" place="2" resultid="8261" />
                    <RANKING order="3" place="3" resultid="5718" />
                    <RANKING order="4" place="4" resultid="6012" />
                    <RANKING order="5" place="5" resultid="8964" />
                    <RANKING order="6" place="6" resultid="6176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9696" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8688" />
                    <RANKING order="2" place="2" resultid="6111" />
                    <RANKING order="3" place="3" resultid="8254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9697" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6458" />
                    <RANKING order="2" place="2" resultid="6410" />
                    <RANKING order="3" place="3" resultid="8793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9698" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9699" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9700" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9701" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9702" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9359" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9360" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9361" daytime="16:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9362" daytime="16:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9363" daytime="17:14" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-06-23" daytime="09:00" number="2">
          <EVENTS>
            <EVENT eventid="1476" daytime="09:14" gender="M" number="11" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9751" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6619" />
                    <RANKING order="2" place="2" resultid="7065" />
                    <RANKING order="3" place="3" resultid="6624" />
                    <RANKING order="4" place="4" resultid="5843" />
                    <RANKING order="5" place="5" resultid="8590" />
                    <RANKING order="6" place="-1" resultid="8317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9752" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7954" />
                    <RANKING order="2" place="2" resultid="7565" />
                    <RANKING order="3" place="3" resultid="6710" />
                    <RANKING order="4" place="4" resultid="8938" />
                    <RANKING order="5" place="4" resultid="8960" />
                    <RANKING order="6" place="6" resultid="7543" />
                    <RANKING order="7" place="7" resultid="7104" />
                    <RANKING order="8" place="-1" resultid="8381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9753" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7199" />
                    <RANKING order="2" place="2" resultid="7924" />
                    <RANKING order="3" place="3" resultid="8323" />
                    <RANKING order="4" place="4" resultid="6147" />
                    <RANKING order="5" place="5" resultid="7538" />
                    <RANKING order="6" place="6" resultid="6775" />
                    <RANKING order="7" place="7" resultid="8340" />
                    <RANKING order="8" place="8" resultid="7730" />
                    <RANKING order="9" place="9" resultid="8599" />
                    <RANKING order="10" place="10" resultid="7476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9754" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8367" />
                    <RANKING order="2" place="2" resultid="6264" />
                    <RANKING order="3" place="3" resultid="6245" />
                    <RANKING order="4" place="4" resultid="8547" />
                    <RANKING order="5" place="5" resultid="8695" />
                    <RANKING order="6" place="6" resultid="5970" />
                    <RANKING order="7" place="7" resultid="6680" />
                    <RANKING order="8" place="8" resultid="6744" />
                    <RANKING order="9" place="-1" resultid="7193" />
                    <RANKING order="10" place="-1" resultid="7322" />
                    <RANKING order="11" place="-1" resultid="8996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9755" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8925" />
                    <RANKING order="2" place="2" resultid="7904" />
                    <RANKING order="3" place="3" resultid="8952" />
                    <RANKING order="4" place="4" resultid="7816" />
                    <RANKING order="5" place="5" resultid="7857" />
                    <RANKING order="6" place="6" resultid="7760" />
                    <RANKING order="7" place="7" resultid="8760" />
                    <RANKING order="8" place="8" resultid="6802" />
                    <RANKING order="9" place="9" resultid="8752" />
                    <RANKING order="10" place="-1" resultid="7774" />
                    <RANKING order="11" place="-1" resultid="5805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9756" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7695" />
                    <RANKING order="2" place="2" resultid="6557" />
                    <RANKING order="3" place="3" resultid="7430" />
                    <RANKING order="4" place="4" resultid="5745" />
                    <RANKING order="5" place="5" resultid="6661" />
                    <RANKING order="6" place="6" resultid="8276" />
                    <RANKING order="7" place="7" resultid="5727" />
                    <RANKING order="8" place="8" resultid="8594" />
                    <RANKING order="9" place="-1" resultid="6428" />
                    <RANKING order="10" place="-1" resultid="7780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9757" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6062" />
                    <RANKING order="2" place="2" resultid="7382" />
                    <RANKING order="3" place="3" resultid="8843" />
                    <RANKING order="4" place="4" resultid="7862" />
                    <RANKING order="5" place="-1" resultid="8014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9758" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6154" />
                    <RANKING order="2" place="2" resultid="6086" />
                    <RANKING order="3" place="3" resultid="7664" />
                    <RANKING order="4" place="4" resultid="6864" />
                    <RANKING order="5" place="5" resultid="6485" />
                    <RANKING order="6" place="6" resultid="6652" />
                    <RANKING order="7" place="7" resultid="6893" />
                    <RANKING order="8" place="8" resultid="8267" />
                    <RANKING order="9" place="9" resultid="7769" />
                    <RANKING order="10" place="10" resultid="7169" />
                    <RANKING order="11" place="11" resultid="6403" />
                    <RANKING order="12" place="12" resultid="7391" />
                    <RANKING order="13" place="-1" resultid="6610" />
                    <RANKING order="14" place="-1" resultid="6832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9759" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8732" />
                    <RANKING order="2" place="2" resultid="6213" />
                    <RANKING order="3" place="3" resultid="8262" />
                    <RANKING order="4" place="4" resultid="5719" />
                    <RANKING order="5" place="5" resultid="6593" />
                    <RANKING order="6" place="6" resultid="6205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9760" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5797" />
                    <RANKING order="2" place="2" resultid="6112" />
                    <RANKING order="3" place="3" resultid="8255" />
                    <RANKING order="4" place="4" resultid="6963" />
                    <RANKING order="5" place="5" resultid="5891" />
                    <RANKING order="6" place="6" resultid="8614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9761" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5697" />
                    <RANKING order="2" place="2" resultid="6876" />
                    <RANKING order="3" place="3" resultid="6191" />
                    <RANKING order="4" place="4" resultid="8250" />
                    <RANKING order="5" place="5" resultid="5683" />
                    <RANKING order="6" place="6" resultid="8633" />
                    <RANKING order="7" place="7" resultid="6959" />
                    <RANKING order="8" place="8" resultid="8794" />
                    <RANKING order="9" place="9" resultid="7144" />
                    <RANKING order="10" place="10" resultid="5709" />
                    <RANKING order="11" place="-1" resultid="6237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9762" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7151" />
                    <RANKING order="2" place="2" resultid="7125" />
                    <RANKING order="3" place="3" resultid="5780" />
                    <RANKING order="4" place="4" resultid="8622" />
                    <RANKING order="5" place="5" resultid="5788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9763" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6139" />
                    <RANKING order="2" place="2" resultid="8247" />
                    <RANKING order="3" place="3" resultid="8629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9764" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5904" />
                    <RANKING order="2" place="2" resultid="5936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9765" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9766" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9447" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9448" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9449" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9450" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9451" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9452" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9453" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9454" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9455" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9456" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9457" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1612" daytime="12:12" gender="M" number="19" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5269" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="5270" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5271" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7984" />
                    <RANKING order="2" place="2" resultid="9002" />
                    <RANKING order="3" place="3" resultid="8700" />
                    <RANKING order="4" place="4" resultid="8386" />
                    <RANKING order="5" place="5" resultid="7443" />
                    <RANKING order="6" place="6" resultid="8601" />
                    <RANKING order="7" place="7" resultid="7983" />
                    <RANKING order="8" place="8" resultid="7509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5272" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9003" />
                    <RANKING order="2" place="2" resultid="7444" />
                    <RANKING order="3" place="3" resultid="7869" />
                    <RANKING order="4" place="4" resultid="7281" />
                    <RANKING order="5" place="5" resultid="6781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5273" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5274" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8294" />
                    <RANKING order="2" place="2" resultid="6283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5275" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6939" />
                    <RANKING order="2" place="2" resultid="8702" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9498" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9499" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="12:04" gender="F" number="18" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5262" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5263" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="5264" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7980" />
                    <RANKING order="2" place="2" resultid="6783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5265" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5266" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6522" />
                    <RANKING order="2" place="2" resultid="9001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5267" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL" />
                <AGEGROUP agegroupid="5268" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6938" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9497" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1544" daytime="10:56" gender="M" number="15" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9815" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8888" />
                    <RANKING order="2" place="2" resultid="6620" />
                    <RANKING order="3" place="3" resultid="7548" />
                    <RANKING order="4" place="4" resultid="5836" />
                    <RANKING order="5" place="5" resultid="7960" />
                    <RANKING order="6" place="6" resultid="6039" />
                    <RANKING order="7" place="7" resultid="5752" />
                    <RANKING order="8" place="8" resultid="6856" />
                    <RANKING order="9" place="9" resultid="8591" />
                    <RANKING order="10" place="10" resultid="8318" />
                    <RANKING order="11" place="11" resultid="8738" />
                    <RANKING order="12" place="12" resultid="8655" />
                    <RANKING order="13" place="13" resultid="5736" />
                    <RANKING order="14" place="14" resultid="8313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9816" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6095" />
                    <RANKING order="2" place="2" resultid="6711" />
                    <RANKING order="3" place="3" resultid="8744" />
                    <RANKING order="4" place="4" resultid="7368" />
                    <RANKING order="5" place="5" resultid="8939" />
                    <RANKING order="6" place="6" resultid="6360" />
                    <RANKING order="7" place="7" resultid="7964" />
                    <RANKING order="8" place="8" resultid="8961" />
                    <RANKING order="9" place="9" resultid="6700" />
                    <RANKING order="10" place="10" resultid="7317" />
                    <RANKING order="11" place="11" resultid="8716" />
                    <RANKING order="12" place="12" resultid="7939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9817" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7894" />
                    <RANKING order="2" place="2" resultid="7932" />
                    <RANKING order="3" place="3" resultid="6148" />
                    <RANKING order="4" place="4" resultid="7206" />
                    <RANKING order="5" place="5" resultid="7463" />
                    <RANKING order="6" place="6" resultid="7200" />
                    <RANKING order="7" place="7" resultid="8541" />
                    <RANKING order="8" place="8" resultid="7974" />
                    <RANKING order="9" place="9" resultid="8341" />
                    <RANKING order="10" place="10" resultid="8600" />
                    <RANKING order="11" place="11" resultid="7477" />
                    <RANKING order="12" place="12" resultid="8584" />
                    <RANKING order="13" place="-1" resultid="7731" />
                    <RANKING order="14" place="-1" resultid="8331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9818" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8548" />
                    <RANKING order="2" place="2" resultid="6246" />
                    <RANKING order="3" place="3" resultid="8918" />
                    <RANKING order="4" place="4" resultid="7300" />
                    <RANKING order="5" place="5" resultid="7831" />
                    <RANKING order="6" place="6" resultid="5767" />
                    <RANKING order="7" place="7" resultid="7950" />
                    <RANKING order="8" place="8" resultid="7470" />
                    <RANKING order="9" place="9" resultid="8648" />
                    <RANKING order="10" place="10" resultid="6756" />
                    <RANKING order="11" place="11" resultid="6745" />
                    <RANKING order="12" place="-1" resultid="6258" />
                    <RANKING order="13" place="-1" resultid="7323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9819" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8775" />
                    <RANKING order="2" place="2" resultid="8821" />
                    <RANKING order="3" place="3" resultid="8926" />
                    <RANKING order="4" place="4" resultid="7236" />
                    <RANKING order="5" place="5" resultid="8813" />
                    <RANKING order="6" place="6" resultid="7414" />
                    <RANKING order="7" place="7" resultid="6803" />
                    <RANKING order="8" place="8" resultid="7437" />
                    <RANKING order="9" place="9" resultid="7900" />
                    <RANKING order="10" place="10" resultid="7944" />
                    <RANKING order="11" place="11" resultid="7823" />
                    <RANKING order="12" place="12" resultid="7257" />
                    <RANKING order="13" place="13" resultid="7775" />
                    <RANKING order="14" place="14" resultid="7457" />
                    <RANKING order="15" place="15" resultid="8761" />
                    <RANKING order="16" place="16" resultid="5662" />
                    <RANKING order="17" place="17" resultid="8576" />
                    <RANKING order="18" place="18" resultid="7765" />
                    <RANKING order="19" place="19" resultid="8753" />
                    <RANKING order="20" place="20" resultid="7911" />
                    <RANKING order="21" place="21" resultid="8557" />
                    <RANKING order="22" place="-1" resultid="5806" />
                    <RANKING order="23" place="-1" resultid="7249" />
                    <RANKING order="24" place="-1" resultid="8946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9820" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7696" />
                    <RANKING order="2" place="2" resultid="5746" />
                    <RANKING order="3" place="3" resultid="6100" />
                    <RANKING order="4" place="4" resultid="6543" />
                    <RANKING order="5" place="5" resultid="7838" />
                    <RANKING order="6" place="6" resultid="8277" />
                    <RANKING order="7" place="7" resultid="7343" />
                    <RANKING order="8" place="8" resultid="7419" />
                    <RANKING order="9" place="9" resultid="6851" />
                    <RANKING order="10" place="-1" resultid="6371" />
                    <RANKING order="11" place="-1" resultid="6871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9821" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7493" />
                    <RANKING order="2" place="2" resultid="7383" />
                    <RANKING order="3" place="3" resultid="8015" />
                    <RANKING order="4" place="4" resultid="6199" />
                    <RANKING order="5" place="5" resultid="9304" />
                    <RANKING order="6" place="6" resultid="6603" />
                    <RANKING order="7" place="7" resultid="7863" />
                    <RANKING order="8" place="-1" resultid="6347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9822" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8870" />
                    <RANKING order="2" place="2" resultid="6087" />
                    <RANKING order="3" place="3" resultid="6865" />
                    <RANKING order="4" place="4" resultid="6833" />
                    <RANKING order="5" place="5" resultid="6894" />
                    <RANKING order="6" place="6" resultid="6404" />
                    <RANKING order="7" place="7" resultid="6006" />
                    <RANKING order="8" place="8" resultid="5999" />
                    <RANKING order="9" place="9" resultid="7392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9823" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6214" />
                    <RANKING order="2" place="2" resultid="8022" />
                    <RANKING order="3" place="3" resultid="5720" />
                    <RANKING order="4" place="4" resultid="8708" />
                    <RANKING order="5" place="5" resultid="6178" />
                    <RANKING order="6" place="6" resultid="5945" />
                    <RANKING order="7" place="7" resultid="6013" />
                    <RANKING order="8" place="8" resultid="5812" />
                    <RANKING order="9" place="9" resultid="6206" />
                    <RANKING order="10" place="10" resultid="6594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9824" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7330" />
                    <RANKING order="2" place="2" resultid="8689" />
                    <RANKING order="3" place="3" resultid="6964" />
                    <RANKING order="4" place="4" resultid="5892" />
                    <RANKING order="5" place="-1" resultid="6113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9825" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6076" />
                    <RANKING order="2" place="2" resultid="6459" />
                    <RANKING order="3" place="3" resultid="7145" />
                    <RANKING order="4" place="4" resultid="8795" />
                    <RANKING order="5" place="-1" resultid="6055" />
                    <RANKING order="6" place="-1" resultid="6238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9826" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6917" />
                    <RANKING order="2" place="2" resultid="7126" />
                    <RANKING order="3" place="3" resultid="5976" />
                    <RANKING order="4" place="4" resultid="7152" />
                    <RANKING order="5" place="5" resultid="8623" />
                    <RANKING order="6" place="6" resultid="5789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9827" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9828" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5905" />
                    <RANKING order="2" place="2" resultid="5937" />
                    <RANKING order="3" place="-1" resultid="8431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9829" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9830" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9477" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9478" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9479" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9480" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9481" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9482" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9483" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9484" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9485" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9486" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9487" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="9488" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="9489" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="9490" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1458" daytime="09:00" gender="F" number="10" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9735" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7591" />
                    <RANKING order="2" place="2" resultid="6720" />
                    <RANKING order="3" place="3" resultid="8970" />
                    <RANKING order="4" place="4" resultid="6563" />
                    <RANKING order="5" place="5" resultid="6106" />
                    <RANKING order="6" place="6" resultid="5825" />
                    <RANKING order="7" place="7" resultid="6571" />
                    <RANKING order="8" place="8" resultid="7115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9736" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6253" />
                    <RANKING order="2" place="2" resultid="6159" />
                    <RANKING order="3" place="3" resultid="8536" />
                    <RANKING order="4" place="4" resultid="7062" />
                    <RANKING order="5" place="5" resultid="7917" />
                    <RANKING order="6" place="6" resultid="6329" />
                    <RANKING order="7" place="7" resultid="7044" />
                    <RANKING order="8" place="8" resultid="6769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9737" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6388" />
                    <RANKING order="2" place="2" resultid="7936" />
                    <RANKING order="3" place="3" resultid="6762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9738" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8566" />
                    <RANKING order="2" place="2" resultid="8768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9739" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7888" />
                    <RANKING order="2" place="2" resultid="7220" />
                    <RANKING order="3" place="3" resultid="7842" />
                    <RANKING order="4" place="4" resultid="8788" />
                    <RANKING order="5" place="5" resultid="7228" />
                    <RANKING order="6" place="6" resultid="7273" />
                    <RANKING order="7" place="7" resultid="7571" />
                    <RANKING order="8" place="-1" resultid="6704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9740" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6230" />
                    <RANKING order="2" place="2" resultid="6672" />
                    <RANKING order="3" place="3" resultid="6436" />
                    <RANKING order="4" place="4" resultid="8354" />
                    <RANKING order="5" place="5" resultid="7211" />
                    <RANKING order="6" place="6" resultid="5920" />
                    <RANKING order="7" place="7" resultid="6694" />
                    <RANKING order="8" place="8" resultid="8667" />
                    <RANKING order="9" place="9" resultid="6493" />
                    <RANKING order="10" place="-1" resultid="6442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9741" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6420" />
                    <RANKING order="2" place="2" resultid="6731" />
                    <RANKING order="3" place="3" resultid="6516" />
                    <RANKING order="4" place="4" resultid="6666" />
                    <RANKING order="5" place="-1" resultid="8862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9742" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6271" />
                    <RANKING order="2" place="2" resultid="6337" />
                    <RANKING order="3" place="3" resultid="7628" />
                    <RANKING order="4" place="4" resultid="7848" />
                    <RANKING order="5" place="5" resultid="5953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9743" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6814" />
                    <RANKING order="2" place="2" resultid="6502" />
                    <RANKING order="3" place="3" resultid="5884" />
                    <RANKING order="4" place="4" resultid="5912" />
                    <RANKING order="5" place="5" resultid="8673" />
                    <RANKING order="6" place="6" resultid="7075" />
                    <RANKING order="7" place="7" resultid="6898" />
                    <RANKING order="8" place="-1" resultid="6725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9744" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8285" />
                    <RANKING order="2" place="2" resultid="7159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9745" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9746" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6921" />
                    <RANKING order="2" place="-1" resultid="8008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9747" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9748" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9749" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9750" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9440" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9441" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9442" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9443" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9444" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9445" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9446" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1561" daytime="11:30" gender="F" number="16" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9831" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8896" />
                    <RANKING order="2" place="2" resultid="7682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9832" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9833" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="9834" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="9835" agemax="44" agemin="40" name="Kat. D" />
                <AGEGROUP agegroupid="9836" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6231" />
                    <RANKING order="2" place="2" resultid="8355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9837" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9838" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6451" />
                    <RANKING order="2" place="2" resultid="6272" />
                    <RANKING order="3" place="3" resultid="6635" />
                    <RANKING order="4" place="4" resultid="6478" />
                    <RANKING order="5" place="-1" resultid="6338" />
                    <RANKING order="6" place="-1" resultid="8903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9839" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6503" />
                    <RANKING order="2" place="-1" resultid="5963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9840" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="9841" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="9842" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9843" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9844" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9845" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9846" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9491" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9492" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1493" daytime="09:34" gender="F" number="12" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9767" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8991" />
                    <RANKING order="2" place="2" resultid="7116" />
                    <RANKING order="3" place="3" resultid="8305" />
                    <RANKING order="4" place="4" resultid="8807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9768" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5926" />
                    <RANKING order="2" place="2" resultid="7558" />
                    <RANKING order="3" place="3" resultid="8977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9769" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8680" />
                    <RANKING order="2" place="2" resultid="7801" />
                    <RANKING order="3" place="3" resultid="8561" />
                    <RANKING order="4" place="4" resultid="7188" />
                    <RANKING order="5" place="-1" resultid="7305" />
                    <RANKING order="6" place="-1" resultid="8375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9770" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7403" />
                    <RANKING order="2" place="2" resultid="8347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9771" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8292" />
                    <RANKING order="2" place="2" resultid="7274" />
                    <RANKING order="3" place="3" resultid="8983" />
                    <RANKING order="4" place="4" resultid="6511" />
                    <RANKING order="5" place="5" resultid="8838" />
                    <RANKING order="6" place="-1" resultid="7640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9772" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6927" />
                    <RANKING order="2" place="2" resultid="7212" />
                    <RANKING order="3" place="3" resultid="7293" />
                    <RANKING order="4" place="4" resultid="6019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9773" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6165" />
                    <RANKING order="2" place="2" resultid="7355" />
                    <RANKING order="3" place="-1" resultid="7528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9774" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6220" />
                    <RANKING order="2" place="2" resultid="8902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9775" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8833" />
                    <RANKING order="2" place="2" resultid="8910" />
                    <RANKING order="3" place="3" resultid="5962" />
                    <RANKING order="4" place="-1" resultid="7076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9776" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8881" />
                    <RANKING order="2" place="2" resultid="5669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9777" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9778" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9779" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9780" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9781" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9782" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9458" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9459" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9460" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9461" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="11:40" gender="M" number="17" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9847" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6366" />
                    <RANKING order="2" place="2" resultid="7703" />
                    <RANKING order="3" place="3" resultid="6396" />
                    <RANKING order="4" place="-1" resultid="6625" />
                    <RANKING order="5" place="-1" resultid="8889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9848" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7566" />
                    <RANKING order="2" place="2" resultid="7048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9849" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5860" />
                    <RANKING order="2" place="2" resultid="8332" />
                    <RANKING order="3" place="3" resultid="8801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9850" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8852" />
                    <RANKING order="2" place="2" resultid="8368" />
                    <RANKING order="3" place="3" resultid="8932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9851" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5994" />
                    <RANKING order="2" place="2" resultid="7426" />
                    <RANKING order="3" place="3" resultid="7258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9852" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6535" />
                    <RANKING order="2" place="2" resultid="6551" />
                    <RANKING order="3" place="3" resultid="6372" />
                    <RANKING order="4" place="4" resultid="5691" />
                    <RANKING order="5" place="5" resultid="6101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9853" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7505" />
                    <RANKING order="2" place="2" resultid="7374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9854" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8826" />
                    <RANKING order="2" place="2" resultid="6122" />
                    <RANKING order="3" place="3" resultid="8875" />
                    <RANKING order="4" place="4" resultid="6611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9855" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7180" />
                    <RANKING order="2" place="2" resultid="6738" />
                    <RANKING order="3" place="-1" resultid="8733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9856" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5798" />
                    <RANKING order="2" place="2" resultid="6586" />
                    <RANKING order="3" place="3" resultid="8615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9857" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6077" />
                    <RANKING order="2" place="2" resultid="7717" />
                    <RANKING order="3" place="3" resultid="6412" />
                    <RANKING order="4" place="4" resultid="5684" />
                    <RANKING order="5" place="-1" resultid="6460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9858" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9859" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9860" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9861" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9862" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9493" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9494" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9495" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9496" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1527" daytime="10:34" gender="F" number="14" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9799" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6572" />
                    <RANKING order="2" place="2" resultid="6564" />
                    <RANKING order="3" place="3" resultid="7592" />
                    <RANKING order="4" place="4" resultid="5826" />
                    <RANKING order="5" place="5" resultid="8971" />
                    <RANKING order="6" place="6" resultid="8992" />
                    <RANKING order="7" place="7" resultid="8306" />
                    <RANKING order="8" place="8" resultid="7554" />
                    <RANKING order="9" place="9" resultid="7140" />
                    <RANKING order="10" place="-1" resultid="8808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9800" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7581" />
                    <RANKING order="2" place="2" resultid="7918" />
                    <RANKING order="3" place="3" resultid="5927" />
                    <RANKING order="4" place="-1" resultid="6254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9801" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6354" />
                    <RANKING order="2" place="2" resultid="8681" />
                    <RANKING order="3" place="3" resultid="7802" />
                    <RANKING order="4" place="4" resultid="5850" />
                    <RANKING order="5" place="5" resultid="6389" />
                    <RANKING order="6" place="6" resultid="7335" />
                    <RANKING order="7" place="7" resultid="7623" />
                    <RANKING order="8" place="8" resultid="6025" />
                    <RANKING order="9" place="9" resultid="6763" />
                    <RANKING order="10" place="10" resultid="6642" />
                    <RANKING order="11" place="11" resultid="6751" />
                    <RANKING order="12" place="-1" resultid="7306" />
                    <RANKING order="13" place="-1" resultid="8376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9802" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7310" />
                    <RANKING order="2" place="2" resultid="6579" />
                    <RANKING order="3" place="3" resultid="8567" />
                    <RANKING order="4" place="4" resultid="8769" />
                    <RANKING order="5" place="5" resultid="8348" />
                    <RANKING order="6" place="6" resultid="7486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9803" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6170" />
                    <RANKING order="2" place="2" resultid="7229" />
                    <RANKING order="3" place="3" resultid="7221" />
                    <RANKING order="4" place="4" resultid="7808" />
                    <RANKING order="5" place="5" resultid="7519" />
                    <RANKING order="6" place="6" resultid="7843" />
                    <RANKING order="7" place="7" resultid="7617" />
                    <RANKING order="8" place="8" resultid="8789" />
                    <RANKING order="9" place="9" resultid="8984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9804" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6437" />
                    <RANKING order="2" place="2" resultid="6695" />
                    <RANKING order="3" place="3" resultid="5921" />
                    <RANKING order="4" place="4" resultid="7294" />
                    <RANKING order="5" place="5" resultid="6494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9805" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6845" />
                    <RANKING order="2" place="2" resultid="6421" />
                    <RANKING order="3" place="3" resultid="6732" />
                    <RANKING order="4" place="4" resultid="7634" />
                    <RANKING order="5" place="5" resultid="8724" />
                    <RANKING order="6" place="6" resultid="6667" />
                    <RANKING order="7" place="-1" resultid="6517" />
                    <RANKING order="8" place="-1" resultid="8863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9806" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6450" />
                    <RANKING order="2" place="2" resultid="7629" />
                    <RANKING order="3" place="3" resultid="5954" />
                    <RANKING order="4" place="4" resultid="7849" />
                    <RANKING order="5" place="5" resultid="6316" />
                    <RANKING order="6" place="6" resultid="6634" />
                    <RANKING order="7" place="7" resultid="6477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9807" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6815" />
                    <RANKING order="2" place="2" resultid="5885" />
                    <RANKING order="3" place="3" resultid="8911" />
                    <RANKING order="4" place="4" resultid="5913" />
                    <RANKING order="5" place="5" resultid="8674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9808" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6902" />
                    <RANKING order="2" place="2" resultid="8882" />
                    <RANKING order="3" place="3" resultid="6186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9809" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9810" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9811" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9812" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9813" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9814" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9469" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9470" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9471" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9472" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9473" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9474" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9475" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9476" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1510" daytime="10:00" gender="M" number="13" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9783" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5844" />
                    <RANKING order="2" place="2" resultid="7514" />
                    <RANKING order="3" place="3" resultid="5676" />
                    <RANKING order="4" place="4" resultid="8312" />
                    <RANKING order="5" place="5" resultid="6395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9784" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8640" />
                    <RANKING order="2" place="2" resultid="7265" />
                    <RANKING order="3" place="3" resultid="8715" />
                    <RANKING order="4" place="-1" resultid="5866" />
                    <RANKING order="5" place="-1" resultid="7105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9785" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8660" />
                    <RANKING order="2" place="2" resultid="8324" />
                    <RANKING order="3" place="3" resultid="6776" />
                    <RANKING order="4" place="4" resultid="8800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9786" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7363" />
                    <RANKING order="2" place="2" resultid="8851" />
                    <RANKING order="3" place="3" resultid="7830" />
                    <RANKING order="4" place="4" resultid="6681" />
                    <RANKING order="5" place="5" resultid="7469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9787" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8820" />
                    <RANKING order="2" place="2" resultid="8945" />
                    <RANKING order="3" place="3" resultid="7425" />
                    <RANKING order="4" place="4" resultid="7749" />
                    <RANKING order="5" place="5" resultid="6129" />
                    <RANKING order="6" place="6" resultid="6069" />
                    <RANKING order="7" place="7" resultid="7248" />
                    <RANKING order="8" place="8" resultid="6688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9788" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6656" />
                    <RANKING order="2" place="2" resultid="7783" />
                    <RANKING order="3" place="3" resultid="6429" />
                    <RANKING order="4" place="4" resultid="7241" />
                    <RANKING order="5" place="5" resultid="5728" />
                    <RANKING order="6" place="6" resultid="6598" />
                    <RANKING order="7" place="7" resultid="7342" />
                    <RANKING order="8" place="8" resultid="8782" />
                    <RANKING order="9" place="9" resultid="7418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9789" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5987" />
                    <RANKING order="2" place="2" resultid="7504" />
                    <RANKING order="3" place="3" resultid="8270" />
                    <RANKING order="4" place="4" resultid="9303" />
                    <RANKING order="5" place="5" resultid="7373" />
                    <RANKING order="6" place="6" resultid="5702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9790" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8027" />
                    <RANKING order="2" place="2" resultid="7499" />
                    <RANKING order="3" place="3" resultid="6824" />
                    <RANKING order="4" place="4" resultid="6260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9791" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7179" />
                    <RANKING order="2" place="2" resultid="6737" />
                    <RANKING order="3" place="3" resultid="6177" />
                    <RANKING order="4" place="-1" resultid="6323" />
                    <RANKING order="5" place="-1" resultid="8241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9792" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7350" />
                    <RANKING order="2" place="2" resultid="7163" />
                    <RANKING order="3" place="3" resultid="7740" />
                    <RANKING order="4" place="4" resultid="6810" />
                    <RANKING order="5" place="5" resultid="6225" />
                    <RANKING order="6" place="6" resultid="6585" />
                    <RANKING order="7" place="7" resultid="5898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9793" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6192" />
                    <RANKING order="2" place="2" resultid="8634" />
                    <RANKING order="3" place="3" resultid="6411" />
                    <RANKING order="4" place="4" resultid="5710" />
                    <RANKING order="5" place="-1" resultid="7788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9794" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9795" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9796" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9797" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9798" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9462" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9463" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9464" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9465" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9466" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9467" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9468" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-06-23" daytime="15:00" endtime="19:05" number="3">
          <EVENTS>
            <EVENT eventid="5399" daytime="16:56" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9975" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8890" />
                    <RANKING order="2" place="2" resultid="7704" />
                    <RANKING order="3" place="3" resultid="7550" />
                    <RANKING order="4" place="4" resultid="6858" />
                    <RANKING order="5" place="5" resultid="8740" />
                    <RANKING order="6" place="6" resultid="5739" />
                    <RANKING order="7" place="-1" resultid="8320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9976" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8746" />
                    <RANKING order="2" place="2" resultid="6362" />
                    <RANKING order="3" place="3" resultid="7370" />
                    <RANKING order="4" place="4" resultid="8941" />
                    <RANKING order="5" place="5" resultid="8718" />
                    <RANKING order="6" place="6" resultid="7941" />
                    <RANKING order="7" place="7" resultid="8554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9977" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7896" />
                    <RANKING order="2" place="2" resultid="7933" />
                    <RANKING order="3" place="3" resultid="8662" />
                    <RANKING order="4" place="4" resultid="8586" />
                    <RANKING order="5" place="-1" resultid="5861" />
                    <RANKING order="6" place="-1" resultid="7733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9978" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8853" />
                    <RANKING order="2" place="2" resultid="7301" />
                    <RANKING order="3" place="3" resultid="5769" />
                    <RANKING order="4" place="4" resultid="7833" />
                    <RANKING order="5" place="5" resultid="7951" />
                    <RANKING order="6" place="6" resultid="8933" />
                    <RANKING order="7" place="7" resultid="8650" />
                    <RANKING order="8" place="8" resultid="7929" />
                    <RANKING order="9" place="9" resultid="6757" />
                    <RANKING order="10" place="-1" resultid="7324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9979" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8776" />
                    <RANKING order="2" place="2" resultid="7237" />
                    <RANKING order="3" place="3" resultid="7415" />
                    <RANKING order="4" place="4" resultid="8954" />
                    <RANKING order="5" place="5" resultid="8814" />
                    <RANKING order="6" place="6" resultid="7438" />
                    <RANKING order="7" place="7" resultid="6805" />
                    <RANKING order="8" place="8" resultid="7825" />
                    <RANKING order="9" place="9" resultid="7901" />
                    <RANKING order="10" place="10" resultid="7259" />
                    <RANKING order="11" place="11" resultid="8763" />
                    <RANKING order="12" place="12" resultid="5664" />
                    <RANKING order="13" place="13" resultid="8578" />
                    <RANKING order="14" place="14" resultid="8755" />
                    <RANKING order="15" place="15" resultid="6690" />
                    <RANKING order="16" place="16" resultid="8558" />
                    <RANKING order="17" place="17" resultid="7913" />
                    <RANKING order="18" place="-1" resultid="7946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9980" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6536" />
                    <RANKING order="2" place="2" resultid="6872" />
                    <RANKING order="3" place="3" resultid="6103" />
                    <RANKING order="4" place="4" resultid="7432" />
                    <RANKING order="5" place="5" resultid="5693" />
                    <RANKING order="6" place="6" resultid="6545" />
                    <RANKING order="7" place="7" resultid="8279" />
                    <RANKING order="8" place="8" resultid="7173" />
                    <RANKING order="9" place="9" resultid="5730" />
                    <RANKING order="10" place="10" resultid="7345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9981" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7494" />
                    <RANKING order="2" place="2" resultid="6647" />
                    <RANKING order="3" place="3" resultid="6064" />
                    <RANKING order="4" place="4" resultid="8845" />
                    <RANKING order="5" place="5" resultid="7670" />
                    <RANKING order="6" place="6" resultid="8017" />
                    <RANKING order="7" place="7" resultid="7376" />
                    <RANKING order="8" place="8" resultid="5704" />
                    <RANKING order="9" place="-1" resultid="6348" />
                    <RANKING order="10" place="-1" resultid="6605" />
                    <RANKING order="11" place="-1" resultid="9306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9982" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8871" />
                    <RANKING order="2" place="2" resultid="6867" />
                    <RANKING order="3" place="3" resultid="6835" />
                    <RANKING order="4" place="4" resultid="6008" />
                    <RANKING order="5" place="5" resultid="8828" />
                    <RANKING order="6" place="6" resultid="7394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9983" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6216" />
                    <RANKING order="2" place="2" resultid="8710" />
                    <RANKING order="3" place="3" resultid="5721" />
                    <RANKING order="4" place="4" resultid="6180" />
                    <RANKING order="5" place="5" resultid="6014" />
                    <RANKING order="6" place="6" resultid="5946" />
                    <RANKING order="7" place="7" resultid="8966" />
                    <RANKING order="8" place="8" resultid="5814" />
                    <RANKING order="9" place="9" resultid="6208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9984" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7332" />
                    <RANKING order="2" place="2" resultid="7741" />
                    <RANKING order="3" place="3" resultid="8691" />
                    <RANKING order="4" place="4" resultid="5894" />
                    <RANKING order="5" place="5" resultid="8616" />
                    <RANKING order="6" place="6" resultid="5900" />
                    <RANKING order="7" place="-1" resultid="6115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9985" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6462" />
                    <RANKING order="2" place="2" resultid="6056" />
                    <RANKING order="3" place="3" resultid="8796" />
                    <RANKING order="4" place="4" resultid="5686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9986" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6918" />
                    <RANKING order="2" place="2" resultid="7128" />
                    <RANKING order="3" place="3" resultid="5978" />
                    <RANKING order="4" place="4" resultid="8625" />
                    <RANKING order="5" place="5" resultid="5791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9987" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9988" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5939" />
                    <RANKING order="2" place="2" resultid="8433" />
                    <RANKING order="3" place="-1" resultid="5907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9989" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9990" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9548" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9549" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9550" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9551" daytime="17:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9552" daytime="17:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9553" daytime="17:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9554" daytime="17:22" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9555" daytime="17:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9556" daytime="17:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9557" daytime="17:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9558" daytime="17:34" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5314" daytime="15:36" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9895" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7593" />
                    <RANKING order="2" place="2" resultid="6565" />
                    <RANKING order="3" place="3" resultid="8972" />
                    <RANKING order="4" place="4" resultid="6573" />
                    <RANKING order="5" place="5" resultid="8809" />
                    <RANKING order="6" place="-1" resultid="6721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9896" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7063" />
                    <RANKING order="2" place="2" resultid="6331" />
                    <RANKING order="3" place="3" resultid="7560" />
                    <RANKING order="4" place="4" resultid="7919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9897" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6355" />
                    <RANKING order="2" place="2" resultid="7409" />
                    <RANKING order="3" place="3" resultid="7336" />
                    <RANKING order="4" place="4" resultid="6390" />
                    <RANKING order="5" place="5" resultid="6026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9898" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6580" />
                    <RANKING order="2" place="2" resultid="7311" />
                    <RANKING order="3" place="3" resultid="7969" />
                    <RANKING order="4" place="4" resultid="8770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9899" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7618" />
                    <RANKING order="2" place="2" resultid="7230" />
                    <RANKING order="3" place="3" resultid="7521" />
                    <RANKING order="4" place="4" resultid="6512" />
                    <RANKING order="5" place="-1" resultid="7642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9900" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6232" />
                    <RANKING order="2" place="2" resultid="6438" />
                    <RANKING order="3" place="3" resultid="6443" />
                    <RANKING order="4" place="4" resultid="6696" />
                    <RANKING order="5" place="5" resultid="6495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9901" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6422" />
                    <RANKING order="2" place="2" resultid="7635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9902" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6273" />
                    <RANKING order="2" place="2" resultid="6452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9903" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7724" />
                    <RANKING order="2" place="2" resultid="5964" />
                    <RANKING order="3" place="3" resultid="5886" />
                    <RANKING order="4" place="4" resultid="5914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9904" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9905" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9906" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9907" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9908" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9909" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9910" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9514" daytime="15:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9515" daytime="15:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9516" daytime="15:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9517" daytime="15:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5279" daytime="15:00" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9863" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8993" />
                    <RANKING order="2" place="2" resultid="7117" />
                    <RANKING order="3" place="3" resultid="8307" />
                    <RANKING order="4" place="4" resultid="7574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9864" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6330" />
                    <RANKING order="2" place="2" resultid="7559" />
                    <RANKING order="3" place="3" resultid="8978" />
                    <RANKING order="4" place="4" resultid="6770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9865" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8682" />
                    <RANKING order="2" place="2" resultid="5851" />
                    <RANKING order="3" place="3" resultid="7307" />
                    <RANKING order="4" place="4" resultid="7803" />
                    <RANKING order="5" place="-1" resultid="7624" />
                    <RANKING order="6" place="-1" resultid="8377" />
                    <RANKING order="7" place="-1" resultid="8562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9866" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8349" />
                    <RANKING order="2" place="2" resultid="7404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9867" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8293" />
                    <RANKING order="2" place="2" resultid="7275" />
                    <RANKING order="3" place="3" resultid="7520" />
                    <RANKING order="4" place="4" resultid="7809" />
                    <RANKING order="5" place="5" resultid="8839" />
                    <RANKING order="6" place="6" resultid="8985" />
                    <RANKING order="7" place="-1" resultid="7641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9868" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6928" />
                    <RANKING order="2" place="2" resultid="7213" />
                    <RANKING order="3" place="3" resultid="7295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9869" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6166" />
                    <RANKING order="2" place="2" resultid="7356" />
                    <RANKING order="3" place="3" resultid="6668" />
                    <RANKING order="4" place="4" resultid="6518" />
                    <RANKING order="5" place="-1" resultid="7529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9870" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6221" />
                    <RANKING order="2" place="2" resultid="8904" />
                    <RANKING order="3" place="3" resultid="5955" />
                    <RANKING order="4" place="4" resultid="7850" />
                    <RANKING order="5" place="5" resultid="6479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9871" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8834" />
                    <RANKING order="2" place="2" resultid="7723" />
                    <RANKING order="3" place="3" resultid="8912" />
                    <RANKING order="4" place="-1" resultid="7077" />
                    <RANKING order="5" place="-1" resultid="6726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9872" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8883" />
                    <RANKING order="2" place="2" resultid="5670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9873" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9874" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9875" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9876" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9877" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9878" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9500" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9501" daytime="15:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9502" daytime="15:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9503" daytime="15:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9504" daytime="15:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5433" daytime="17:42" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5491" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="5492" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7981" />
                    <RANKING order="2" place="-1" resultid="7599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5493" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7441" />
                    <RANKING order="2" place="2" resultid="8387" />
                    <RANKING order="3" place="3" resultid="8701" />
                    <RANKING order="4" place="4" resultid="7982" />
                    <RANKING order="5" place="5" resultid="8602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5494" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9005" />
                    <RANKING order="2" place="2" resultid="9010" />
                    <RANKING order="3" place="3" resultid="7871" />
                    <RANKING order="4" place="4" resultid="7282" />
                    <RANKING order="5" place="5" resultid="6782" />
                    <RANKING order="6" place="-1" resultid="7508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5495" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5496" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5497" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6941" />
                    <RANKING order="2" place="2" resultid="8703" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9560" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9561" daytime="17:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5450" daytime="17:50" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9991" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8994" />
                    <RANKING order="2" place="2" resultid="7683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9992" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9993" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7804" />
                    <RANKING order="2" place="-1" resultid="7410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9994" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="8350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9995" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6378" />
                    <RANKING order="2" place="2" resultid="7276" />
                    <RANKING order="3" place="3" resultid="7620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9996" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8357" />
                    <RANKING order="2" place="2" resultid="6444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9997" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7525" />
                    <RANKING order="2" place="2" resultid="6519" />
                    <RANKING order="3" place="3" resultid="8726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9998" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6340" />
                    <RANKING order="2" place="2" resultid="7851" />
                    <RANKING order="3" place="3" resultid="8905" />
                    <RANKING order="4" place="4" resultid="6637" />
                    <RANKING order="5" place="5" resultid="6480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9999" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10000" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="10001" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="10002" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="10003" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10004" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10005" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10006" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9562" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9563" daytime="18:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5416" daytime="17:38" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5484" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5485" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL" />
                <AGEGROUP agegroupid="5486" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7979" />
                    <RANKING order="2" place="2" resultid="6780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5487" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7870" />
                    <RANKING order="2" place="2" resultid="9006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5488" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5489" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5490" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6940" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9559" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5382" daytime="16:30" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9959" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7594" />
                    <RANKING order="2" place="2" resultid="6574" />
                    <RANKING order="3" place="3" resultid="6566" />
                    <RANKING order="4" place="4" resultid="5828" />
                    <RANKING order="5" place="5" resultid="8810" />
                    <RANKING order="6" place="-1" resultid="8308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9960" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5928" />
                    <RANKING order="2" place="2" resultid="7059" />
                    <RANKING order="3" place="3" resultid="8979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9961" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8683" />
                    <RANKING order="2" place="2" resultid="7337" />
                    <RANKING order="3" place="3" resultid="7190" />
                    <RANKING order="4" place="4" resultid="6027" />
                    <RANKING order="5" place="5" resultid="6643" />
                    <RANKING order="6" place="6" resultid="6752" />
                    <RANKING order="7" place="-1" resultid="6765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9962" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6312" />
                    <RANKING order="2" place="2" resultid="8569" />
                    <RANKING order="3" place="3" resultid="7487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9963" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6171" />
                    <RANKING order="2" place="2" resultid="7223" />
                    <RANKING order="3" place="3" resultid="6384" />
                    <RANKING order="4" place="4" resultid="7231" />
                    <RANKING order="5" place="5" resultid="7810" />
                    <RANKING order="6" place="6" resultid="6513" />
                    <RANKING order="7" place="-1" resultid="7619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9964" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6929" />
                    <RANKING order="2" place="2" resultid="7214" />
                    <RANKING order="3" place="3" resultid="5922" />
                    <RANKING order="4" place="4" resultid="7296" />
                    <RANKING order="5" place="5" resultid="6020" />
                    <RANKING order="6" place="-1" resultid="6496" />
                    <RANKING order="7" place="-1" resultid="6697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9965" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6846" />
                    <RANKING order="2" place="2" resultid="8725" />
                    <RANKING order="3" place="3" resultid="7357" />
                    <RANKING order="4" place="4" resultid="7636" />
                    <RANKING order="5" place="5" resultid="6669" />
                    <RANKING order="6" place="-1" resultid="8865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9966" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7630" />
                    <RANKING order="2" place="2" resultid="6453" />
                    <RANKING order="3" place="3" resultid="6222" />
                    <RANKING order="4" place="4" resultid="5956" />
                    <RANKING order="5" place="-1" resultid="6318" />
                    <RANKING order="6" place="-1" resultid="6636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9967" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6817" />
                    <RANKING order="2" place="2" resultid="5965" />
                    <RANKING order="3" place="3" resultid="5915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9968" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8287" />
                    <RANKING order="2" place="2" resultid="6187" />
                    <RANKING order="3" place="3" resultid="7398" />
                    <RANKING order="4" place="-1" resultid="6903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9969" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="9970" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="9971" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9972" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9973" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9974" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9542" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9543" daytime="16:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9544" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9545" daytime="16:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9546" daytime="16:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9547" daytime="16:52" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5467" daytime="18:08" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10007" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7705" />
                    <RANKING order="2" place="2" resultid="6397" />
                    <RANKING order="3" place="-1" resultid="8891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10008" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8642" />
                    <RANKING order="2" place="2" resultid="7049" />
                    <RANKING order="3" place="-1" resultid="5856" />
                    <RANKING order="4" place="-1" resultid="7267" />
                    <RANKING order="5" place="-1" resultid="7568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10009" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6134" />
                    <RANKING order="2" place="2" resultid="8334" />
                    <RANKING order="3" place="3" resultid="8326" />
                    <RANKING order="4" place="-1" resultid="5862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10010" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8854" />
                    <RANKING order="2" place="2" resultid="6683" />
                    <RANKING order="3" place="-1" resultid="7325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10011" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8777" />
                    <RANKING order="2" place="2" resultid="8815" />
                    <RANKING order="3" place="3" resultid="5995" />
                    <RANKING order="4" place="4" resultid="7762" />
                    <RANKING order="5" place="5" resultid="7751" />
                    <RANKING order="6" place="6" resultid="7260" />
                    <RANKING order="7" place="-1" resultid="6048" />
                    <RANKING order="8" place="-1" resultid="7427" />
                    <RANKING order="9" place="-1" resultid="7818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10012" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6537" />
                    <RANKING order="2" place="2" resultid="7698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10013" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7495" />
                    <RANKING order="2" place="2" resultid="7506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10014" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6124" />
                    <RANKING order="2" place="2" resultid="6044" />
                    <RANKING order="3" place="3" resultid="6613" />
                    <RANKING order="4" place="4" resultid="6000" />
                    <RANKING order="5" place="-1" resultid="8876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10015" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7182" />
                    <RANKING order="2" place="2" resultid="8264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10016" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7742" />
                    <RANKING order="2" place="2" resultid="7352" />
                    <RANKING order="3" place="3" resultid="5800" />
                    <RANKING order="4" place="4" resultid="8617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10017" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6079" />
                    <RANKING order="2" place="2" resultid="7718" />
                    <RANKING order="3" place="3" resultid="6414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10018" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10019" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10020" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10021" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10022" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9564" daytime="18:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9565" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9566" daytime="18:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9567" daytime="18:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9568" daytime="18:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5297" daytime="15:14" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9879" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7515" />
                    <RANKING order="2" place="2" resultid="5845" />
                    <RANKING order="3" place="3" resultid="5837" />
                    <RANKING order="4" place="4" resultid="5753" />
                    <RANKING order="5" place="5" resultid="5677" />
                    <RANKING order="6" place="6" resultid="5737" />
                    <RANKING order="7" place="7" resultid="8314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9880" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7755" />
                    <RANKING order="2" place="2" resultid="5867" />
                    <RANKING order="3" place="3" resultid="8641" />
                    <RANKING order="4" place="4" resultid="7965" />
                    <RANKING order="5" place="5" resultid="6361" />
                    <RANKING order="6" place="5" resultid="7481" />
                    <RANKING order="7" place="7" resultid="7266" />
                    <RANKING order="8" place="-1" resultid="7106" />
                    <RANKING order="9" place="-1" resultid="7544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9881" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6031" />
                    <RANKING order="2" place="2" resultid="8661" />
                    <RANKING order="3" place="3" resultid="8333" />
                    <RANKING order="4" place="4" resultid="7539" />
                    <RANKING order="5" place="5" resultid="8542" />
                    <RANKING order="6" place="6" resultid="6777" />
                    <RANKING order="7" place="7" resultid="8802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9882" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8919" />
                    <RANKING order="2" place="2" resultid="6247" />
                    <RANKING order="3" place="3" resultid="7364" />
                    <RANKING order="4" place="4" resultid="7832" />
                    <RANKING order="5" place="5" resultid="7471" />
                    <RANKING order="6" place="6" resultid="6746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9883" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8822" />
                    <RANKING order="2" place="2" resultid="8947" />
                    <RANKING order="3" place="3" resultid="7905" />
                    <RANKING order="4" place="4" resultid="7750" />
                    <RANKING order="5" place="5" resultid="6130" />
                    <RANKING order="6" place="6" resultid="6070" />
                    <RANKING order="7" place="7" resultid="7250" />
                    <RANKING order="8" place="8" resultid="6689" />
                    <RANKING order="9" place="9" resultid="7458" />
                    <RANKING order="10" place="10" resultid="7766" />
                    <RANKING order="11" place="-1" resultid="7134" />
                    <RANKING order="12" place="-1" resultid="7824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9884" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6657" />
                    <RANKING order="2" place="2" resultid="7784" />
                    <RANKING order="3" place="3" resultid="7242" />
                    <RANKING order="4" place="4" resultid="6430" />
                    <RANKING order="5" place="5" resultid="7344" />
                    <RANKING order="6" place="6" resultid="6599" />
                    <RANKING order="7" place="7" resultid="7420" />
                    <RANKING order="8" place="-1" resultid="7781" />
                    <RANKING order="9" place="-1" resultid="8783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9885" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6307" />
                    <RANKING order="2" place="2" resultid="8271" />
                    <RANKING order="3" place="3" resultid="5988" />
                    <RANKING order="4" place="4" resultid="7669" />
                    <RANKING order="5" place="5" resultid="7375" />
                    <RANKING order="6" place="6" resultid="6604" />
                    <RANKING order="7" place="7" resultid="5703" />
                    <RANKING order="8" place="-1" resultid="9305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9886" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8028" />
                    <RANKING order="2" place="2" resultid="7500" />
                    <RANKING order="3" place="3" resultid="6825" />
                    <RANKING order="4" place="4" resultid="6261" />
                    <RANKING order="5" place="5" resultid="6405" />
                    <RANKING order="6" place="-1" resultid="8298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9887" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7181" />
                    <RANKING order="2" place="2" resultid="6739" />
                    <RANKING order="3" place="3" resultid="6324" />
                    <RANKING order="4" place="4" resultid="6179" />
                    <RANKING order="5" place="5" resultid="8242" />
                    <RANKING order="6" place="6" resultid="8965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9888" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7351" />
                    <RANKING order="2" place="2" resultid="7164" />
                    <RANKING order="3" place="3" resultid="6811" />
                    <RANKING order="4" place="4" resultid="6226" />
                    <RANKING order="5" place="5" resultid="6587" />
                    <RANKING order="6" place="6" resultid="5899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9889" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6193" />
                    <RANKING order="2" place="2" resultid="8635" />
                    <RANKING order="3" place="3" resultid="5711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9890" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6907" />
                    <RANKING order="2" place="2" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9891" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9892" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5906" />
                    <RANKING order="2" place="2" resultid="8432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9893" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9894" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9505" daytime="15:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9506" daytime="15:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9507" daytime="15:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9508" daytime="15:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9509" daytime="15:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9510" daytime="15:28" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9511" daytime="15:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9512" daytime="15:32" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9513" daytime="15:34" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5331" daytime="15:44" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9911" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6621" />
                    <RANKING order="2" place="2" resultid="7549" />
                    <RANKING order="3" place="3" resultid="7961" />
                    <RANKING order="4" place="4" resultid="6367" />
                    <RANKING order="5" place="5" resultid="5838" />
                    <RANKING order="6" place="6" resultid="6626" />
                    <RANKING order="7" place="7" resultid="5846" />
                    <RANKING order="8" place="8" resultid="6040" />
                    <RANKING order="9" place="9" resultid="6857" />
                    <RANKING order="10" place="10" resultid="8739" />
                    <RANKING order="11" place="11" resultid="5754" />
                    <RANKING order="12" place="12" resultid="8656" />
                    <RANKING order="13" place="13" resultid="5678" />
                    <RANKING order="14" place="14" resultid="5738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9912" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7589" />
                    <RANKING order="2" place="2" resultid="8745" />
                    <RANKING order="3" place="3" resultid="7955" />
                    <RANKING order="4" place="4" resultid="6712" />
                    <RANKING order="5" place="5" resultid="7369" />
                    <RANKING order="6" place="6" resultid="8940" />
                    <RANKING order="7" place="7" resultid="7318" />
                    <RANKING order="8" place="8" resultid="6701" />
                    <RANKING order="9" place="9" resultid="8717" />
                    <RANKING order="10" place="10" resultid="7482" />
                    <RANKING order="11" place="11" resultid="7940" />
                    <RANKING order="12" place="-1" resultid="7756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9913" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7895" />
                    <RANKING order="2" place="2" resultid="7534" />
                    <RANKING order="3" place="3" resultid="7925" />
                    <RANKING order="4" place="4" resultid="7201" />
                    <RANKING order="5" place="5" resultid="7464" />
                    <RANKING order="6" place="6" resultid="8342" />
                    <RANKING order="7" place="7" resultid="7975" />
                    <RANKING order="8" place="8" resultid="7478" />
                    <RANKING order="9" place="9" resultid="8803" />
                    <RANKING order="10" place="10" resultid="8385" />
                    <RANKING order="11" place="-1" resultid="6149" />
                    <RANKING order="12" place="-1" resultid="8585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9914" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8369" />
                    <RANKING order="2" place="2" resultid="8920" />
                    <RANKING order="3" place="3" resultid="6265" />
                    <RANKING order="4" place="4" resultid="6248" />
                    <RANKING order="5" place="5" resultid="8549" />
                    <RANKING order="6" place="6" resultid="7070" />
                    <RANKING order="7" place="7" resultid="5971" />
                    <RANKING order="8" place="8" resultid="8649" />
                    <RANKING order="9" place="9" resultid="5768" />
                    <RANKING order="10" place="10" resultid="7472" />
                    <RANKING order="11" place="11" resultid="7928" />
                    <RANKING order="12" place="12" resultid="6747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9915" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8823" />
                    <RANKING order="2" place="2" resultid="7135" />
                    <RANKING order="3" place="3" resultid="8948" />
                    <RANKING order="4" place="4" resultid="7945" />
                    <RANKING order="5" place="5" resultid="5763" />
                    <RANKING order="6" place="6" resultid="5775" />
                    <RANKING order="7" place="7" resultid="8577" />
                    <RANKING order="8" place="8" resultid="5663" />
                    <RANKING order="9" place="9" resultid="7459" />
                    <RANKING order="10" place="10" resultid="8754" />
                    <RANKING order="11" place="11" resultid="7912" />
                    <RANKING order="12" place="-1" resultid="5807" />
                    <RANKING order="13" place="-1" resultid="7251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9916" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6552" />
                    <RANKING order="2" place="2" resultid="6658" />
                    <RANKING order="3" place="3" resultid="7431" />
                    <RANKING order="4" place="4" resultid="5692" />
                    <RANKING order="5" place="5" resultid="6102" />
                    <RANKING order="6" place="6" resultid="6373" />
                    <RANKING order="7" place="7" resultid="6662" />
                    <RANKING order="8" place="8" resultid="6544" />
                    <RANKING order="9" place="9" resultid="8278" />
                    <RANKING order="10" place="10" resultid="7839" />
                    <RANKING order="11" place="11" resultid="5729" />
                    <RANKING order="12" place="12" resultid="7172" />
                    <RANKING order="13" place="13" resultid="7421" />
                    <RANKING order="14" place="-1" resultid="7243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9917" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6063" />
                    <RANKING order="2" place="2" resultid="7384" />
                    <RANKING order="3" place="3" resultid="6200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9918" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6088" />
                    <RANKING order="2" place="2" resultid="6486" />
                    <RANKING order="3" place="3" resultid="6866" />
                    <RANKING order="4" place="4" resultid="8827" />
                    <RANKING order="5" place="5" resultid="6007" />
                    <RANKING order="6" place="6" resultid="7393" />
                    <RANKING order="7" place="-1" resultid="6123" />
                    <RANKING order="8" place="-1" resultid="8299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9919" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8023" />
                    <RANKING order="2" place="2" resultid="6215" />
                    <RANKING order="3" place="3" resultid="9300" />
                    <RANKING order="4" place="4" resultid="5813" />
                    <RANKING order="5" place="5" resultid="6595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9920" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8690" />
                    <RANKING order="2" place="2" resultid="6965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9921" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6078" />
                    <RANKING order="2" place="2" resultid="6461" />
                    <RANKING order="3" place="3" resultid="7146" />
                    <RANKING order="4" place="4" resultid="5685" />
                    <RANKING order="5" place="5" resultid="6960" />
                    <RANKING order="6" place="-1" resultid="6239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9922" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7127" />
                    <RANKING order="2" place="2" resultid="5977" />
                    <RANKING order="3" place="3" resultid="7154" />
                    <RANKING order="4" place="4" resultid="5782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9923" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9924" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9925" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9926" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9518" daytime="15:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9519" daytime="15:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9520" daytime="15:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9521" daytime="15:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9522" daytime="15:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9523" daytime="15:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9524" daytime="15:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9525" daytime="15:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9526" daytime="15:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="9527" daytime="15:54" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="9528" daytime="15:56" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5365" daytime="16:12" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9943" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7066" />
                    <RANKING order="2" place="2" resultid="6627" />
                    <RANKING order="3" place="3" resultid="8319" />
                    <RANKING order="4" place="-1" resultid="8592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9944" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7956" />
                    <RANKING order="2" place="2" resultid="6713" />
                    <RANKING order="3" place="-1" resultid="7107" />
                    <RANKING order="4" place="-1" resultid="7567" />
                    <RANKING order="5" place="-1" resultid="8382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9945" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8325" />
                    <RANKING order="2" place="2" resultid="7202" />
                    <RANKING order="3" place="3" resultid="6150" />
                    <RANKING order="4" place="4" resultid="6778" />
                    <RANKING order="5" place="5" resultid="8343" />
                    <RANKING order="6" place="-1" resultid="7732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9946" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7194" />
                    <RANKING order="2" place="2" resultid="8370" />
                    <RANKING order="3" place="3" resultid="6266" />
                    <RANKING order="4" place="4" resultid="8550" />
                    <RANKING order="5" place="5" resultid="8696" />
                    <RANKING order="6" place="6" resultid="6682" />
                    <RANKING order="7" place="-1" resultid="5972" />
                    <RANKING order="8" place="-1" resultid="8997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9947" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8927" />
                    <RANKING order="2" place="2" resultid="8953" />
                    <RANKING order="3" place="3" resultid="7906" />
                    <RANKING order="4" place="4" resultid="7817" />
                    <RANKING order="5" place="5" resultid="7761" />
                    <RANKING order="6" place="6" resultid="7858" />
                    <RANKING order="7" place="7" resultid="8762" />
                    <RANKING order="8" place="8" resultid="7776" />
                    <RANKING order="9" place="-1" resultid="5808" />
                    <RANKING order="10" place="-1" resultid="6047" />
                    <RANKING order="11" place="-1" resultid="6804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9948" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7697" />
                    <RANKING order="2" place="2" resultid="5747" />
                    <RANKING order="3" place="3" resultid="6663" />
                    <RANKING order="4" place="-1" resultid="6431" />
                    <RANKING order="5" place="-1" resultid="8595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9949" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7385" />
                    <RANKING order="2" place="2" resultid="8844" />
                    <RANKING order="3" place="3" resultid="5989" />
                    <RANKING order="4" place="4" resultid="8016" />
                    <RANKING order="5" place="5" resultid="7864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9950" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6155" />
                    <RANKING order="2" place="2" resultid="6487" />
                    <RANKING order="3" place="3" resultid="7665" />
                    <RANKING order="4" place="4" resultid="6089" />
                    <RANKING order="5" place="5" resultid="6653" />
                    <RANKING order="6" place="6" resultid="6895" />
                    <RANKING order="7" place="7" resultid="6043" />
                    <RANKING order="8" place="8" resultid="8268" />
                    <RANKING order="9" place="-1" resultid="6612" />
                    <RANKING order="10" place="-1" resultid="6834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9951" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8734" />
                    <RANKING order="2" place="2" resultid="6740" />
                    <RANKING order="3" place="3" resultid="8263" />
                    <RANKING order="4" place="4" resultid="6207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9952" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7331" />
                    <RANKING order="2" place="2" resultid="5799" />
                    <RANKING order="3" place="3" resultid="6114" />
                    <RANKING order="4" place="4" resultid="8256" />
                    <RANKING order="5" place="5" resultid="5893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9953" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6194" />
                    <RANKING order="2" place="2" resultid="6877" />
                    <RANKING order="3" place="3" resultid="5698" />
                    <RANKING order="4" place="4" resultid="8251" />
                    <RANKING order="5" place="5" resultid="6413" />
                    <RANKING order="6" place="6" resultid="5712" />
                    <RANKING order="7" place="-1" resultid="6240" />
                    <RANKING order="8" place="-1" resultid="7789" />
                    <RANKING order="9" place="-1" resultid="8636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9954" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8624" />
                    <RANKING order="2" place="2" resultid="5790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9955" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9956" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9957" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9958" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9534" daytime="16:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9535" daytime="16:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9536" daytime="16:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9537" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9538" daytime="16:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9539" daytime="16:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9540" daytime="16:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9541" daytime="16:28" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5348" daytime="15:58" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9927" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6722" />
                    <RANKING order="2" place="2" resultid="8973" />
                    <RANKING order="3" place="3" resultid="5827" />
                    <RANKING order="4" place="4" resultid="6107" />
                    <RANKING order="5" place="-1" resultid="7118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9928" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6160" />
                    <RANKING order="2" place="2" resultid="8537" />
                    <RANKING order="3" place="3" resultid="7045" />
                    <RANKING order="4" place="-1" resultid="6771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9929" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6391" />
                    <RANKING order="2" place="2" resultid="7189" />
                    <RANKING order="3" place="3" resultid="6764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9930" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8568" />
                    <RANKING order="2" place="2" resultid="8771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9931" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7889" />
                    <RANKING order="2" place="2" resultid="7222" />
                    <RANKING order="3" place="3" resultid="7844" />
                    <RANKING order="4" place="4" resultid="8790" />
                    <RANKING order="5" place="-1" resultid="6705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9932" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6233" />
                    <RANKING order="2" place="2" resultid="8356" />
                    <RANKING order="3" place="3" resultid="6673" />
                    <RANKING order="4" place="4" resultid="8668" />
                    <RANKING order="5" place="-1" resultid="6439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9933" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6423" />
                    <RANKING order="2" place="2" resultid="6733" />
                    <RANKING order="3" place="3" resultid="8864" />
                    <RANKING order="4" place="-1" resultid="7530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9934" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6339" />
                    <RANKING order="2" place="2" resultid="6274" />
                    <RANKING order="3" place="3" resultid="6317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9935" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6816" />
                    <RANKING order="2" place="2" resultid="6504" />
                    <RANKING order="3" place="3" resultid="5887" />
                    <RANKING order="4" place="4" resultid="8675" />
                    <RANKING order="5" place="5" resultid="8913" />
                    <RANKING order="6" place="6" resultid="7078" />
                    <RANKING order="7" place="-1" resultid="6727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9936" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9937" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="9938" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6923" />
                    <RANKING order="2" place="-1" resultid="8009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9939" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="9940" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="9941" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="9942" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9529" daytime="15:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9530" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9531" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9532" daytime="16:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9533" daytime="16:08" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-06-24" daytime="09:00" endtime="12:47" number="4">
          <EVENTS>
            <EVENT eventid="5517" daytime="09:08" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10039" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7962" />
                    <RANKING order="2" place="2" resultid="7551" />
                    <RANKING order="3" place="3" resultid="8892" />
                    <RANKING order="4" place="4" resultid="7706" />
                    <RANKING order="5" place="5" resultid="8741" />
                    <RANKING order="6" place="6" resultid="6628" />
                    <RANKING order="7" place="7" resultid="5740" />
                    <RANKING order="8" place="8" resultid="8657" />
                    <RANKING order="9" place="9" resultid="6399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10040" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7957" />
                    <RANKING order="2" place="2" resultid="8747" />
                    <RANKING order="3" place="3" resultid="6714" />
                    <RANKING order="4" place="4" resultid="8942" />
                    <RANKING order="5" place="5" resultid="8719" />
                    <RANKING order="6" place="-1" resultid="7050" />
                    <RANKING order="7" place="-1" resultid="7371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10041" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8335" />
                    <RANKING order="2" place="2" resultid="7897" />
                    <RANKING order="3" place="3" resultid="5863" />
                    <RANKING order="4" place="4" resultid="8362" />
                    <RANKING order="5" place="-1" resultid="8543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10042" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8371" />
                    <RANKING order="2" place="2" resultid="8855" />
                    <RANKING order="3" place="3" resultid="6267" />
                    <RANKING order="4" place="4" resultid="8551" />
                    <RANKING order="5" place="5" resultid="8934" />
                    <RANKING order="6" place="6" resultid="8651" />
                    <RANKING order="7" place="7" resultid="5770" />
                    <RANKING order="8" place="-1" resultid="6249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10043" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8778" />
                    <RANKING order="2" place="2" resultid="7763" />
                    <RANKING order="3" place="3" resultid="8579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10044" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6538" />
                    <RANKING order="2" place="2" resultid="6553" />
                    <RANKING order="3" place="3" resultid="5694" />
                    <RANKING order="4" place="-1" resultid="6374" />
                    <RANKING order="5" place="-1" resultid="6546" />
                    <RANKING order="6" place="-1" resultid="7174" />
                    <RANKING order="7" place="-1" resultid="7433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10045" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6065" />
                    <RANKING order="2" place="2" resultid="7386" />
                    <RANKING order="3" place="3" resultid="7507" />
                    <RANKING order="4" place="4" resultid="7377" />
                    <RANKING order="5" place="-1" resultid="6201" />
                    <RANKING order="6" place="-1" resultid="6648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10046" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6090" />
                    <RANKING order="2" place="2" resultid="6488" />
                    <RANKING order="3" place="3" resultid="6827" />
                    <RANKING order="4" place="4" resultid="8829" />
                    <RANKING order="5" place="-1" resultid="6125" />
                    <RANKING order="6" place="-1" resultid="8300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10047" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8735" />
                    <RANKING order="2" place="2" resultid="8024" />
                    <RANKING order="3" place="3" resultid="7183" />
                    <RANKING order="4" place="4" resultid="6741" />
                    <RANKING order="5" place="5" resultid="5815" />
                    <RANKING order="6" place="6" resultid="6596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10048" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7743" />
                    <RANKING order="2" place="2" resultid="8692" />
                    <RANKING order="3" place="3" resultid="5801" />
                    <RANKING order="4" place="4" resultid="8618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10049" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6080" />
                    <RANKING order="2" place="2" resultid="6463" />
                    <RANKING order="3" place="3" resultid="6415" />
                    <RANKING order="4" place="4" resultid="5687" />
                    <RANKING order="5" place="-1" resultid="6241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10050" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7129" />
                    <RANKING order="2" place="2" resultid="5784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10051" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10052" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10053" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10054" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9572" daytime="09:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9573" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9574" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9575" daytime="09:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9576" daytime="09:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9577" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9578" daytime="09:22" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5602" daytime="10:44" gender="X" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5653" agemax="99" agemin="80" name="Kat. 0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9007" />
                    <RANKING order="2" place="-1" resultid="7597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5654" agemax="119" agemin="100" name="Kat. A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7072" />
                    <RANKING order="2" place="-1" resultid="7595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5655" agemax="159" agemin="120" name="Kat. B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7977" />
                    <RANKING order="2" place="2" resultid="8603" />
                    <RANKING order="3" place="3" resultid="8389" />
                    <RANKING order="4" place="4" resultid="7872" />
                    <RANKING order="5" place="5" resultid="8360" />
                    <RANKING order="6" place="-1" resultid="7978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5656" agemax="199" agemin="160" name="Kat. C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7442" />
                    <RANKING order="2" place="2" resultid="6675" />
                    <RANKING order="3" place="3" resultid="7280" />
                    <RANKING order="4" place="4" resultid="6785" />
                    <RANKING order="5" place="5" resultid="9008" />
                    <RANKING order="6" place="6" resultid="7873" />
                    <RANKING order="7" place="-1" resultid="7510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5657" agemax="239" agemin="200" name="Kat. D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6525" />
                    <RANKING order="2" place="2" resultid="9009" />
                    <RANKING order="3" place="3" resultid="8699" />
                    <RANKING order="4" place="-1" resultid="5980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5658" agemax="279" agemin="240" name="Kat. E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5659" agemax="400" agemin="280" name="Kat. F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6942" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9606" daytime="10:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9607" daytime="10:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9608" daytime="10:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5551" daytime="09:44" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10071" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7067" />
                    <RANKING order="2" place="2" resultid="8859" />
                    <RANKING order="3" place="3" resultid="6629" />
                    <RANKING order="4" place="4" resultid="6398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10072" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5857" />
                    <RANKING order="2" place="2" resultid="6715" />
                    <RANKING order="3" place="3" resultid="7108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10073" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6135" />
                    <RANKING order="2" place="2" resultid="8327" />
                    <RANKING order="3" place="3" resultid="6151" />
                    <RANKING order="4" place="4" resultid="8344" />
                    <RANKING order="5" place="-1" resultid="7734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10074" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7195" />
                    <RANKING order="2" place="2" resultid="6268" />
                    <RANKING order="3" place="3" resultid="8372" />
                    <RANKING order="4" place="4" resultid="8697" />
                    <RANKING order="5" place="5" resultid="6684" />
                    <RANKING order="6" place="6" resultid="8572" />
                    <RANKING order="7" place="-1" resultid="7326" />
                    <RANKING order="8" place="-1" resultid="8998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10075" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8928" />
                    <RANKING order="2" place="2" resultid="8955" />
                    <RANKING order="3" place="3" resultid="6806" />
                    <RANKING order="4" place="4" resultid="8816" />
                    <RANKING order="5" place="5" resultid="7819" />
                    <RANKING order="6" place="6" resultid="7859" />
                    <RANKING order="7" place="7" resultid="8764" />
                    <RANKING order="8" place="8" resultid="7261" />
                    <RANKING order="9" place="9" resultid="7777" />
                    <RANKING order="10" place="10" resultid="8756" />
                    <RANKING order="11" place="-1" resultid="5809" />
                    <RANKING order="12" place="-1" resultid="6049" />
                    <RANKING order="13" place="-1" resultid="7752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10076" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7699" />
                    <RANKING order="2" place="2" resultid="6558" />
                    <RANKING order="3" place="3" resultid="5748" />
                    <RANKING order="4" place="4" resultid="6664" />
                    <RANKING order="5" place="5" resultid="8280" />
                    <RANKING order="6" place="-1" resultid="6432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10077" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7387" />
                    <RANKING order="2" place="2" resultid="8846" />
                    <RANKING order="3" place="3" resultid="5990" />
                    <RANKING order="4" place="4" resultid="8018" />
                    <RANKING order="5" place="5" resultid="7865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10078" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6156" />
                    <RANKING order="2" place="2" resultid="6654" />
                    <RANKING order="3" place="3" resultid="6896" />
                    <RANKING order="4" place="4" resultid="6009" />
                    <RANKING order="5" place="-1" resultid="6045" />
                    <RANKING order="6" place="-1" resultid="6614" />
                    <RANKING order="7" place="-1" resultid="6828" />
                    <RANKING order="8" place="-1" resultid="6836" />
                    <RANKING order="9" place="-1" resultid="8877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10079" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6217" />
                    <RANKING order="2" place="2" resultid="8265" />
                    <RANKING order="3" place="3" resultid="5947" />
                    <RANKING order="4" place="4" resultid="6209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10080" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7333" />
                    <RANKING order="2" place="2" resultid="5802" />
                    <RANKING order="3" place="3" resultid="6116" />
                    <RANKING order="4" place="-1" resultid="5895" />
                    <RANKING order="5" place="-1" resultid="8257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10081" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6195" />
                    <RANKING order="2" place="2" resultid="6878" />
                    <RANKING order="3" place="3" resultid="5699" />
                    <RANKING order="4" place="4" resultid="8252" />
                    <RANKING order="5" place="5" resultid="6416" />
                    <RANKING order="6" place="6" resultid="5713" />
                    <RANKING order="7" place="-1" resultid="7719" />
                    <RANKING order="8" place="-1" resultid="7790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10082" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7155" />
                    <RANKING order="2" place="2" resultid="7130" />
                    <RANKING order="3" place="3" resultid="5785" />
                    <RANKING order="4" place="4" resultid="8626" />
                    <RANKING order="5" place="5" resultid="5792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10083" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10084" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10085" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10086" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9583" daytime="09:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9584" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9585" daytime="09:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9586" daytime="10:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9587" daytime="10:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9588" daytime="10:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9589" daytime="10:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9590" daytime="10:16" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5499" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10023" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10024" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10025" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7338" />
                    <RANKING order="2" place="2" resultid="6392" />
                    <RANKING order="3" place="3" resultid="6028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10026" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7312" />
                    <RANKING order="2" place="2" resultid="6581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10027" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7232" />
                    <RANKING order="2" place="2" resultid="6379" />
                    <RANKING order="3" place="3" resultid="7277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10028" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6234" />
                    <RANKING order="2" place="2" resultid="6440" />
                    <RANKING order="3" place="3" resultid="6445" />
                    <RANKING order="4" place="4" resultid="6497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10029" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6520" />
                    <RANKING order="2" place="2" resultid="7526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10030" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6275" />
                    <RANKING order="2" place="2" resultid="6454" />
                    <RANKING order="3" place="3" resultid="8906" />
                    <RANKING order="4" place="4" resultid="6481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10031" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6506" />
                    <RANKING order="2" place="2" resultid="5966" />
                    <RANKING order="3" place="3" resultid="5888" />
                    <RANKING order="4" place="4" resultid="5916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10032" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="10033" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="10034" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10035" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10036" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10037" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10038" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9569" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9570" daytime="09:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9571" daytime="09:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5534" daytime="09:24" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10055" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6723" />
                    <RANKING order="2" place="2" resultid="8898" />
                    <RANKING order="3" place="-1" resultid="5829" />
                    <RANKING order="4" place="-1" resultid="7119" />
                    <RANKING order="5" place="-1" resultid="8974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10056" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10057" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6393" />
                    <RANKING order="2" place="2" resultid="7191" />
                    <RANKING order="3" place="3" resultid="6766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10058" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8570" />
                    <RANKING order="2" place="-1" resultid="7970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10059" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7224" />
                    <RANKING order="2" place="2" resultid="7890" />
                    <RANKING order="3" place="3" resultid="7845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10060" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8358" />
                    <RANKING order="2" place="2" resultid="6674" />
                    <RANKING order="3" place="3" resultid="8669" />
                    <RANKING order="4" place="4" resultid="6446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10061" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6847" />
                    <RANKING order="2" place="2" resultid="8727" />
                    <RANKING order="3" place="3" resultid="8866" />
                    <RANKING order="4" place="-1" resultid="7531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10062" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6341" />
                    <RANKING order="2" place="2" resultid="7852" />
                    <RANKING order="3" place="3" resultid="5957" />
                    <RANKING order="4" place="-1" resultid="6319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10063" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6818" />
                    <RANKING order="2" place="2" resultid="5889" />
                    <RANKING order="3" place="3" resultid="8676" />
                    <RANKING order="4" place="4" resultid="7079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10064" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8288" />
                    <RANKING order="2" place="-1" resultid="6904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10065" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="10066" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6924" />
                    <RANKING order="2" place="-1" resultid="8010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10067" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10068" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10069" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10070" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9579" daytime="09:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9580" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9581" daytime="09:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9582" daytime="09:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5619" daytime="10:56" gender="F" number="39" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10119" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6568" />
                    <RANKING order="2" place="2" resultid="5830" />
                    <RANKING order="3" place="3" resultid="7684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10120" agemax="29" agemin="25" name="Kat. A" />
                <AGEGROUP agegroupid="10121" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7339" />
                    <RANKING order="2" place="2" resultid="6644" />
                    <RANKING order="3" place="3" resultid="6767" />
                    <RANKING order="4" place="4" resultid="6753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10122" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6313" />
                    <RANKING order="2" place="2" resultid="7489" />
                    <RANKING order="3" place="3" resultid="8352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10123" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6172" />
                    <RANKING order="2" place="2" resultid="7225" />
                    <RANKING order="3" place="3" resultid="6385" />
                    <RANKING order="4" place="4" resultid="7621" />
                    <RANKING order="5" place="5" resultid="7812" />
                    <RANKING order="6" place="6" resultid="8987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10124" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6931" />
                    <RANKING order="2" place="2" resultid="7216" />
                    <RANKING order="3" place="3" resultid="8359" />
                    <RANKING order="4" place="4" resultid="8670" />
                    <RANKING order="5" place="5" resultid="6021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10125" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6848" />
                    <RANKING order="2" place="2" resultid="8728" />
                    <RANKING order="3" place="3" resultid="7637" />
                    <RANKING order="4" place="4" resultid="7359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10126" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7631" />
                    <RANKING order="2" place="2" resultid="6455" />
                    <RANKING order="3" place="3" resultid="6342" />
                    <RANKING order="4" place="4" resultid="7853" />
                    <RANKING order="5" place="5" resultid="6320" />
                    <RANKING order="6" place="6" resultid="6482" />
                    <RANKING order="7" place="-1" resultid="6638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10127" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6819" />
                    <RANKING order="2" place="2" resultid="6507" />
                    <RANKING order="3" place="3" resultid="5917" />
                    <RANKING order="4" place="4" resultid="8915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10128" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8289" />
                    <RANKING order="2" place="2" resultid="6188" />
                    <RANKING order="3" place="3" resultid="7399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10129" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="10130" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="10131" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10132" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10133" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10134" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9609" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9610" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9611" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9612" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5636" daytime="11:02" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10135" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6860" />
                    <RANKING order="2" place="2" resultid="5840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10136" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8644" />
                    <RANKING order="2" place="2" resultid="7041" />
                    <RANKING order="3" place="3" resultid="8748" />
                    <RANKING order="4" place="4" resultid="8555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10137" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6136" />
                    <RANKING order="2" place="2" resultid="7898" />
                    <RANKING order="3" place="3" resultid="8664" />
                    <RANKING order="4" place="4" resultid="8588" />
                    <RANKING order="5" place="-1" resultid="5821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10138" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8856" />
                    <RANKING order="2" place="2" resultid="7302" />
                    <RANKING order="3" place="3" resultid="5771" />
                    <RANKING order="4" place="4" resultid="7835" />
                    <RANKING order="5" place="5" resultid="8935" />
                    <RANKING order="6" place="6" resultid="5973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10139" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8779" />
                    <RANKING order="2" place="2" resultid="8956" />
                    <RANKING order="3" place="3" resultid="8817" />
                    <RANKING order="4" place="4" resultid="7416" />
                    <RANKING order="5" place="5" resultid="5996" />
                    <RANKING order="6" place="6" resultid="7439" />
                    <RANKING order="7" place="7" resultid="7827" />
                    <RANKING order="8" place="8" resultid="7820" />
                    <RANKING order="9" place="9" resultid="7262" />
                    <RANKING order="10" place="10" resultid="7902" />
                    <RANKING order="11" place="11" resultid="6692" />
                    <RANKING order="12" place="12" resultid="8757" />
                    <RANKING order="13" place="13" resultid="8559" />
                    <RANKING order="14" place="-1" resultid="7914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10140" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6539" />
                    <RANKING order="2" place="2" resultid="6873" />
                    <RANKING order="3" place="3" resultid="6554" />
                    <RANKING order="4" place="4" resultid="6547" />
                    <RANKING order="5" place="5" resultid="8281" />
                    <RANKING order="6" place="6" resultid="5732" />
                    <RANKING order="7" place="7" resultid="7347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10141" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6066" />
                    <RANKING order="2" place="2" resultid="6649" />
                    <RANKING order="3" place="3" resultid="7497" />
                    <RANKING order="4" place="4" resultid="8847" />
                    <RANKING order="5" place="5" resultid="7672" />
                    <RANKING order="6" place="6" resultid="8019" />
                    <RANKING order="7" place="7" resultid="5706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10142" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6837" />
                    <RANKING order="2" place="2" resultid="6126" />
                    <RANKING order="3" place="3" resultid="6001" />
                    <RANKING order="4" place="4" resultid="8830" />
                    <RANKING order="5" place="5" resultid="7395" />
                    <RANKING order="6" place="6" resultid="6615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10143" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8736" />
                    <RANKING order="2" place="2" resultid="8709" />
                    <RANKING order="3" place="3" resultid="6326" />
                    <RANKING order="4" place="4" resultid="5722" />
                    <RANKING order="5" place="5" resultid="6182" />
                    <RANKING order="6" place="6" resultid="8967" />
                    <RANKING order="7" place="7" resultid="6015" />
                    <RANKING order="8" place="8" resultid="5948" />
                    <RANKING order="9" place="9" resultid="5816" />
                    <RANKING order="10" place="10" resultid="6210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10144" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7744" />
                    <RANKING order="2" place="2" resultid="8693" />
                    <RANKING order="3" place="3" resultid="6117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10145" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9620" />
                    <RANKING order="2" place="2" resultid="6081" />
                    <RANKING order="3" place="3" resultid="6057" />
                    <RANKING order="4" place="4" resultid="8797" />
                    <RANKING order="5" place="5" resultid="9622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10146" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10147" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="10148" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5941" />
                    <RANKING order="2" place="2" resultid="8435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10149" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10150" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9613" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9614" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9615" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9616" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9617" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9618" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9619" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9621" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5568" daytime="10:20" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10087" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6567" />
                    <RANKING order="2" place="2" resultid="7120" />
                    <RANKING order="3" place="3" resultid="7575" />
                    <RANKING order="4" place="4" resultid="7555" />
                    <RANKING order="5" place="-1" resultid="7650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10088" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6332" />
                    <RANKING order="2" place="2" resultid="5931" />
                    <RANKING order="3" place="3" resultid="7920" />
                    <RANKING order="4" place="4" resultid="7561" />
                    <RANKING order="5" place="5" resultid="8980" />
                    <RANKING order="6" place="6" resultid="8538" />
                    <RANKING order="7" place="7" resultid="6772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10089" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8684" />
                    <RANKING order="2" place="2" resultid="7308" />
                    <RANKING order="3" place="3" resultid="5852" />
                    <RANKING order="4" place="4" resultid="6356" />
                    <RANKING order="5" place="5" resultid="7805" />
                    <RANKING order="6" place="-1" resultid="8378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10090" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7313" />
                    <RANKING order="2" place="2" resultid="7405" />
                    <RANKING order="3" place="3" resultid="8351" />
                    <RANKING order="4" place="4" resultid="7488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10091" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7522" />
                    <RANKING order="2" place="2" resultid="7278" />
                    <RANKING order="3" place="3" resultid="7233" />
                    <RANKING order="4" place="4" resultid="7811" />
                    <RANKING order="5" place="5" resultid="8840" />
                    <RANKING order="6" place="6" resultid="8986" />
                    <RANKING order="7" place="-1" resultid="7643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10092" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6930" />
                    <RANKING order="2" place="2" resultid="7215" />
                    <RANKING order="3" place="3" resultid="6498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10093" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6167" />
                    <RANKING order="2" place="2" resultid="6424" />
                    <RANKING order="3" place="3" resultid="7358" />
                    <RANKING order="4" place="4" resultid="6670" />
                    <RANKING order="5" place="-1" resultid="6521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10094" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6223" />
                    <RANKING order="2" place="2" resultid="8907" />
                    <RANKING order="3" place="3" resultid="5958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10095" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8835" />
                    <RANKING order="2" place="2" resultid="5967" />
                    <RANKING order="3" place="3" resultid="8914" />
                    <RANKING order="4" place="4" resultid="6899" />
                    <RANKING order="5" place="-1" resultid="6728" />
                    <RANKING order="6" place="-1" resultid="7725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10096" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8884" />
                    <RANKING order="2" place="2" resultid="7161" />
                    <RANKING order="3" place="-1" resultid="5671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10097" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6891" />
                    <RANKING order="2" place="2" resultid="6472" />
                    <RANKING order="3" place="-1" resultid="5983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10098" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10099" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10100" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="10101" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10102" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9591" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9592" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9593" daytime="10:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9594" daytime="10:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9595" daytime="10:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9596" daytime="10:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5585" daytime="10:32" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10103" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5839" />
                    <RANKING order="2" place="2" resultid="6622" />
                    <RANKING order="3" place="3" resultid="5847" />
                    <RANKING order="4" place="4" resultid="7516" />
                    <RANKING order="5" place="5" resultid="5755" />
                    <RANKING order="6" place="6" resultid="5679" />
                    <RANKING order="7" place="7" resultid="7707" />
                    <RANKING order="8" place="8" resultid="6859" />
                    <RANKING order="9" place="9" resultid="5741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10104" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5833" />
                    <RANKING order="2" place="2" resultid="7757" />
                    <RANKING order="3" place="3" resultid="8643" />
                    <RANKING order="4" place="4" resultid="7966" />
                    <RANKING order="5" place="5" resultid="5868" />
                    <RANKING order="6" place="6" resultid="6363" />
                    <RANKING order="7" place="7" resultid="7268" />
                    <RANKING order="8" place="8" resultid="7483" />
                    <RANKING order="9" place="9" resultid="7109" />
                    <RANKING order="10" place="10" resultid="8720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10105" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6032" />
                    <RANKING order="2" place="2" resultid="8663" />
                    <RANKING order="3" place="3" resultid="8336" />
                    <RANKING order="4" place="4" resultid="7540" />
                    <RANKING order="5" place="5" resultid="6779" />
                    <RANKING order="6" place="6" resultid="7203" />
                    <RANKING order="7" place="7" resultid="8363" />
                    <RANKING order="8" place="7" resultid="8544" />
                    <RANKING order="9" place="9" resultid="8345" />
                    <RANKING order="10" place="10" resultid="8587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10106" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8921" />
                    <RANKING order="2" place="2" resultid="6250" />
                    <RANKING order="3" place="3" resultid="7365" />
                    <RANKING order="4" place="4" resultid="8552" />
                    <RANKING order="5" place="5" resultid="7834" />
                    <RANKING order="6" place="6" resultid="6685" />
                    <RANKING order="7" place="7" resultid="7473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10107" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8949" />
                    <RANKING order="2" place="2" resultid="7907" />
                    <RANKING order="3" place="3" resultid="7136" />
                    <RANKING order="4" place="4" resultid="6131" />
                    <RANKING order="5" place="5" resultid="8929" />
                    <RANKING order="6" place="6" resultid="6071" />
                    <RANKING order="7" place="7" resultid="7252" />
                    <RANKING order="8" place="8" resultid="7826" />
                    <RANKING order="9" place="8" resultid="8580" />
                    <RANKING order="10" place="10" resultid="6691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10108" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6659" />
                    <RANKING order="2" place="2" resultid="7244" />
                    <RANKING order="3" place="3" resultid="6433" />
                    <RANKING order="4" place="4" resultid="7346" />
                    <RANKING order="5" place="5" resultid="5731" />
                    <RANKING order="6" place="6" resultid="6600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10109" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6308" />
                    <RANKING order="2" place="2" resultid="7671" />
                    <RANKING order="3" place="3" resultid="8272" />
                    <RANKING order="4" place="4" resultid="7496" />
                    <RANKING order="5" place="5" resultid="7378" />
                    <RANKING order="6" place="6" resultid="6606" />
                    <RANKING order="7" place="7" resultid="5705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10110" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8029" />
                    <RANKING order="2" place="2" resultid="6091" />
                    <RANKING order="3" place="3" resultid="7501" />
                    <RANKING order="4" place="4" resultid="6489" />
                    <RANKING order="5" place="5" resultid="7770" />
                    <RANKING order="6" place="6" resultid="6406" />
                    <RANKING order="7" place="-1" resultid="6046" />
                    <RANKING order="8" place="-1" resultid="6262" />
                    <RANKING order="9" place="-1" resultid="8301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10111" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7184" />
                    <RANKING order="2" place="2" resultid="6325" />
                    <RANKING order="3" place="3" resultid="6742" />
                    <RANKING order="4" place="4" resultid="6181" />
                    <RANKING order="5" place="-1" resultid="8243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10112" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7353" />
                    <RANKING order="2" place="2" resultid="6812" />
                    <RANKING order="3" place="3" resultid="7165" />
                    <RANKING order="4" place="4" resultid="6227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10113" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6196" />
                    <RANKING order="2" place="2" resultid="8637" />
                    <RANKING order="3" place="3" resultid="5714" />
                    <RANKING order="4" place="4" resultid="7147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10114" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6908" />
                    <RANKING order="2" place="2" resultid="7156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10115" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8248" />
                    <RANKING order="2" place="2" resultid="6144" />
                    <RANKING order="3" place="3" resultid="8630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10116" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5908" />
                    <RANKING order="2" place="2" resultid="8434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10117" agemax="94" agemin="90" name="Kat. N" />
                <AGEGROUP agegroupid="10118" agemax="99" agemin="95" name="Kat. O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="9597" daytime="10:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9598" daytime="10:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9599" daytime="10:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9600" daytime="10:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="9601" daytime="10:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="9602" daytime="10:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9603" daytime="10:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="9604" daytime="10:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9605" daytime="10:42" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="3WAT" nation="POL" clubid="7518" name="Akademia Sportów Wodnych 3 WATERS">
          <ATHLETES>
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="7517">
              <RESULTS>
                <RESULT eventid="1527" points="304" reactiontime="+74" swimtime="00:01:16.87" resultid="7519" heatid="9474" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="263" reactiontime="+76" swimtime="00:01:40.04" resultid="7520" heatid="9502" lane="3" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="238" reactiontime="+82" swimtime="00:00:39.38" resultid="7521" heatid="9515" lane="2" entrytime="00:00:38.50" />
                <RESULT eventid="5568" points="312" reactiontime="+82" swimtime="00:00:43.32" resultid="7522" heatid="9594" lane="6" entrytime="00:00:43.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-15" firstname="Krystyna" gender="F" lastname="Noskiewicz-Czarnecka" nation="POL" athleteid="7523">
              <RESULTS>
                <RESULT eventid="1561" points="232" reactiontime="+95" swimtime="00:03:18.02" resultid="7524" heatid="9492" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="150" swimtime="00:02:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="287" reactiontime="+87" swimtime="00:06:43.68" resultid="7525" heatid="9563" lane="8" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:33.97" />
                    <SPLIT distance="150" swimtime="00:02:27.55" />
                    <SPLIT distance="200" swimtime="00:03:21.43" />
                    <SPLIT distance="250" swimtime="00:04:18.83" />
                    <SPLIT distance="300" swimtime="00:05:16.98" />
                    <SPLIT distance="350" swimtime="00:06:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="249" reactiontime="+80" swimtime="00:01:28.09" resultid="7526" heatid="9571" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-20" firstname="Agnieszka" gender="F" lastname="Bernat" nation="POL" athleteid="7527">
              <RESULTS>
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="7528" heatid="9460" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="7529" heatid="9501" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="7530" heatid="9531" lane="2" entrytime="00:01:35.00" />
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="7531" heatid="9581" lane="2" entrytime="00:03:05.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WSB" nation="POL" clubid="7101" name="Akademia WSB">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="7100">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="7102" heatid="9330" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="7103" heatid="9345" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="1476" points="260" reactiontime="+73" swimtime="00:00:37.65" resultid="7104" heatid="9456" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1510" status="DNS" swimtime="00:00:00.00" resultid="7105" heatid="9466" lane="4" entrytime="00:03:00.00" />
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="7106" heatid="9506" lane="3" entrytime="00:01:50.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="7107" heatid="9535" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="5551" points="244" reactiontime="+74" swimtime="00:02:58.98" resultid="7108" heatid="9587" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:01:25.35" />
                    <SPLIT distance="150" swimtime="00:02:12.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="358" reactiontime="+70" swimtime="00:00:36.54" resultid="7109" heatid="9598" lane="0" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AMO" nation="POL" clubid="8436" name="Aquasfera Masters Olsztyn">
          <CONTACT name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="8811">
              <RESULTS>
                <RESULT eventid="1314" points="397" swimtime="00:19:45.04" resultid="8812" heatid="9365" lane="9" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                    <SPLIT distance="200" swimtime="00:02:37.54" />
                    <SPLIT distance="250" swimtime="00:03:18.38" />
                    <SPLIT distance="300" swimtime="00:03:59.67" />
                    <SPLIT distance="350" swimtime="00:04:40.88" />
                    <SPLIT distance="400" swimtime="00:05:21.37" />
                    <SPLIT distance="450" swimtime="00:06:01.21" />
                    <SPLIT distance="500" swimtime="00:06:40.70" />
                    <SPLIT distance="550" swimtime="00:07:20.31" />
                    <SPLIT distance="600" swimtime="00:08:00.06" />
                    <SPLIT distance="650" swimtime="00:08:39.78" />
                    <SPLIT distance="700" swimtime="00:09:18.97" />
                    <SPLIT distance="750" swimtime="00:09:58.88" />
                    <SPLIT distance="800" swimtime="00:10:38.40" />
                    <SPLIT distance="850" swimtime="00:11:18.05" />
                    <SPLIT distance="900" swimtime="00:11:57.42" />
                    <SPLIT distance="950" swimtime="00:12:36.69" />
                    <SPLIT distance="1000" swimtime="00:13:15.93" />
                    <SPLIT distance="1050" swimtime="00:13:55.68" />
                    <SPLIT distance="1100" swimtime="00:14:34.77" />
                    <SPLIT distance="1150" swimtime="00:15:13.96" />
                    <SPLIT distance="1200" swimtime="00:15:53.30" />
                    <SPLIT distance="1250" swimtime="00:16:32.86" />
                    <SPLIT distance="1300" swimtime="00:17:11.77" />
                    <SPLIT distance="1350" swimtime="00:17:50.85" />
                    <SPLIT distance="1400" swimtime="00:18:29.37" />
                    <SPLIT distance="1450" swimtime="00:19:08.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="424" swimtime="00:01:02.42" resultid="8813" heatid="9485" lane="9" entrytime="00:01:04.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="399" swimtime="00:02:18.54" resultid="8814" heatid="9555" lane="6" entrytime="00:02:23.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="343" swimtime="00:05:48.10" resultid="8815" heatid="9567" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:08.31" />
                    <SPLIT distance="200" swimtime="00:02:53.11" />
                    <SPLIT distance="250" swimtime="00:03:43.49" />
                    <SPLIT distance="300" swimtime="00:04:33.45" />
                    <SPLIT distance="350" swimtime="00:05:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="307" reactiontime="+68" swimtime="00:02:45.87" resultid="8816" heatid="9588" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:02:04.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="419" reactiontime="+74" swimtime="00:04:53.88" resultid="8817" heatid="9614" lane="0" entrytime="00:05:04.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:47.53" />
                    <SPLIT distance="200" swimtime="00:02:25.55" />
                    <SPLIT distance="250" swimtime="00:03:03.19" />
                    <SPLIT distance="300" swimtime="00:03:41.25" />
                    <SPLIT distance="350" swimtime="00:04:18.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="8785">
              <RESULTS>
                <RESULT eventid="1133" points="266" reactiontime="+89" swimtime="00:00:36.79" resultid="8786" heatid="9311" lane="2" entrytime="00:00:36.55" />
                <RESULT eventid="1458" points="305" reactiontime="+86" swimtime="00:00:40.19" resultid="8788" heatid="9444" lane="9" entrytime="00:00:40.04" />
                <RESULT eventid="1527" points="213" swimtime="00:01:26.57" resultid="8789" heatid="9472" lane="9" entrytime="00:01:25.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="225" reactiontime="+71" swimtime="00:01:35.44" resultid="8790" heatid="9531" lane="4" entrytime="00:01:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-28" firstname="Maciej" gender="M" lastname="Zembrzuski" nation="POL" athleteid="8742">
              <RESULTS>
                <RESULT eventid="1195" points="590" reactiontime="+82" swimtime="00:00:24.92" resultid="8743" heatid="9332" lane="1" entrytime="00:00:24.45" />
                <RESULT eventid="1544" points="625" reactiontime="+78" swimtime="00:00:54.85" resultid="8744" heatid="9490" lane="2" entrytime="00:00:54.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="671" reactiontime="+86" swimtime="00:00:25.62" resultid="8745" heatid="9528" lane="6" entrytime="00:00:25.36" />
                <RESULT eventid="5399" points="502" reactiontime="+81" swimtime="00:02:08.34" resultid="8746" heatid="9558" lane="3" entrytime="00:02:03.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="584" reactiontime="+80" swimtime="00:00:59.57" resultid="8747" heatid="9578" lane="7" entrytime="00:01:01.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="426" reactiontime="+80" swimtime="00:04:52.46" resultid="8748" heatid="9613" lane="0" entrytime="00:04:41.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:42.07" />
                    <SPLIT distance="200" swimtime="00:02:18.23" />
                    <SPLIT distance="250" swimtime="00:02:55.22" />
                    <SPLIT distance="300" swimtime="00:03:34.34" />
                    <SPLIT distance="350" swimtime="00:04:14.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-09" firstname="Aleksandra" gender="F" lastname="Milewska" nation="POL" athleteid="8804">
              <RESULTS>
                <RESULT eventid="1133" points="395" reactiontime="+88" swimtime="00:00:32.26" resultid="8805" heatid="9313" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1212" points="311" swimtime="00:03:06.09" resultid="8806" heatid="9339" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="150" swimtime="00:02:20.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="285" reactiontime="+84" swimtime="00:03:31.18" resultid="8807" heatid="9458" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:42.96" />
                    <SPLIT distance="150" swimtime="00:02:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="8808" heatid="9474" lane="6" entrytime="00:01:12.00" />
                <RESULT eventid="5314" points="325" reactiontime="+84" swimtime="00:00:35.51" resultid="8809" heatid="9516" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="5382" points="302" swimtime="00:02:48.36" resultid="8810" heatid="9546" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-14" firstname="Paweł" gender="M" lastname="Dąbrowski" nation="POL" athleteid="8758">
              <RESULTS>
                <RESULT eventid="1195" points="333" reactiontime="+93" swimtime="00:00:30.16" resultid="8759" heatid="9323" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1476" points="302" reactiontime="+72" swimtime="00:00:35.81" resultid="8760" heatid="9447" lane="2" />
                <RESULT eventid="1544" points="312" reactiontime="+90" swimtime="00:01:09.12" resultid="8761" heatid="9482" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="275" reactiontime="+73" swimtime="00:01:19.72" resultid="8762" heatid="9534" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="260" swimtime="00:02:39.72" resultid="8763" heatid="9553" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:16.54" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="246" reactiontime="+80" swimtime="00:02:58.58" resultid="8764" heatid="9583" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="8721">
              <RESULTS>
                <RESULT eventid="1133" points="295" reactiontime="+80" swimtime="00:00:35.55" resultid="8722" heatid="9312" lane="0" entrytime="00:00:34.50" />
                <RESULT eventid="1297" points="309" reactiontime="+89" swimtime="00:22:47.83" resultid="8723" heatid="9364" lane="4" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:27.12" />
                    <SPLIT distance="150" swimtime="00:02:13.93" />
                    <SPLIT distance="200" swimtime="00:03:00.95" />
                    <SPLIT distance="250" swimtime="00:03:47.63" />
                    <SPLIT distance="300" swimtime="00:04:34.02" />
                    <SPLIT distance="350" swimtime="00:05:20.53" />
                    <SPLIT distance="400" swimtime="00:06:07.05" />
                    <SPLIT distance="450" swimtime="00:06:53.10" />
                    <SPLIT distance="500" swimtime="00:07:39.23" />
                    <SPLIT distance="550" swimtime="00:08:25.17" />
                    <SPLIT distance="600" swimtime="00:09:10.64" />
                    <SPLIT distance="650" swimtime="00:09:55.77" />
                    <SPLIT distance="700" swimtime="00:10:41.65" />
                    <SPLIT distance="750" swimtime="00:11:27.14" />
                    <SPLIT distance="800" swimtime="00:12:13.07" />
                    <SPLIT distance="850" swimtime="00:12:58.62" />
                    <SPLIT distance="900" swimtime="00:13:44.36" />
                    <SPLIT distance="950" swimtime="00:14:29.65" />
                    <SPLIT distance="1000" swimtime="00:15:15.30" />
                    <SPLIT distance="1050" swimtime="00:16:00.60" />
                    <SPLIT distance="1100" swimtime="00:16:46.03" />
                    <SPLIT distance="1150" swimtime="00:17:31.14" />
                    <SPLIT distance="1200" swimtime="00:18:16.77" />
                    <SPLIT distance="1250" swimtime="00:19:02.34" />
                    <SPLIT distance="1300" swimtime="00:19:47.80" />
                    <SPLIT distance="1350" swimtime="00:20:32.97" />
                    <SPLIT distance="1400" swimtime="00:21:18.79" />
                    <SPLIT distance="1450" swimtime="00:22:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="307" reactiontime="+80" swimtime="00:01:16.64" resultid="8724" heatid="9473" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="320" swimtime="00:02:45.14" resultid="8725" heatid="9544" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="247" reactiontime="+88" swimtime="00:07:04.35" resultid="8726" heatid="9562" lane="4" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:51.91" />
                    <SPLIT distance="150" swimtime="00:02:46.97" />
                    <SPLIT distance="200" swimtime="00:03:42.37" />
                    <SPLIT distance="250" swimtime="00:04:38.55" />
                    <SPLIT distance="300" swimtime="00:05:36.37" />
                    <SPLIT distance="350" swimtime="00:06:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="206" reactiontime="+80" swimtime="00:03:30.00" resultid="8727" heatid="9580" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:01:41.84" />
                    <SPLIT distance="150" swimtime="00:02:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="306" reactiontime="+88" swimtime="00:05:50.86" resultid="8728" heatid="9609" lane="0" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:22.78" />
                    <SPLIT distance="150" swimtime="00:02:07.05" />
                    <SPLIT distance="200" swimtime="00:02:52.39" />
                    <SPLIT distance="250" swimtime="00:03:36.98" />
                    <SPLIT distance="300" swimtime="00:04:22.20" />
                    <SPLIT distance="350" swimtime="00:05:06.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Zdzisław" gender="M" lastname="Choroszewski" nation="POL" athleteid="8791">
              <RESULTS>
                <RESULT eventid="1195" points="122" reactiontime="+101" swimtime="00:00:42.10" resultid="8792" heatid="9318" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1280" points="88" reactiontime="+93" swimtime="00:16:53.47" resultid="8793" heatid="9363" lane="5" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.77" />
                    <SPLIT distance="100" swimtime="00:02:01.76" />
                    <SPLIT distance="150" swimtime="00:03:06.60" />
                    <SPLIT distance="200" swimtime="00:04:11.35" />
                    <SPLIT distance="250" swimtime="00:05:16.81" />
                    <SPLIT distance="300" swimtime="00:06:20.71" />
                    <SPLIT distance="350" swimtime="00:07:27.68" />
                    <SPLIT distance="400" swimtime="00:08:31.37" />
                    <SPLIT distance="450" swimtime="00:09:34.66" />
                    <SPLIT distance="500" swimtime="00:10:37.93" />
                    <SPLIT distance="550" swimtime="00:11:41.52" />
                    <SPLIT distance="600" swimtime="00:12:46.18" />
                    <SPLIT distance="650" swimtime="00:13:49.18" />
                    <SPLIT distance="700" swimtime="00:14:51.03" />
                    <SPLIT distance="750" swimtime="00:15:54.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="56" reactiontime="+96" swimtime="00:01:02.78" resultid="8794" heatid="9447" lane="6" />
                <RESULT eventid="1544" points="84" reactiontime="+86" swimtime="00:01:46.84" resultid="8795" heatid="9477" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="79" reactiontime="+89" swimtime="00:03:56.93" resultid="8796" heatid="9549" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.49" />
                    <SPLIT distance="100" swimtime="00:01:57.13" />
                    <SPLIT distance="150" swimtime="00:03:01.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="78" reactiontime="+94" swimtime="00:08:34.77" resultid="8797" heatid="9619" lane="7" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                    <SPLIT distance="100" swimtime="00:02:04.52" />
                    <SPLIT distance="150" swimtime="00:03:11.95" />
                    <SPLIT distance="200" swimtime="00:04:19.43" />
                    <SPLIT distance="250" swimtime="00:05:24.84" />
                    <SPLIT distance="300" swimtime="00:06:29.55" />
                    <SPLIT distance="350" swimtime="00:07:34.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="8798">
              <RESULTS>
                <RESULT eventid="1229" points="286" reactiontime="+69" swimtime="00:02:52.94" resultid="8799" heatid="9346" lane="4" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:11.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="274" reactiontime="+70" swimtime="00:03:14.93" resultid="8800" heatid="9467" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:21.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="225" reactiontime="+80" swimtime="00:03:03.15" resultid="8801" heatid="9495" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="263" swimtime="00:01:29.06" resultid="8802" heatid="9511" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="287" reactiontime="+78" swimtime="00:00:33.97" resultid="8803" heatid="9525" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-25" firstname="Adam" gender="M" lastname="Matusiak Vel Matuszewski" nation="POL" athleteid="8749">
              <RESULTS>
                <RESULT eventid="1195" points="209" reactiontime="+83" swimtime="00:00:35.22" resultid="8750" heatid="9320" lane="4" entrytime="00:00:35.11" />
                <RESULT eventid="1280" points="215" reactiontime="+90" swimtime="00:12:34.61" resultid="8751" heatid="9361" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:28.52" />
                    <SPLIT distance="150" swimtime="00:02:15.70" />
                    <SPLIT distance="200" swimtime="00:03:03.07" />
                    <SPLIT distance="250" swimtime="00:03:50.59" />
                    <SPLIT distance="300" swimtime="00:04:38.21" />
                    <SPLIT distance="350" swimtime="00:05:25.84" />
                    <SPLIT distance="400" swimtime="00:06:14.60" />
                    <SPLIT distance="450" swimtime="00:07:02.89" />
                    <SPLIT distance="500" swimtime="00:07:51.32" />
                    <SPLIT distance="550" swimtime="00:08:39.36" />
                    <SPLIT distance="600" swimtime="00:09:27.40" />
                    <SPLIT distance="650" swimtime="00:10:15.72" />
                    <SPLIT distance="700" swimtime="00:11:03.71" />
                    <SPLIT distance="750" swimtime="00:11:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="168" reactiontime="+74" swimtime="00:00:43.49" resultid="8752" heatid="9449" lane="4" entrytime="00:00:46.68" />
                <RESULT eventid="1544" points="216" reactiontime="+81" swimtime="00:01:18.16" resultid="8753" heatid="9480" lane="7" entrytime="00:01:20.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="170" reactiontime="+88" swimtime="00:00:40.45" resultid="8754" heatid="9520" lane="8" entrytime="00:00:43.28" />
                <RESULT eventid="5399" points="208" swimtime="00:02:52.02" resultid="8755" heatid="9552" lane="6" entrytime="00:02:48.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="131" reactiontime="+74" swimtime="00:03:40.11" resultid="8756" heatid="9583" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.37" />
                    <SPLIT distance="100" swimtime="00:01:47.05" />
                    <SPLIT distance="150" swimtime="00:02:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="193" swimtime="00:06:20.74" resultid="8757" heatid="9617" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:32.89" />
                    <SPLIT distance="150" swimtime="00:02:22.17" />
                    <SPLIT distance="200" swimtime="00:03:10.45" />
                    <SPLIT distance="250" swimtime="00:03:59.25" />
                    <SPLIT distance="300" swimtime="00:04:47.55" />
                    <SPLIT distance="350" swimtime="00:05:35.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-28" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="8729">
              <RESULTS>
                <RESULT eventid="1195" points="345" reactiontime="+90" swimtime="00:00:29.81" resultid="8730" heatid="9326" lane="0" entrytime="00:00:29.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski 800 i 400 dow" eventid="1280" points="373" reactiontime="+91" swimtime="00:10:27.97" resultid="8731" heatid="9359" lane="8" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:35.37" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:54.54" />
                    <SPLIT distance="350" swimtime="00:04:34.06" />
                    <SPLIT distance="400" swimtime="00:05:13.48" />
                    <SPLIT distance="450" swimtime="00:05:53.25" />
                    <SPLIT distance="500" swimtime="00:06:32.95" />
                    <SPLIT distance="550" swimtime="00:07:12.82" />
                    <SPLIT distance="600" swimtime="00:07:52.32" />
                    <SPLIT distance="650" swimtime="00:08:32.32" />
                    <SPLIT distance="700" swimtime="00:09:11.75" />
                    <SPLIT distance="750" swimtime="00:09:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1476" points="328" reactiontime="+84" swimtime="00:00:34.85" resultid="8732" heatid="9454" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8733" heatid="9495" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="5365" points="295" reactiontime="+84" swimtime="00:01:17.83" resultid="8734" heatid="9538" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5517" points="317" swimtime="00:01:12.99" resultid="8735" heatid="9576" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5636" points="380" reactiontime="+92" swimtime="00:05:03.62" resultid="8736" heatid="9615" lane="4" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:12.85" />
                    <SPLIT distance="150" swimtime="00:01:50.89" />
                    <SPLIT distance="200" swimtime="00:02:29.54" />
                    <SPLIT distance="250" swimtime="00:03:08.61" />
                    <SPLIT distance="300" swimtime="00:03:47.53" />
                    <SPLIT distance="350" swimtime="00:04:26.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="8765">
              <RESULTS>
                <RESULT eventid="1133" points="376" reactiontime="+82" swimtime="00:00:32.78" resultid="8766" heatid="9312" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="1212" points="313" reactiontime="+82" swimtime="00:03:05.64" resultid="8767" heatid="9339" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:29.36" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="302" reactiontime="+80" swimtime="00:00:40.29" resultid="8768" heatid="9444" lane="2" entrytime="00:00:39.50" />
                <RESULT eventid="1527" points="346" reactiontime="+71" swimtime="00:01:13.62" resultid="8769" heatid="9474" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="318" reactiontime="+75" swimtime="00:00:35.76" resultid="8770" heatid="9515" lane="5" entrytime="00:00:36.60" />
                <RESULT eventid="5348" points="276" reactiontime="+77" swimtime="00:01:29.20" resultid="8771" heatid="9532" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="8772">
              <RESULTS>
                <RESULT eventid="1229" points="475" reactiontime="+70" swimtime="00:02:26.10" resultid="8773" heatid="9348" lane="7" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:52.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="490" reactiontime="+77" swimtime="00:09:33.32" resultid="8774" heatid="9359" lane="3" entrytime="00:09:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                    <SPLIT distance="200" swimtime="00:02:18.34" />
                    <SPLIT distance="250" swimtime="00:02:54.45" />
                    <SPLIT distance="300" swimtime="00:03:30.62" />
                    <SPLIT distance="350" swimtime="00:04:07.09" />
                    <SPLIT distance="400" swimtime="00:04:43.49" />
                    <SPLIT distance="450" swimtime="00:05:19.84" />
                    <SPLIT distance="500" swimtime="00:05:56.39" />
                    <SPLIT distance="550" swimtime="00:06:32.85" />
                    <SPLIT distance="600" swimtime="00:07:09.25" />
                    <SPLIT distance="650" swimtime="00:07:45.31" />
                    <SPLIT distance="700" swimtime="00:08:21.75" />
                    <SPLIT distance="750" swimtime="00:08:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="539" swimtime="00:00:57.64" resultid="8775" heatid="9489" lane="9" entrytime="00:00:58.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="524" swimtime="00:02:06.47" resultid="8776" heatid="9558" lane="9" entrytime="00:02:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="150" swimtime="00:01:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="417" swimtime="00:05:26.26" resultid="8777" heatid="9567" lane="6" entrytime="00:05:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:59.47" />
                    <SPLIT distance="200" swimtime="00:02:41.40" />
                    <SPLIT distance="250" swimtime="00:03:27.55" />
                    <SPLIT distance="300" swimtime="00:04:14.03" />
                    <SPLIT distance="350" swimtime="00:04:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="471" swimtime="00:01:04.00" resultid="8778" heatid="9577" lane="1" entrytime="00:01:05.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="505" swimtime="00:04:36.32" resultid="8779" heatid="9613" lane="1" entrytime="00:04:38.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.35" />
                    <SPLIT distance="150" swimtime="00:01:41.63" />
                    <SPLIT distance="200" swimtime="00:02:17.42" />
                    <SPLIT distance="250" swimtime="00:02:53.17" />
                    <SPLIT distance="300" swimtime="00:03:28.92" />
                    <SPLIT distance="350" swimtime="00:04:04.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-18" firstname="Bogdan" gender="M" lastname="Milewski" nation="POL" athleteid="8780">
              <RESULTS>
                <RESULT eventid="1229" points="199" swimtime="00:03:15.04" resultid="8781" heatid="9342" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:02:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="208" reactiontime="+83" swimtime="00:03:33.62" resultid="8782" heatid="9465" lane="8" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="8783" heatid="9509" lane="9" entrytime="00:01:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-10-03" firstname="Bartosz" gender="M" lastname="Wolak" nation="POL" athleteid="8737">
              <RESULTS>
                <RESULT eventid="1544" points="436" reactiontime="+66" swimtime="00:01:01.83" resultid="8738" heatid="9488" lane="4" entrytime="00:00:58.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="428" reactiontime="+78" swimtime="00:00:29.75" resultid="8739" heatid="9526" lane="6" entrytime="00:00:28.90" />
                <RESULT eventid="5399" points="341" reactiontime="+70" swimtime="00:02:25.86" resultid="8740" heatid="9556" lane="5" entrytime="00:02:17.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="407" reactiontime="+70" swimtime="00:01:07.19" resultid="8741" heatid="9577" lane="0" entrytime="00:01:06.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASG" nation="POL" clubid="7131" name="AquaStars Gdynia">
          <CONTACT email="mariuszgolon5@wp.pl" name="Golon Mariusz" phone="609649755" />
          <ATHLETES>
            <ATHLETE birthdate="1978-11-20" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="7132">
              <RESULTS>
                <RESULT eventid="1280" points="241" reactiontime="+84" swimtime="00:12:06.27" resultid="7133" heatid="9360" lane="0" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:57.76" />
                    <SPLIT distance="200" swimtime="00:02:40.98" />
                    <SPLIT distance="250" swimtime="00:03:25.73" />
                    <SPLIT distance="300" swimtime="00:04:10.47" />
                    <SPLIT distance="350" swimtime="00:04:56.53" />
                    <SPLIT distance="400" swimtime="00:05:43.58" />
                    <SPLIT distance="450" swimtime="00:06:31.65" />
                    <SPLIT distance="500" swimtime="00:07:19.60" />
                    <SPLIT distance="550" swimtime="00:08:07.96" />
                    <SPLIT distance="600" swimtime="00:08:56.24" />
                    <SPLIT distance="650" swimtime="00:09:44.41" />
                    <SPLIT distance="700" swimtime="00:10:32.77" />
                    <SPLIT distance="750" swimtime="00:11:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="7134" heatid="9506" lane="5" entrytime="00:01:50.00" />
                <RESULT eventid="5331" points="468" reactiontime="+81" swimtime="00:00:28.88" resultid="7135" heatid="9524" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="5585" points="412" reactiontime="+84" swimtime="00:00:34.85" resultid="7136" heatid="9598" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="409635" nation="AUS" clubid="7737" name="Australia">
          <ATHLETES>
            <ATHLETE birthdate="1952-12-13" firstname="Maciej" gender="M" lastname="Slugocki" nation="POL" athleteid="7736" externalid="409635">
              <RESULTS>
                <RESULT eventid="1229" points="245" reactiontime="+85" swimtime="00:03:02.16" resultid="7738" heatid="9345" lane="0" entrytime="00:03:03.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:27.09" />
                    <SPLIT distance="150" swimtime="00:02:19.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="313" swimtime="00:21:21.58" resultid="7739" heatid="9366" lane="6" entrytime="00:22:10.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:22.68" />
                    <SPLIT distance="150" swimtime="00:02:05.08" />
                    <SPLIT distance="200" swimtime="00:02:48.37" />
                    <SPLIT distance="250" swimtime="00:03:31.32" />
                    <SPLIT distance="300" swimtime="00:04:14.56" />
                    <SPLIT distance="350" swimtime="00:04:57.40" />
                    <SPLIT distance="400" swimtime="00:05:40.46" />
                    <SPLIT distance="450" swimtime="00:06:23.30" />
                    <SPLIT distance="500" swimtime="00:07:06.29" />
                    <SPLIT distance="550" swimtime="00:07:49.07" />
                    <SPLIT distance="600" swimtime="00:08:32.08" />
                    <SPLIT distance="650" swimtime="00:09:14.73" />
                    <SPLIT distance="700" swimtime="00:09:58.22" />
                    <SPLIT distance="750" swimtime="00:10:41.17" />
                    <SPLIT distance="800" swimtime="00:11:24.45" />
                    <SPLIT distance="850" swimtime="00:12:07.54" />
                    <SPLIT distance="900" swimtime="00:12:50.44" />
                    <SPLIT distance="950" swimtime="00:13:33.50" />
                    <SPLIT distance="1000" swimtime="00:14:16.16" />
                    <SPLIT distance="1050" swimtime="00:14:58.92" />
                    <SPLIT distance="1100" swimtime="00:15:42.14" />
                    <SPLIT distance="1150" swimtime="00:16:25.18" />
                    <SPLIT distance="1200" swimtime="00:17:08.17" />
                    <SPLIT distance="1250" swimtime="00:17:50.96" />
                    <SPLIT distance="1300" swimtime="00:18:34.14" />
                    <SPLIT distance="1350" swimtime="00:19:16.89" />
                    <SPLIT distance="1400" swimtime="00:19:59.75" />
                    <SPLIT distance="1450" swimtime="00:20:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="209" reactiontime="+86" swimtime="00:03:33.12" resultid="7740" heatid="9464" lane="8" entrytime="00:03:34.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                    <SPLIT distance="100" swimtime="00:01:42.84" />
                    <SPLIT distance="150" swimtime="00:02:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="266" reactiontime="+95" swimtime="00:02:38.43" resultid="7741" heatid="9553" lane="7" entrytime="00:02:35.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:01:59.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="219" reactiontime="+101" swimtime="00:06:44.20" resultid="7742" heatid="9566" lane="8" entrytime="00:06:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:39.91" />
                    <SPLIT distance="150" swimtime="00:02:32.93" />
                    <SPLIT distance="200" swimtime="00:03:23.85" />
                    <SPLIT distance="250" swimtime="00:04:21.82" />
                    <SPLIT distance="300" swimtime="00:05:19.48" />
                    <SPLIT distance="350" swimtime="00:06:02.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="186" reactiontime="+102" swimtime="00:01:27.25" resultid="7743" heatid="9573" lane="5" entrytime="00:01:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="305" swimtime="00:05:26.68" resultid="7744" heatid="9616" lane="6" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:02.13" />
                    <SPLIT distance="200" swimtime="00:02:44.01" />
                    <SPLIT distance="250" swimtime="00:03:25.36" />
                    <SPLIT distance="300" swimtime="00:04:07.03" />
                    <SPLIT distance="350" swimtime="00:04:48.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="8417" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501370222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" license="100611700315" athleteid="8427">
              <RESULTS>
                <RESULT eventid="1195" points="35" reactiontime="+121" swimtime="00:01:03.71" resultid="8428" heatid="9318" lane="0" entrytime="00:00:58.48" />
                <RESULT eventid="1314" points="27" swimtime="00:48:00.47" resultid="8429" heatid="9368" lane="6" entrytime="00:44:33.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.46" />
                    <SPLIT distance="100" swimtime="00:02:46.39" />
                    <SPLIT distance="150" swimtime="00:04:19.49" />
                    <SPLIT distance="200" swimtime="00:05:51.72" />
                    <SPLIT distance="250" swimtime="00:07:24.55" />
                    <SPLIT distance="300" swimtime="00:08:59.12" />
                    <SPLIT distance="350" swimtime="00:10:33.95" />
                    <SPLIT distance="400" swimtime="00:12:09.62" />
                    <SPLIT distance="450" swimtime="00:13:46.56" />
                    <SPLIT distance="500" swimtime="00:15:20.87" />
                    <SPLIT distance="550" swimtime="00:16:59.27" />
                    <SPLIT distance="600" swimtime="00:18:34.61" />
                    <SPLIT distance="650" swimtime="00:20:13.02" />
                    <SPLIT distance="700" swimtime="00:21:48.35" />
                    <SPLIT distance="750" swimtime="00:23:27.09" />
                    <SPLIT distance="800" swimtime="00:25:02.38" />
                    <SPLIT distance="850" swimtime="00:26:41.98" />
                    <SPLIT distance="900" swimtime="00:28:17.03" />
                    <SPLIT distance="950" swimtime="00:29:57.66" />
                    <SPLIT distance="1000" swimtime="00:31:39.29" />
                    <SPLIT distance="1050" swimtime="00:33:19.42" />
                    <SPLIT distance="1100" swimtime="00:34:57.54" />
                    <SPLIT distance="1150" swimtime="00:36:41.01" />
                    <SPLIT distance="1200" swimtime="00:38:19.28" />
                    <SPLIT distance="1250" swimtime="00:40:00.34" />
                    <SPLIT distance="1300" swimtime="00:41:39.47" />
                    <SPLIT distance="1350" swimtime="00:43:20.07" />
                    <SPLIT distance="1400" swimtime="00:44:57.13" />
                    <SPLIT distance="1450" swimtime="00:46:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="34" reactiontime="+100" swimtime="00:06:30.49" resultid="8430" heatid="9462" lane="3" entrytime="00:05:52.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.33" />
                    <SPLIT distance="100" swimtime="00:03:09.21" />
                    <SPLIT distance="150" swimtime="00:04:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="8431" heatid="9477" lane="6" entrytime="00:02:32.20" />
                <RESULT eventid="5297" points="31" reactiontime="+114" swimtime="00:03:00.01" resultid="8432" heatid="9505" lane="4" entrytime="00:02:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="31" reactiontime="+96" swimtime="00:05:24.68" resultid="8433" heatid="9548" lane="4" entrytime="00:05:15.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.43" />
                    <SPLIT distance="100" swimtime="00:02:42.56" />
                    <SPLIT distance="150" swimtime="00:04:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="38" swimtime="00:01:17.15" resultid="8434" heatid="9597" lane="1" entrytime="00:01:08.57" />
                <RESULT eventid="5636" points="33" reactiontime="+112" swimtime="00:11:24.12" resultid="8435" heatid="9619" lane="0" entrytime="00:10:21.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.93" />
                    <SPLIT distance="100" swimtime="00:02:43.82" />
                    <SPLIT distance="150" swimtime="00:04:12.89" />
                    <SPLIT distance="200" swimtime="00:05:41.40" />
                    <SPLIT distance="250" swimtime="00:07:09.49" />
                    <SPLIT distance="300" swimtime="00:08:38.15" />
                    <SPLIT distance="350" swimtime="00:10:03.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS" nation="POL" clubid="6357" name="AZS KU Uniwersytetu Warszawskiego" shortname="AZS KU Uniwersytetu Warszawski">
          <CONTACT city="Warszawa" email="mbaranowski@fuw.edu.pl" internet="azs@uw.edu.pl" name="Baranowski Marek" phone="602445201" state="MAZ" street="ul. Dobra 56/66, p. 162" zip="00-312" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" athleteid="6358">
              <RESULTS>
                <RESULT eventid="1195" points="487" reactiontime="+71" swimtime="00:00:26.56" resultid="6359" heatid="9330" lane="5" entrytime="00:00:25.80" entrycourse="LCM" />
                <RESULT eventid="1544" points="545" reactiontime="+68" swimtime="00:00:57.40" resultid="6360" heatid="9489" lane="4" entrytime="00:00:56.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="426" swimtime="00:01:15.91" resultid="6361" heatid="9512" lane="6" entrytime="00:01:12.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="495" reactiontime="+67" swimtime="00:02:08.91" resultid="6362" heatid="9558" lane="8" entrytime="00:02:08.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:03.30" />
                    <SPLIT distance="150" swimtime="00:01:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="438" reactiontime="+69" swimtime="00:00:34.16" resultid="6363" heatid="9603" lane="0" entrytime="00:00:34.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-05" firstname="Yauheni" gender="M" lastname="Puzan" nation="POL" athleteid="6364">
              <RESULTS>
                <RESULT eventid="1195" points="571" reactiontime="+68" swimtime="00:00:25.20" resultid="6365" heatid="9331" lane="0" entrytime="00:00:25.50" entrycourse="LCM" />
                <RESULT eventid="1578" points="549" reactiontime="+76" swimtime="00:02:16.11" resultid="6366" heatid="9496" lane="2" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:03.32" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="629" reactiontime="+74" swimtime="00:00:26.17" resultid="6367" heatid="9528" lane="7" entrytime="00:00:25.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS PWSZ R" nation="POL" region="SLA" clubid="7176" name="AZS PWSZ Racibórz">
          <CONTACT city="Racibórz" email="adip45@poczta.onet.pl" name="PIECHULA" state="ŚLĄSK" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="7177">
              <RESULTS>
                <RESULT eventid="1229" points="229" reactiontime="+84" swimtime="00:03:06.07" resultid="7178" heatid="9344" lane="3" entrytime="00:03:10.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:26.50" />
                    <SPLIT distance="150" swimtime="00:02:20.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="238" reactiontime="+78" swimtime="00:03:24.38" resultid="7179" heatid="9464" lane="3" entrytime="00:03:23.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:37.87" />
                    <SPLIT distance="150" swimtime="00:02:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="165" reactiontime="+98" swimtime="00:03:23.03" resultid="7180" heatid="9494" lane="3" entrytime="00:03:13.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="237" reactiontime="+84" swimtime="00:01:32.25" resultid="7181" heatid="9508" lane="4" entrytime="00:01:29.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="207" reactiontime="+95" swimtime="00:06:52.11" resultid="7182" heatid="9566" lane="0" entrytime="00:06:40.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:38.26" />
                    <SPLIT distance="150" swimtime="00:02:33.97" />
                    <SPLIT distance="200" swimtime="00:03:28.32" />
                    <SPLIT distance="250" swimtime="00:04:25.71" />
                    <SPLIT distance="300" swimtime="00:05:21.57" />
                    <SPLIT distance="350" swimtime="00:06:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="173" reactiontime="+82" swimtime="00:01:29.26" resultid="7183" heatid="9574" lane="7" entrytime="00:01:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="277" reactiontime="+91" swimtime="00:00:39.78" resultid="7184" heatid="9600" lane="7" entrytime="00:00:39.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BB" nation="POL" region="PDL" clubid="7745" name="Barracuda Białystok">
          <CONTACT name="Milewski" phone="606365708" />
          <ATHLETES>
            <ATHLETE birthdate="1977-08-19" firstname="Hubert" gender="M" lastname="Milewski" nation="POL" athleteid="7746">
              <RESULTS>
                <RESULT eventid="1229" points="310" reactiontime="+102" swimtime="00:02:48.32" resultid="7747" heatid="9345" lane="2" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:05.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" reactiontime="+115" status="OTL" swimtime="00:22:48.44" resultid="7748" heatid="9366" lane="2" entrytime="00:22:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:02:01.28" />
                    <SPLIT distance="200" swimtime="00:02:44.89" />
                    <SPLIT distance="250" swimtime="00:03:28.81" />
                    <SPLIT distance="300" swimtime="00:04:13.95" />
                    <SPLIT distance="350" swimtime="00:04:59.84" />
                    <SPLIT distance="400" swimtime="00:05:45.94" />
                    <SPLIT distance="450" swimtime="00:06:32.27" />
                    <SPLIT distance="500" swimtime="00:07:18.41" />
                    <SPLIT distance="550" swimtime="00:08:04.57" />
                    <SPLIT distance="600" swimtime="00:08:51.16" />
                    <SPLIT distance="650" swimtime="00:09:37.83" />
                    <SPLIT distance="700" swimtime="00:10:22.83" />
                    <SPLIT distance="750" swimtime="00:11:10.06" />
                    <SPLIT distance="800" swimtime="00:11:55.53" />
                    <SPLIT distance="850" swimtime="00:12:42.70" />
                    <SPLIT distance="900" swimtime="00:13:28.31" />
                    <SPLIT distance="950" swimtime="00:14:15.86" />
                    <SPLIT distance="1000" swimtime="00:15:01.54" />
                    <SPLIT distance="1050" swimtime="00:15:48.73" />
                    <SPLIT distance="1100" swimtime="00:16:35.19" />
                    <SPLIT distance="1150" swimtime="00:17:22.77" />
                    <SPLIT distance="1200" swimtime="00:18:10.02" />
                    <SPLIT distance="1250" swimtime="00:18:57.08" />
                    <SPLIT distance="1300" swimtime="00:19:43.91" />
                    <SPLIT distance="1350" swimtime="00:20:31.31" />
                    <SPLIT distance="1400" swimtime="00:21:18.24" />
                    <SPLIT distance="1450" swimtime="00:22:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="341" reactiontime="+110" swimtime="00:03:01.24" resultid="7749" heatid="9465" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:27.23" />
                    <SPLIT distance="150" swimtime="00:02:14.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="359" reactiontime="+101" swimtime="00:01:20.33" resultid="7750" heatid="9510" lane="0" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="285" reactiontime="+110" swimtime="00:06:10.14" resultid="7751" heatid="9567" lane="8" entrytime="00:05:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:02:14.68" />
                    <SPLIT distance="200" swimtime="00:03:03.31" />
                    <SPLIT distance="250" swimtime="00:03:51.12" />
                    <SPLIT distance="300" swimtime="00:04:40.18" />
                    <SPLIT distance="350" swimtime="00:05:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="7752" heatid="9586" lane="5" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CP" nation="POL" clubid="7604" name="Cityzen Poznań">
          <CONTACT name="Gołembiewski Tadeusz" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="7615">
              <RESULTS>
                <RESULT eventid="1263" points="265" swimtime="00:12:33.83" resultid="7616" heatid="9356" lane="6" entrytime="00:12:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:11.15" />
                    <SPLIT distance="200" swimtime="00:02:57.85" />
                    <SPLIT distance="250" swimtime="00:03:44.54" />
                    <SPLIT distance="300" swimtime="00:04:32.35" />
                    <SPLIT distance="350" swimtime="00:05:20.39" />
                    <SPLIT distance="400" swimtime="00:06:08.65" />
                    <SPLIT distance="450" swimtime="00:06:57.21" />
                    <SPLIT distance="500" swimtime="00:07:46.17" />
                    <SPLIT distance="550" swimtime="00:08:34.87" />
                    <SPLIT distance="600" swimtime="00:09:23.93" />
                    <SPLIT distance="650" swimtime="00:10:12.65" />
                    <SPLIT distance="700" swimtime="00:11:01.05" />
                    <SPLIT distance="750" swimtime="00:11:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="267" reactiontime="+87" swimtime="00:01:20.21" resultid="7617" heatid="9473" lane="8" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="246" swimtime="00:00:38.95" resultid="7618" heatid="9514" lane="5" entrytime="00:00:47.50" entrycourse="LCM" />
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="7619" heatid="9545" lane="8" entrytime="00:02:58.00" entrycourse="LCM" />
                <RESULT eventid="5450" points="246" reactiontime="+98" swimtime="00:07:04.93" resultid="7620" heatid="9562" lane="5" entrytime="00:07:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:39.95" />
                    <SPLIT distance="150" swimtime="00:02:37.72" />
                    <SPLIT distance="200" swimtime="00:03:33.51" />
                    <SPLIT distance="250" swimtime="00:04:32.08" />
                    <SPLIT distance="300" swimtime="00:05:31.59" />
                    <SPLIT distance="350" swimtime="00:06:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="261" reactiontime="+88" swimtime="00:06:09.62" resultid="7621" heatid="9610" lane="8" entrytime="00:06:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:12.07" />
                    <SPLIT distance="200" swimtime="00:02:59.63" />
                    <SPLIT distance="250" swimtime="00:03:47.64" />
                    <SPLIT distance="300" swimtime="00:04:35.40" />
                    <SPLIT distance="350" swimtime="00:05:23.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-30" firstname="Małgorzata" gender="F" lastname="Rabiega" nation="POL" athleteid="7622">
              <RESULTS>
                <RESULT eventid="1527" points="240" reactiontime="+82" swimtime="00:01:23.18" resultid="7623" heatid="9472" lane="2" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="7624" heatid="9500" lane="7" entrytime="00:03:30.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CMUJ" nation="POL" clubid="7052" name="CMUJ Masters Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="7051">
              <RESULTS>
                <RESULT eventid="1229" points="153" swimtime="00:03:33.00" resultid="7053" heatid="9344" lane="0" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:44.38" />
                    <SPLIT distance="150" swimtime="00:02:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="209" swimtime="00:24:26.52" resultid="7054" heatid="9367" lane="4" entrytime="00:24:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                    <SPLIT distance="200" swimtime="00:03:03.42" />
                    <SPLIT distance="250" swimtime="00:03:51.41" />
                    <SPLIT distance="300" swimtime="00:04:40.63" />
                    <SPLIT distance="350" swimtime="00:05:29.24" />
                    <SPLIT distance="400" swimtime="00:06:19.00" />
                    <SPLIT distance="450" swimtime="00:07:08.26" />
                    <SPLIT distance="500" swimtime="00:07:57.53" />
                    <SPLIT distance="550" swimtime="00:08:47.16" />
                    <SPLIT distance="600" swimtime="00:09:36.99" />
                    <SPLIT distance="650" swimtime="00:10:26.91" />
                    <SPLIT distance="700" swimtime="00:11:15.98" />
                    <SPLIT distance="750" swimtime="00:12:05.59" />
                    <SPLIT distance="800" swimtime="00:12:54.80" />
                    <SPLIT distance="850" swimtime="00:13:44.57" />
                    <SPLIT distance="900" swimtime="00:16:14.51" />
                    <SPLIT distance="950" swimtime="00:15:25.02" />
                    <SPLIT distance="1000" swimtime="00:17:53.61" />
                    <SPLIT distance="1050" swimtime="00:17:04.01" />
                    <SPLIT distance="1100" swimtime="00:19:33.06" />
                    <SPLIT distance="1150" swimtime="00:18:43.51" />
                    <SPLIT distance="1200" swimtime="00:21:13.05" />
                    <SPLIT distance="1250" swimtime="00:20:23.06" />
                    <SPLIT distance="1300" swimtime="00:22:53.64" />
                    <SPLIT distance="1350" swimtime="00:22:03.13" />
                    <SPLIT distance="1400" swimtime="00:24:26.55" />
                    <SPLIT distance="1450" swimtime="00:23:42.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="6616" name="CSIR MOS Dąbrowa Górnicza">
          <CONTACT name="Waliczek Mariusz" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="6623">
              <RESULTS>
                <RESULT eventid="1476" points="436" reactiontime="+69" swimtime="00:00:31.69" resultid="6624" heatid="9456" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6625" heatid="9495" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="5331" points="529" reactiontime="+76" swimtime="00:00:27.73" resultid="6626" heatid="9527" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="5365" points="421" reactiontime="+71" swimtime="00:01:09.18" resultid="6627" heatid="9540" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="382" reactiontime="+75" swimtime="00:01:08.61" resultid="6628" heatid="9578" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="351" reactiontime="+70" swimtime="00:02:38.57" resultid="6629" heatid="9590" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:15.75" />
                    <SPLIT distance="150" swimtime="00:01:56.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-01" firstname="Dawid" gender="M" lastname="Nowodworski" nation="POL" license="102711700137" athleteid="6617">
              <RESULTS>
                <RESULT eventid="1195" points="626" reactiontime="+71" swimtime="00:00:24.44" resultid="6618" heatid="9332" lane="5" entrytime="00:00:23.70" />
                <RESULT eventid="1476" points="597" reactiontime="+79" swimtime="00:00:28.54" resultid="6619" heatid="9457" lane="5" entrytime="00:00:27.81" />
                <RESULT eventid="1544" points="644" swimtime="00:00:54.31" resultid="6620" heatid="9490" lane="1" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="676" reactiontime="+68" swimtime="00:00:25.55" resultid="6621" heatid="9528" lane="5" entrytime="00:00:25.00" />
                <RESULT eventid="5585" points="661" reactiontime="+75" swimtime="00:00:29.78" resultid="6622" heatid="9605" lane="5" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DT" nation="POL" clubid="7513" name="DEEMTEAM">
          <ATHLETES>
            <ATHLETE birthdate="1995-01-14" firstname="Mateusz" gender="M" lastname="Szot" nation="POL" athleteid="7512">
              <RESULTS>
                <RESULT eventid="1510" points="498" swimtime="00:02:39.76" resultid="7514" heatid="9468" lane="9" entrytime="00:02:45.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="593" reactiontime="+69" swimtime="00:01:07.98" resultid="7515" heatid="9511" lane="5" entrytime="00:01:15.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="624" reactiontime="+74" swimtime="00:00:30.36" resultid="7516" heatid="9604" lane="3" entrytime="00:00:32.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="D92" nation="POL" clubid="5707" name="Delfin 92 Gliwice">
          <CONTACT email="cupialsport@op.pl" name="Cupiał Jarosław" phone="605065587" />
          <ATHLETES>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="5708">
              <RESULTS>
                <RESULT eventid="1476" points="52" reactiontime="+122" swimtime="00:01:04.12" resultid="5709" heatid="9448" lane="8" entrytime="00:01:03.80" />
                <RESULT eventid="1510" points="56" reactiontime="+101" swimtime="00:05:30.81" resultid="5710" heatid="9462" lane="5" entrytime="00:05:21.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.76" />
                    <SPLIT distance="100" swimtime="00:02:38.29" />
                    <SPLIT distance="150" swimtime="00:04:07.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="59" swimtime="00:02:26.71" resultid="5711" heatid="9506" lane="9" entrytime="00:02:22.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="47" reactiontime="+106" swimtime="00:02:22.92" resultid="5712" heatid="9534" lane="4" entrytime="00:02:23.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="37" reactiontime="+79" swimtime="00:05:33.60" resultid="5713" heatid="9583" lane="5" entrytime="00:05:48.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.88" />
                    <SPLIT distance="100" swimtime="00:02:42.44" />
                    <SPLIT distance="150" swimtime="00:04:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="78" reactiontime="+131" swimtime="00:01:00.65" resultid="5714" heatid="9597" lane="7" entrytime="00:01:03.98" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DD" nation="POL" clubid="5690" name="Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Wawrzyniec" gender="M" lastname="Mańczak" nation="POL" athleteid="5695">
              <RESULTS>
                <RESULT eventid="1195" points="194" reactiontime="+102" swimtime="00:00:36.09" resultid="5696" heatid="9320" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1476" points="185" reactiontime="+91" swimtime="00:00:42.14" resultid="5697" heatid="9450" lane="6" entrytime="00:00:44.50" />
                <RESULT eventid="5365" points="141" reactiontime="+86" swimtime="00:01:39.55" resultid="5698" heatid="9535" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="117" reactiontime="+105" swimtime="00:03:48.37" resultid="5699" heatid="9585" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:50.58" />
                    <SPLIT distance="150" swimtime="00:02:51.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" athleteid="5689">
              <RESULTS>
                <RESULT eventid="1578" points="236" swimtime="00:03:00.29" resultid="5691" heatid="9495" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="398" reactiontime="+81" swimtime="00:00:30.47" resultid="5692" heatid="9525" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="5399" points="328" reactiontime="+77" swimtime="00:02:27.83" resultid="5693" heatid="9554" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="318" reactiontime="+79" swimtime="00:01:12.93" resultid="5694" heatid="9576" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="381" reactiontime="+76" swimtime="00:00:28.84" resultid="6400" heatid="9325" lane="6" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HUN" nation="HUN" clubid="8712" name="Dr. Regele Károly Szenior Úszóklub">
          <ATHLETES>
            <ATHLETE birthdate="1989-02-05" firstname="Ferenc" gender="M" lastname="Bagdi" nation="HUN" athleteid="8711">
              <RESULTS>
                <RESULT eventid="1280" points="299" reactiontime="+96" swimtime="00:11:16.08" resultid="8713" heatid="9360" lane="3" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:54.80" />
                    <SPLIT distance="200" swimtime="00:02:37.29" />
                    <SPLIT distance="250" swimtime="00:03:20.72" />
                    <SPLIT distance="300" swimtime="00:04:03.85" />
                    <SPLIT distance="350" swimtime="00:04:47.85" />
                    <SPLIT distance="400" swimtime="00:05:31.91" />
                    <SPLIT distance="450" swimtime="00:06:15.80" />
                    <SPLIT distance="500" swimtime="00:06:58.90" />
                    <SPLIT distance="550" swimtime="00:07:42.14" />
                    <SPLIT distance="600" swimtime="00:08:25.36" />
                    <SPLIT distance="650" swimtime="00:09:08.92" />
                    <SPLIT distance="700" swimtime="00:09:52.35" />
                    <SPLIT distance="750" swimtime="00:10:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1229" points="344" swimtime="00:02:42.61" resultid="8714" heatid="9347" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:02:03.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="327" reactiontime="+87" swimtime="00:03:03.69" resultid="8715" heatid="9466" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:26.05" />
                    <SPLIT distance="150" swimtime="00:02:15.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="394" swimtime="00:01:03.97" resultid="8716" heatid="9484" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="385" reactiontime="+94" swimtime="00:00:30.82" resultid="8717" heatid="9524" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="5399" points="355" reactiontime="+84" swimtime="00:02:23.92" resultid="8718" heatid="9555" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="376" swimtime="00:01:08.99" resultid="8719" heatid="9576" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="322" reactiontime="+98" swimtime="00:00:37.85" resultid="8720" heatid="9601" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GM" nation="POL" clubid="7141" name="Gdynia Masters">
          <CONTACT email="kasiiamysiak@gdynia.pl" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="7148">
              <RESULTS>
                <RESULT eventid="1195" points="124" reactiontime="+109" swimtime="00:00:41.84" resultid="7149" heatid="9319" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1229" points="86" swimtime="00:04:17.58" resultid="7150" heatid="9343" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.96" />
                    <SPLIT distance="100" swimtime="00:02:14.78" />
                    <SPLIT distance="150" swimtime="00:03:24.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="95" reactiontime="+99" swimtime="00:00:52.55" resultid="7151" heatid="9449" lane="3" entrytime="00:00:49.50" />
                <RESULT eventid="1544" points="96" reactiontime="+105" swimtime="00:01:42.38" resultid="7152" heatid="9478" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="103" swimtime="00:02:01.52" resultid="7153" heatid="9507" lane="9" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="51" reactiontime="+114" swimtime="00:01:00.33" resultid="7154" heatid="9519" lane="7" entrytime="00:00:49.50" />
                <RESULT eventid="5551" points="62" reactiontime="+91" swimtime="00:04:42.56" resultid="7155" heatid="9584" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.56" />
                    <SPLIT distance="100" swimtime="00:02:17.25" />
                    <SPLIT distance="150" swimtime="00:03:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="134" reactiontime="+116" swimtime="00:00:50.65" resultid="7156" heatid="9598" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="7157">
              <RESULTS>
                <RESULT eventid="1133" points="162" reactiontime="+87" swimtime="00:00:43.41" resultid="7158" heatid="9310" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="1458" points="113" reactiontime="+80" swimtime="00:00:55.88" resultid="7159" heatid="9441" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="5348" points="104" reactiontime="+81" swimtime="00:02:03.25" resultid="7160" heatid="9530" lane="5" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="119" reactiontime="+97" swimtime="00:00:59.70" resultid="7161" heatid="9592" lane="2" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Jan" gender="M" lastname="Boboli" nation="POL" athleteid="7142">
              <RESULTS>
                <RESULT eventid="1195" points="148" reactiontime="+94" swimtime="00:00:39.50" resultid="7143" heatid="9320" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1476" points="52" reactiontime="+87" swimtime="00:01:04.01" resultid="7144" heatid="9448" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="1544" points="112" swimtime="00:01:37.25" resultid="7145" heatid="9479" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="79" reactiontime="+100" swimtime="00:00:52.10" resultid="7146" heatid="9520" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="5585" points="47" reactiontime="+108" swimtime="00:01:11.90" resultid="7147" heatid="9597" lane="3" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="7162">
              <RESULTS>
                <RESULT eventid="1510" points="228" reactiontime="+98" swimtime="00:03:27.16" resultid="7163" heatid="9464" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="240" swimtime="00:01:31.86" resultid="7164" heatid="9508" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="248" reactiontime="+102" swimtime="00:00:41.25" resultid="7165" heatid="9599" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKS" nation="POL" clubid="6096" name="IKS Konstancin">
          <CONTACT email="rafal@juchno.com" name="Juchno" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="6097">
              <RESULTS>
                <RESULT eventid="1195" points="389" reactiontime="+73" swimtime="00:00:28.63" resultid="6098" heatid="9328" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1280" points="339" reactiontime="+80" swimtime="00:10:48.13" resultid="6099" heatid="9360" lane="2" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                    <SPLIT distance="200" swimtime="00:02:35.49" />
                    <SPLIT distance="250" swimtime="00:03:16.78" />
                    <SPLIT distance="300" swimtime="00:03:58.36" />
                    <SPLIT distance="350" swimtime="00:04:40.12" />
                    <SPLIT distance="400" swimtime="00:05:22.04" />
                    <SPLIT distance="450" swimtime="00:06:04.19" />
                    <SPLIT distance="500" swimtime="00:06:45.66" />
                    <SPLIT distance="550" swimtime="00:07:27.32" />
                    <SPLIT distance="600" swimtime="00:08:09.22" />
                    <SPLIT distance="650" swimtime="00:08:50.57" />
                    <SPLIT distance="700" swimtime="00:09:31.98" />
                    <SPLIT distance="750" swimtime="00:10:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="440" reactiontime="+70" swimtime="00:01:01.64" resultid="6100" heatid="9487" lane="0" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="185" reactiontime="+81" swimtime="00:03:15.57" resultid="6101" heatid="9495" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:30.11" />
                    <SPLIT distance="150" swimtime="00:02:21.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="381" reactiontime="+79" swimtime="00:00:30.92" resultid="6102" heatid="9521" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="5399" points="404" swimtime="00:02:17.97" resultid="6103" heatid="9556" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-02-23" firstname="Maciej" gender="M" lastname="Piłatowicz" nation="POL" license="103714700120" athleteid="7170">
              <RESULTS>
                <RESULT eventid="1314" points="243" reactiontime="+86" swimtime="00:23:15.21" resultid="7171" heatid="9366" lane="8" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:01:27.68" />
                    <SPLIT distance="150" swimtime="00:02:14.88" />
                    <SPLIT distance="200" swimtime="00:03:02.99" />
                    <SPLIT distance="250" swimtime="00:03:50.64" />
                    <SPLIT distance="300" swimtime="00:04:37.21" />
                    <SPLIT distance="350" swimtime="00:05:24.37" />
                    <SPLIT distance="400" swimtime="00:06:11.68" />
                    <SPLIT distance="450" swimtime="00:06:59.05" />
                    <SPLIT distance="500" swimtime="00:07:46.01" />
                    <SPLIT distance="550" swimtime="00:08:32.60" />
                    <SPLIT distance="600" swimtime="00:09:18.89" />
                    <SPLIT distance="650" swimtime="00:10:05.06" />
                    <SPLIT distance="700" swimtime="00:10:51.30" />
                    <SPLIT distance="750" swimtime="00:11:37.68" />
                    <SPLIT distance="800" swimtime="00:12:23.54" />
                    <SPLIT distance="850" swimtime="00:13:10.56" />
                    <SPLIT distance="900" swimtime="00:13:56.64" />
                    <SPLIT distance="950" swimtime="00:14:43.67" />
                    <SPLIT distance="1000" swimtime="00:15:30.87" />
                    <SPLIT distance="1050" swimtime="00:16:17.42" />
                    <SPLIT distance="1100" swimtime="00:17:03.99" />
                    <SPLIT distance="1150" swimtime="00:17:50.69" />
                    <SPLIT distance="1200" swimtime="00:18:37.50" />
                    <SPLIT distance="1250" swimtime="00:19:24.33" />
                    <SPLIT distance="1300" swimtime="00:20:11.27" />
                    <SPLIT distance="1350" swimtime="00:20:58.49" />
                    <SPLIT distance="1400" swimtime="00:21:45.04" />
                    <SPLIT distance="1450" swimtime="00:22:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="262" reactiontime="+87" swimtime="00:00:35.03" resultid="7172" heatid="9522" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="5399" points="272" swimtime="00:02:37.26" resultid="7173" heatid="9554" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="7174" heatid="9575" lane="8" entrytime="00:01:19.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-03" firstname="Rafal" gender="M" lastname="Juchno" nation="POL" license="103714700087" athleteid="7455">
              <RESULTS>
                <RESULT eventid="1195" points="371" reactiontime="+93" swimtime="00:00:29.10" resultid="7456" heatid="9324" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1544" points="317" swimtime="00:01:08.76" resultid="7457" heatid="9482" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="250" reactiontime="+90" swimtime="00:01:30.58" resultid="7458" heatid="9508" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="231" reactiontime="+108" swimtime="00:00:36.55" resultid="7459" heatid="9521" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="6002" name="K.S.niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="6010">
              <RESULTS>
                <RESULT eventid="1195" points="142" reactiontime="+104" swimtime="00:00:40.06" resultid="6011" heatid="9317" lane="5" />
                <RESULT eventid="1280" points="142" reactiontime="+109" swimtime="00:14:25.09" resultid="6012" heatid="9362" lane="2" entrytime="00:14:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:30.24" />
                    <SPLIT distance="200" swimtime="00:03:25.07" />
                    <SPLIT distance="250" swimtime="00:04:19.71" />
                    <SPLIT distance="300" swimtime="00:05:14.58" />
                    <SPLIT distance="350" swimtime="00:06:09.88" />
                    <SPLIT distance="400" swimtime="00:07:04.40" />
                    <SPLIT distance="450" swimtime="00:07:59.66" />
                    <SPLIT distance="500" swimtime="00:08:54.23" />
                    <SPLIT distance="550" swimtime="00:09:49.88" />
                    <SPLIT distance="600" swimtime="00:10:45.71" />
                    <SPLIT distance="650" swimtime="00:11:42.49" />
                    <SPLIT distance="700" swimtime="00:12:38.47" />
                    <SPLIT distance="750" swimtime="00:13:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="131" reactiontime="+113" swimtime="00:01:32.31" resultid="6013" heatid="9477" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="137" reactiontime="+105" swimtime="00:03:17.86" resultid="6014" heatid="9550" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:37.12" />
                    <SPLIT distance="150" swimtime="00:02:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="139" reactiontime="+103" swimtime="00:07:04.07" resultid="6015" heatid="9618" lane="2" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:38.14" />
                    <SPLIT distance="150" swimtime="00:02:32.29" />
                    <SPLIT distance="200" swimtime="00:03:27.16" />
                    <SPLIT distance="250" swimtime="00:04:22.70" />
                    <SPLIT distance="300" swimtime="00:05:17.93" />
                    <SPLIT distance="350" swimtime="00:06:12.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="6016">
              <RESULTS>
                <RESULT eventid="1133" points="173" reactiontime="+84" swimtime="00:00:42.42" resultid="6017" heatid="9309" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="1212" points="137" swimtime="00:04:04.33" resultid="6018" heatid="9338" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.38" />
                    <SPLIT distance="100" swimtime="00:02:12.02" />
                    <SPLIT distance="150" swimtime="00:03:13.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="190" swimtime="00:04:01.86" resultid="6019" heatid="9459" lane="7" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.30" />
                    <SPLIT distance="100" swimtime="00:01:57.36" />
                    <SPLIT distance="150" swimtime="00:03:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="156" reactiontime="+96" swimtime="00:03:29.51" resultid="6020" heatid="9543" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:40.24" />
                    <SPLIT distance="150" swimtime="00:02:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="152" reactiontime="+95" swimtime="00:07:23.00" resultid="6021" heatid="9612" lane="4" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                    <SPLIT distance="100" swimtime="00:01:41.57" />
                    <SPLIT distance="150" swimtime="00:02:38.76" />
                    <SPLIT distance="200" swimtime="00:03:35.78" />
                    <SPLIT distance="250" swimtime="00:04:33.08" />
                    <SPLIT distance="300" swimtime="00:05:32.01" />
                    <SPLIT distance="350" swimtime="00:06:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="6003">
              <RESULTS>
                <RESULT eventid="1195" points="210" reactiontime="+92" swimtime="00:00:35.13" resultid="6004" heatid="9320" lane="5" entrytime="00:00:35.30" />
                <RESULT eventid="1280" points="198" swimtime="00:12:54.46" resultid="6005" heatid="9361" lane="1" entrytime="00:13:14.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:20.71" />
                    <SPLIT distance="200" swimtime="00:03:11.25" />
                    <SPLIT distance="250" swimtime="00:04:02.11" />
                    <SPLIT distance="300" swimtime="00:04:52.41" />
                    <SPLIT distance="350" swimtime="00:05:42.53" />
                    <SPLIT distance="400" swimtime="00:06:32.10" />
                    <SPLIT distance="450" swimtime="00:07:21.93" />
                    <SPLIT distance="500" swimtime="00:08:11.08" />
                    <SPLIT distance="550" swimtime="00:08:59.77" />
                    <SPLIT distance="600" swimtime="00:09:47.75" />
                    <SPLIT distance="650" swimtime="00:10:36.00" />
                    <SPLIT distance="700" swimtime="00:11:24.23" />
                    <SPLIT distance="750" swimtime="00:12:11.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="205" reactiontime="+100" swimtime="00:01:19.55" resultid="6006" heatid="9480" lane="4" entrytime="00:01:18.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="135" reactiontime="+108" swimtime="00:00:43.67" resultid="6007" heatid="9519" lane="4" entrytime="00:00:44.43" />
                <RESULT eventid="5399" points="187" swimtime="00:02:58.29" resultid="6008" heatid="9552" lane="9" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="150" swimtime="00:02:14.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="180" reactiontime="+71" swimtime="00:03:18.09" resultid="6009" heatid="9586" lane="7" entrytime="00:03:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                    <SPLIT distance="100" swimtime="00:01:37.44" />
                    <SPLIT distance="150" swimtime="00:02:29.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KAUNO" nation="LTU" clubid="6548" name="Kauno Takas">
          <CONTACT city="Kaunas" email="kaunotakas@gmail.com" name="Romaldas Bickauskas" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1972-02-06" firstname="Vedestas" gender="M" lastname="Sefleris" nation="LTU" athleteid="6549">
              <RESULTS>
                <RESULT eventid="1195" points="457" reactiontime="+67" swimtime="00:00:27.14" resultid="6550" heatid="9328" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1578" points="396" reactiontime="+67" swimtime="00:02:31.77" resultid="6551" heatid="9495" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:48.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="491" reactiontime="+70" swimtime="00:00:28.43" resultid="6552" heatid="9526" lane="4" entrytime="00:00:28.12" />
                <RESULT eventid="5517" points="467" reactiontime="+71" swimtime="00:01:04.17" resultid="6553" heatid="9577" lane="4" entrytime="00:01:02.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="445" reactiontime="+75" swimtime="00:04:48.14" resultid="6554" heatid="9615" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:46.02" />
                    <SPLIT distance="200" swimtime="00:02:22.87" />
                    <SPLIT distance="250" swimtime="00:03:00.02" />
                    <SPLIT distance="300" swimtime="00:03:37.17" />
                    <SPLIT distance="350" swimtime="00:04:14.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="Kersevicius" nation="LTU" athleteid="6555">
              <RESULTS>
                <RESULT eventid="1229" points="340" reactiontime="+85" swimtime="00:02:43.28" resultid="6556" heatid="9346" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:02:03.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="399" reactiontime="+86" swimtime="00:00:32.65" resultid="6557" heatid="9455" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="5551" points="383" reactiontime="+86" swimtime="00:02:34.07" resultid="6558" heatid="9589" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KRO" nation="POL" region="PDK" clubid="7726" name="Klub Pływacki Masters Krosno">
          <CONTACT city="Krosno" email="masters@masters.krosoft.pl" internet="masters.krosoft.pl" name="Szydło" phone="531304943" state="PDK" street="Sportowa 8" zip="38-400" />
          <ATHLETES>
            <ATHLETE birthdate="1986-03-13" firstname="Konrad" gender="M" lastname="Szydło" nation="POL" athleteid="7727">
              <RESULTS>
                <RESULT eventid="1195" points="323" reactiontime="+88" swimtime="00:00:30.47" resultid="7728" heatid="9324" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1314" reactiontime="+91" status="OTL" swimtime="00:20:53.49" resultid="7729" heatid="9365" lane="8" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="150" swimtime="00:01:55.71" />
                    <SPLIT distance="200" swimtime="00:02:36.94" />
                    <SPLIT distance="250" swimtime="00:03:18.64" />
                    <SPLIT distance="300" swimtime="00:04:00.67" />
                    <SPLIT distance="350" swimtime="00:04:42.06" />
                    <SPLIT distance="400" swimtime="00:05:23.29" />
                    <SPLIT distance="450" swimtime="00:06:05.26" />
                    <SPLIT distance="500" swimtime="00:06:46.67" />
                    <SPLIT distance="550" swimtime="00:07:28.80" />
                    <SPLIT distance="600" swimtime="00:08:10.68" />
                    <SPLIT distance="650" swimtime="00:08:53.37" />
                    <SPLIT distance="700" swimtime="00:09:34.88" />
                    <SPLIT distance="750" swimtime="00:10:17.37" />
                    <SPLIT distance="800" swimtime="00:10:59.07" />
                    <SPLIT distance="850" swimtime="00:11:41.75" />
                    <SPLIT distance="900" swimtime="00:12:23.94" />
                    <SPLIT distance="950" swimtime="00:13:05.80" />
                    <SPLIT distance="1000" swimtime="00:13:47.84" />
                    <SPLIT distance="1050" swimtime="00:14:30.96" />
                    <SPLIT distance="1100" swimtime="00:15:13.22" />
                    <SPLIT distance="1150" swimtime="00:15:57.01" />
                    <SPLIT distance="1200" swimtime="00:16:40.23" />
                    <SPLIT distance="1250" swimtime="00:17:23.11" />
                    <SPLIT distance="1300" swimtime="00:18:05.61" />
                    <SPLIT distance="1350" swimtime="00:18:48.52" />
                    <SPLIT distance="1400" swimtime="00:19:30.54" />
                    <SPLIT distance="1450" swimtime="00:20:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="270" reactiontime="+73" swimtime="00:00:37.18" resultid="7730" heatid="9452" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="7731" heatid="9483" lane="0" entrytime="00:01:09.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="7732" heatid="9537" lane="3" entrytime="00:01:25.00" />
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="7733" heatid="9554" lane="5" entrytime="00:02:30.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="7734" heatid="9588" lane="9" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKO" nation="POL" region="WAR" clubid="6022" name="Klub Sportowy MAKO">
          <CONTACT email="annadabrowska@ksmako.pl" name="Anna Dąbrowska" phone="601 480 280" />
          <ATHLETES>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="6029">
              <RESULTS>
                <RESULT eventid="1195" points="636" reactiontime="+74" swimtime="00:00:24.31" resultid="6030" heatid="9332" lane="7" entrytime="00:00:24.37" />
                <RESULT eventid="5297" points="631" swimtime="00:01:06.60" resultid="6031" heatid="9513" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5585" points="694" reactiontime="+73" swimtime="00:00:29.31" resultid="6032" heatid="9605" lane="3" entrytime="00:00:29.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Dąbrowska" nation="POL" athleteid="6023">
              <RESULTS>
                <RESULT eventid="1133" points="245" reactiontime="+85" swimtime="00:00:37.82" resultid="6024" heatid="9311" lane="9" entrytime="00:00:38.01" />
                <RESULT eventid="1527" points="221" reactiontime="+93" swimtime="00:01:25.47" resultid="6025" heatid="9472" lane="0" entrytime="00:01:25.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="177" reactiontime="+120" swimtime="00:00:43.43" resultid="6026" heatid="9515" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="5382" points="211" swimtime="00:03:09.67" resultid="6027" heatid="9544" lane="7" entrytime="00:03:09.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                    <SPLIT distance="150" swimtime="00:02:23.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="165" swimtime="00:01:41.03" resultid="6028" heatid="9570" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="8030" name="Klub Sportowy Warta Poznań">
          <CONTACT city="POZNAŃ" email="jacekthiem@gmail.com" name="THIEM JACEK" phone="502 499 565" state="WIE" street="OSIEDE DĘBINA 19 M 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1962-03-22" firstname="Piotr" gender="M" lastname="Burzyński" nation="POL" athleteid="8873">
              <RESULTS>
                <RESULT eventid="1314" status="OTL" swimtime="00:27:35.27" resultid="8874" heatid="9366" lane="9" entrytime="00:24:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:33.88" />
                    <SPLIT distance="150" swimtime="00:02:26.08" />
                    <SPLIT distance="200" swimtime="00:03:18.32" />
                    <SPLIT distance="250" swimtime="00:04:13.52" />
                    <SPLIT distance="300" swimtime="00:05:07.36" />
                    <SPLIT distance="350" swimtime="00:06:01.96" />
                    <SPLIT distance="400" swimtime="00:06:56.13" />
                    <SPLIT distance="450" swimtime="00:07:51.24" />
                    <SPLIT distance="500" swimtime="00:08:46.34" />
                    <SPLIT distance="550" swimtime="00:09:41.80" />
                    <SPLIT distance="600" swimtime="00:10:36.90" />
                    <SPLIT distance="650" swimtime="00:11:32.30" />
                    <SPLIT distance="700" swimtime="00:12:27.57" />
                    <SPLIT distance="750" swimtime="00:13:25.28" />
                    <SPLIT distance="800" swimtime="00:14:20.16" />
                    <SPLIT distance="850" swimtime="00:15:16.23" />
                    <SPLIT distance="900" swimtime="00:16:12.26" />
                    <SPLIT distance="950" swimtime="00:17:09.57" />
                    <SPLIT distance="1000" swimtime="00:18:04.90" />
                    <SPLIT distance="1050" swimtime="00:19:01.79" />
                    <SPLIT distance="1100" swimtime="00:19:57.31" />
                    <SPLIT distance="1150" swimtime="00:20:54.47" />
                    <SPLIT distance="1200" swimtime="00:21:50.29" />
                    <SPLIT distance="1250" swimtime="00:22:47.67" />
                    <SPLIT distance="1300" swimtime="00:23:44.29" />
                    <SPLIT distance="1350" swimtime="00:24:42.91" />
                    <SPLIT distance="1400" swimtime="00:25:39.24" />
                    <SPLIT distance="1450" swimtime="00:26:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="79" swimtime="00:04:18.82" resultid="8875" heatid="9494" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.47" />
                    <SPLIT distance="100" swimtime="00:02:02.22" />
                    <SPLIT distance="150" swimtime="00:03:10.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="8876" heatid="9565" lane="1" entrytime="00:07:45.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="8877" heatid="9585" lane="6" entrytime="00:03:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-17" firstname="Magdalena" gender="F" lastname="Zajączek" nation="POL" license="500115600524" athleteid="8981">
              <RESULTS>
                <RESULT eventid="1133" points="74" swimtime="00:00:56.29" resultid="8982" heatid="9309" lane="8" entrytime="00:00:57.81" />
                <RESULT eventid="1493" points="141" swimtime="00:04:27.06" resultid="8983" heatid="9458" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.93" />
                    <SPLIT distance="100" swimtime="00:02:09.35" />
                    <SPLIT distance="150" swimtime="00:03:18.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="64" swimtime="00:02:08.78" resultid="8984" heatid="9469" lane="4" entrytime="00:02:06.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="128" swimtime="00:02:07.18" resultid="8985" heatid="9501" lane="1" entrytime="00:02:06.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="128" swimtime="00:00:58.25" resultid="8986" heatid="9592" lane="3" entrytime="00:00:57.45" />
                <RESULT eventid="5619" points="83" swimtime="00:09:01.14" resultid="8987" heatid="9612" lane="8" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.33" />
                    <SPLIT distance="100" swimtime="00:02:08.97" />
                    <SPLIT distance="150" swimtime="00:03:19.05" />
                    <SPLIT distance="200" swimtime="00:04:29.99" />
                    <SPLIT distance="250" swimtime="00:05:39.29" />
                    <SPLIT distance="300" swimtime="00:06:48.83" />
                    <SPLIT distance="350" swimtime="00:07:55.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-08" firstname="Tomasz" gender="M" lastname="Śron" nation="POL" athleteid="8957">
              <RESULTS>
                <RESULT eventid="1195" points="473" reactiontime="+63" swimtime="00:00:26.83" resultid="8958" heatid="9329" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1229" points="382" swimtime="00:02:37.07" resultid="8959" heatid="9349" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="448" reactiontime="+62" swimtime="00:00:31.41" resultid="8960" heatid="9457" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1544" points="525" swimtime="00:00:58.13" resultid="8961" heatid="9489" lane="1" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" license="500115600520" athleteid="8879">
              <RESULTS>
                <RESULT eventid="1133" points="135" reactiontime="+107" swimtime="00:00:46.10" resultid="8880" heatid="9309" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1493" points="164" reactiontime="+118" swimtime="00:04:13.99" resultid="8881" heatid="9459" lane="8" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.71" />
                    <SPLIT distance="100" swimtime="00:02:04.01" />
                    <SPLIT distance="150" swimtime="00:03:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="106" reactiontime="+119" swimtime="00:01:49.22" resultid="8882" heatid="9470" lane="5" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="171" reactiontime="+113" swimtime="00:01:55.50" resultid="8883" heatid="9501" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="188" reactiontime="+110" swimtime="00:00:51.31" resultid="8884" heatid="9593" lane="1" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="8995">
              <RESULTS>
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="8996" heatid="9450" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="8997" heatid="9537" lane="9" entrytime="00:01:30.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="8998" heatid="9587" lane="6" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-07-13" firstname="Paulina" gender="F" lastname="Mendowska" nation="POL" athleteid="8894">
              <RESULTS>
                <RESULT eventid="1212" points="511" reactiontime="+68" swimtime="00:02:37.69" resultid="8895" heatid="9340" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="439" reactiontime="+68" swimtime="00:02:40.16" resultid="8896" heatid="9492" lane="4" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                    <SPLIT distance="150" swimtime="00:01:56.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="488" reactiontime="+72" swimtime="00:01:10.46" resultid="8897" heatid="9571" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="441" reactiontime="+74" swimtime="00:02:42.93" resultid="8898" heatid="9582" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:02.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="Kuca" nation="POL" athleteid="8885">
              <RESULTS>
                <RESULT eventid="1195" points="611" reactiontime="+68" swimtime="00:00:24.63" resultid="8886" heatid="9331" lane="4" entrytime="00:00:24.80" />
                <RESULT eventid="1229" points="599" reactiontime="+64" swimtime="00:02:15.22" resultid="8887" heatid="9349" lane="3" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="650" reactiontime="+62" swimtime="00:00:54.13" resultid="8888" heatid="9490" lane="7" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="8889" heatid="9496" lane="5" entrytime="00:02:15.00" />
                <RESULT eventid="5399" points="593" reactiontime="+64" swimtime="00:02:01.37" resultid="8890" heatid="9558" lane="5" entrytime="00:02:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="100" swimtime="00:00:58.52" />
                    <SPLIT distance="150" swimtime="00:01:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="8891" heatid="9568" lane="2" entrytime="00:05:00.00" />
                <RESULT eventid="5517" points="571" swimtime="00:01:00.03" resultid="8892" heatid="9578" lane="6" entrytime="00:00:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="8848">
              <RESULTS>
                <RESULT eventid="1229" points="502" reactiontime="+63" swimtime="00:02:23.40" resultid="8849" heatid="9349" lane="2" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="465" reactiontime="+64" swimtime="00:09:43.51" resultid="8850" heatid="9359" lane="5" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:43.89" />
                    <SPLIT distance="200" swimtime="00:02:20.60" />
                    <SPLIT distance="250" swimtime="00:02:57.52" />
                    <SPLIT distance="300" swimtime="00:03:34.74" />
                    <SPLIT distance="350" swimtime="00:04:12.15" />
                    <SPLIT distance="400" swimtime="00:04:49.83" />
                    <SPLIT distance="450" swimtime="00:05:27.69" />
                    <SPLIT distance="500" swimtime="00:06:05.38" />
                    <SPLIT distance="550" swimtime="00:06:43.39" />
                    <SPLIT distance="600" swimtime="00:07:21.43" />
                    <SPLIT distance="650" swimtime="00:07:59.46" />
                    <SPLIT distance="700" swimtime="00:08:36.96" />
                    <SPLIT distance="750" swimtime="00:09:12.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="456" swimtime="00:02:44.46" resultid="8851" heatid="9468" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="438" reactiontime="+67" swimtime="00:02:26.83" resultid="8852" heatid="9496" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="486" swimtime="00:02:09.73" resultid="8853" heatid="9558" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:03.48" />
                    <SPLIT distance="150" swimtime="00:01:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="485" swimtime="00:05:10.18" resultid="8854" heatid="9568" lane="1" entrytime="00:05:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:50.82" />
                    <SPLIT distance="200" swimtime="00:02:32.60" />
                    <SPLIT distance="250" swimtime="00:03:16.90" />
                    <SPLIT distance="300" swimtime="00:04:01.82" />
                    <SPLIT distance="350" swimtime="00:04:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="469" reactiontime="+68" swimtime="00:01:04.10" resultid="8855" heatid="9577" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="510" reactiontime="+70" swimtime="00:04:35.36" resultid="8856" heatid="9613" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                    <SPLIT distance="200" swimtime="00:02:15.94" />
                    <SPLIT distance="250" swimtime="00:02:51.72" />
                    <SPLIT distance="300" swimtime="00:03:26.97" />
                    <SPLIT distance="350" swimtime="00:04:02.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-08" firstname="Błażej" gender="M" lastname="Wachowski" nation="POL" athleteid="8930">
              <RESULTS>
                <RESULT eventid="1280" points="273" swimtime="00:11:36.26" resultid="8931" heatid="9360" lane="1" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.97" />
                    <SPLIT distance="200" swimtime="00:02:47.01" />
                    <SPLIT distance="250" swimtime="00:03:30.91" />
                    <SPLIT distance="300" swimtime="00:04:15.31" />
                    <SPLIT distance="350" swimtime="00:04:59.96" />
                    <SPLIT distance="400" swimtime="00:05:44.42" />
                    <SPLIT distance="450" swimtime="00:06:28.64" />
                    <SPLIT distance="500" swimtime="00:07:12.81" />
                    <SPLIT distance="550" swimtime="00:07:57.25" />
                    <SPLIT distance="600" swimtime="00:08:41.29" />
                    <SPLIT distance="650" swimtime="00:09:25.57" />
                    <SPLIT distance="700" swimtime="00:10:09.93" />
                    <SPLIT distance="750" swimtime="00:10:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="224" reactiontime="+99" swimtime="00:03:03.40" resultid="8932" heatid="9495" lane="8" entrytime="00:02:59.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:02:13.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="262" reactiontime="+95" swimtime="00:02:39.21" resultid="8933" heatid="9554" lane="4" entrytime="00:02:29.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="224" reactiontime="+91" swimtime="00:01:21.99" resultid="8934" heatid="9574" lane="2" entrytime="00:01:25.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="278" swimtime="00:05:37.05" resultid="8935" heatid="9615" lane="1" entrytime="00:05:19.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                    <SPLIT distance="200" swimtime="00:02:47.97" />
                    <SPLIT distance="250" swimtime="00:03:31.27" />
                    <SPLIT distance="300" swimtime="00:04:14.82" />
                    <SPLIT distance="350" swimtime="00:04:57.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" license="500115600462" athleteid="8899">
              <RESULTS>
                <RESULT eventid="1212" points="148" reactiontime="+85" swimtime="00:03:58.22" resultid="8900" heatid="9338" lane="8" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.76" />
                    <SPLIT distance="100" swimtime="00:01:58.96" />
                    <SPLIT distance="150" swimtime="00:03:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="179" swimtime="00:04:06.76" resultid="8902" heatid="9459" lane="1" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                    <SPLIT distance="100" swimtime="00:01:56.35" />
                    <SPLIT distance="150" swimtime="00:03:01.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" status="DNS" swimtime="00:00:00.00" resultid="8903" heatid="9491" lane="4" entrytime="00:04:25.00" />
                <RESULT eventid="5279" points="209" reactiontime="+82" swimtime="00:01:47.95" resultid="8904" heatid="9501" lane="2" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="154" swimtime="00:08:16.50" resultid="8905" heatid="9562" lane="7" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.36" />
                    <SPLIT distance="100" swimtime="00:02:02.83" />
                    <SPLIT distance="150" swimtime="00:03:08.48" />
                    <SPLIT distance="200" swimtime="00:04:11.14" />
                    <SPLIT distance="250" swimtime="00:05:16.01" />
                    <SPLIT distance="300" swimtime="00:06:19.62" />
                    <SPLIT distance="350" swimtime="00:07:19.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="95" reactiontime="+95" swimtime="00:02:01.46" resultid="8906" heatid="9569" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="251" reactiontime="+88" swimtime="00:00:46.56" resultid="8907" heatid="9593" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1297" points="128" reactiontime="+99" swimtime="00:30:36.10" resultid="9436" heatid="9364" lane="8" late="yes" entrytime="00:32:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:46.30" />
                    <SPLIT distance="150" swimtime="00:02:45.33" />
                    <SPLIT distance="200" swimtime="00:03:46.23" />
                    <SPLIT distance="250" swimtime="00:04:48.86" />
                    <SPLIT distance="300" swimtime="00:05:51.45" />
                    <SPLIT distance="350" swimtime="00:08:58.72" />
                    <SPLIT distance="400" swimtime="00:07:55.96" />
                    <SPLIT distance="450" swimtime="00:11:03.89" />
                    <SPLIT distance="500" swimtime="00:10:01.33" />
                    <SPLIT distance="550" swimtime="00:13:07.14" />
                    <SPLIT distance="600" swimtime="00:12:04.46" />
                    <SPLIT distance="650" swimtime="00:15:10.67" />
                    <SPLIT distance="700" swimtime="00:14:08.46" />
                    <SPLIT distance="750" swimtime="00:17:15.59" />
                    <SPLIT distance="800" swimtime="00:16:13.02" />
                    <SPLIT distance="850" swimtime="00:19:19.38" />
                    <SPLIT distance="900" swimtime="00:18:16.76" />
                    <SPLIT distance="950" swimtime="00:23:26.80" />
                    <SPLIT distance="1000" swimtime="00:20:20.49" />
                    <SPLIT distance="1050" swimtime="00:27:35.85" />
                    <SPLIT distance="1100" swimtime="00:22:25.28" />
                    <SPLIT distance="1200" swimtime="00:24:28.93" />
                    <SPLIT distance="1300" swimtime="00:26:33.44" />
                    <SPLIT distance="1400" swimtime="00:28:37.23" />
                    <SPLIT distance="1450" swimtime="00:29:37.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="8841">
              <RESULTS>
                <RESULT eventid="1280" points="338" reactiontime="+92" swimtime="00:10:49.01" resultid="8842" heatid="9360" lane="4" entrytime="00:10:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:54.63" />
                    <SPLIT distance="200" swimtime="00:02:34.99" />
                    <SPLIT distance="250" swimtime="00:03:15.85" />
                    <SPLIT distance="300" swimtime="00:03:56.90" />
                    <SPLIT distance="350" swimtime="00:04:38.03" />
                    <SPLIT distance="400" swimtime="00:05:19.60" />
                    <SPLIT distance="450" swimtime="00:06:00.88" />
                    <SPLIT distance="500" swimtime="00:06:42.77" />
                    <SPLIT distance="550" swimtime="00:07:24.20" />
                    <SPLIT distance="600" swimtime="00:08:05.99" />
                    <SPLIT distance="650" swimtime="00:08:47.44" />
                    <SPLIT distance="700" swimtime="00:09:29.50" />
                    <SPLIT distance="750" swimtime="00:10:09.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="374" reactiontime="+73" swimtime="00:00:33.34" resultid="8843" heatid="9454" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="5365" points="354" reactiontime="+81" swimtime="00:01:13.29" resultid="8844" heatid="9539" lane="3" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="322" reactiontime="+85" swimtime="00:02:28.67" resultid="8845" heatid="9555" lane="2" entrytime="00:02:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="330" reactiontime="+83" swimtime="00:02:41.83" resultid="8846" heatid="9589" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:00.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="343" swimtime="00:05:14.32" resultid="8847" heatid="9614" lane="9" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.48" />
                    <SPLIT distance="150" swimtime="00:01:52.95" />
                    <SPLIT distance="200" swimtime="00:02:33.60" />
                    <SPLIT distance="250" swimtime="00:03:14.38" />
                    <SPLIT distance="300" swimtime="00:03:56.56" />
                    <SPLIT distance="350" swimtime="00:04:36.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-12" firstname="Włodzimierz" gender="M" lastname="Wiatr" nation="POL" athleteid="8962">
              <RESULTS>
                <RESULT eventid="1229" points="104" reactiontime="+95" swimtime="00:04:01.90" resultid="8963" heatid="9343" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.71" />
                    <SPLIT distance="100" swimtime="00:02:02.70" />
                    <SPLIT distance="150" swimtime="00:03:10.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="142" swimtime="00:14:25.75" resultid="8964" heatid="9362" lane="1" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                    <SPLIT distance="150" swimtime="00:02:36.00" />
                    <SPLIT distance="200" swimtime="00:03:31.16" />
                    <SPLIT distance="250" swimtime="00:04:26.18" />
                    <SPLIT distance="300" swimtime="00:05:21.98" />
                    <SPLIT distance="350" swimtime="00:06:17.47" />
                    <SPLIT distance="400" swimtime="00:07:12.30" />
                    <SPLIT distance="450" swimtime="00:08:07.80" />
                    <SPLIT distance="500" swimtime="00:09:03.20" />
                    <SPLIT distance="550" swimtime="00:09:57.29" />
                    <SPLIT distance="600" swimtime="00:10:53.08" />
                    <SPLIT distance="650" swimtime="00:11:47.03" />
                    <SPLIT distance="700" swimtime="00:12:41.05" />
                    <SPLIT distance="750" swimtime="00:13:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="135" swimtime="00:01:51.14" resultid="8965" heatid="9506" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="122" reactiontime="+94" swimtime="00:03:25.34" resultid="8966" heatid="9550" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:36.82" />
                    <SPLIT distance="150" swimtime="00:02:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="141" reactiontime="+106" swimtime="00:07:02.70" resultid="8967" heatid="9619" lane="4" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                    <SPLIT distance="150" swimtime="00:02:33.41" />
                    <SPLIT distance="200" swimtime="00:03:28.22" />
                    <SPLIT distance="250" swimtime="00:04:21.24" />
                    <SPLIT distance="300" swimtime="00:05:16.29" />
                    <SPLIT distance="350" swimtime="00:06:10.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-01" firstname="Paula" gender="F" lastname="Owczarzak" nation="POL" athleteid="8975">
              <RESULTS>
                <RESULT eventid="1263" points="233" reactiontime="+92" swimtime="00:13:06.87" resultid="8976" heatid="9355" lane="0" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:02:04.36" />
                    <SPLIT distance="200" swimtime="00:02:53.23" />
                    <SPLIT distance="250" swimtime="00:03:44.40" />
                    <SPLIT distance="300" swimtime="00:04:36.38" />
                    <SPLIT distance="350" swimtime="00:05:27.51" />
                    <SPLIT distance="400" swimtime="00:06:18.60" />
                    <SPLIT distance="450" swimtime="00:07:09.65" />
                    <SPLIT distance="500" swimtime="00:08:00.74" />
                    <SPLIT distance="550" swimtime="00:08:52.18" />
                    <SPLIT distance="600" swimtime="00:09:44.88" />
                    <SPLIT distance="650" swimtime="00:10:36.89" />
                    <SPLIT distance="700" swimtime="00:11:27.14" />
                    <SPLIT distance="750" swimtime="00:12:18.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="332" reactiontime="+81" swimtime="00:03:20.87" resultid="8977" heatid="9460" lane="5" entrytime="00:03:15.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:33.07" />
                    <SPLIT distance="150" swimtime="00:02:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="340" reactiontime="+84" swimtime="00:01:31.88" resultid="8978" heatid="9503" lane="2" entrytime="00:01:32.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="287" reactiontime="+83" swimtime="00:02:51.27" resultid="8979" heatid="9546" lane="2" entrytime="00:02:45.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="338" reactiontime="+92" swimtime="00:00:42.19" resultid="8980" heatid="9593" lane="6" entrytime="00:00:47.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="8860">
              <RESULTS>
                <RESULT eventid="1263" points="210" swimtime="00:13:35.19" resultid="8861" heatid="9356" lane="8" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:30.47" />
                    <SPLIT distance="150" swimtime="00:02:19.61" />
                    <SPLIT distance="200" swimtime="00:03:09.74" />
                    <SPLIT distance="250" swimtime="00:04:00.61" />
                    <SPLIT distance="300" swimtime="00:04:52.25" />
                    <SPLIT distance="350" swimtime="00:05:44.53" />
                    <SPLIT distance="400" swimtime="00:06:37.24" />
                    <SPLIT distance="450" swimtime="00:07:28.87" />
                    <SPLIT distance="500" swimtime="00:08:20.67" />
                    <SPLIT distance="550" swimtime="00:09:13.21" />
                    <SPLIT distance="600" swimtime="00:10:06.50" />
                    <SPLIT distance="650" swimtime="00:10:59.16" />
                    <SPLIT distance="700" swimtime="00:11:51.53" />
                    <SPLIT distance="750" swimtime="00:12:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" status="DNS" swimtime="00:00:00.00" resultid="8862" heatid="9442" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="8863" heatid="9471" lane="6" entrytime="00:01:27.00" />
                <RESULT eventid="5348" points="179" reactiontime="+114" swimtime="00:01:42.95" resultid="8864" heatid="9531" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="8865" heatid="9544" lane="4" entrytime="00:03:01.00" />
                <RESULT eventid="5534" points="190" reactiontime="+119" swimtime="00:03:35.73" resultid="8866" heatid="9580" lane="6" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                    <SPLIT distance="100" swimtime="00:01:45.79" />
                    <SPLIT distance="150" swimtime="00:02:41.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-31" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" license="500115700461" athleteid="8943">
              <RESULTS>
                <RESULT eventid="1195" points="448" reactiontime="+81" swimtime="00:00:27.32" resultid="8944" heatid="9328" lane="6" entrytime="00:00:27.27" />
                <RESULT eventid="1510" points="456" reactiontime="+73" swimtime="00:02:44.48" resultid="8945" heatid="9467" lane="4" entrytime="00:02:49.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:02:01.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="8946" heatid="9487" lane="9" entrytime="00:01:01.89" />
                <RESULT eventid="5297" points="477" reactiontime="+78" swimtime="00:01:13.08" resultid="8947" heatid="9512" lane="8" entrytime="00:01:14.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="392" reactiontime="+80" swimtime="00:00:30.63" resultid="8948" heatid="9525" lane="4" entrytime="00:00:29.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5585" points="515" reactiontime="+76" swimtime="00:00:32.36" resultid="8949" heatid="9604" lane="1" entrytime="00:00:32.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-11" firstname="Piotr" gender="M" lastname="Witt" nation="POL" athleteid="8936">
              <RESULTS>
                <RESULT eventid="1195" points="553" reactiontime="+76" swimtime="00:00:25.47" resultid="8937" heatid="9331" lane="7" entrytime="00:00:25.21" />
                <RESULT eventid="1476" points="448" reactiontime="+79" swimtime="00:00:31.41" resultid="8938" heatid="9456" lane="3" entrytime="00:00:30.89" />
                <RESULT eventid="1544" points="565" swimtime="00:00:56.74" resultid="8939" heatid="9489" lane="6" entrytime="00:00:57.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="512" reactiontime="+79" swimtime="00:00:28.02" resultid="8940" heatid="9527" lane="8" entrytime="00:00:27.77" />
                <RESULT eventid="5399" points="476" reactiontime="+74" swimtime="00:02:10.58" resultid="8941" heatid="9557" lane="3" entrytime="00:02:11.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="100" swimtime="00:01:01.74" />
                    <SPLIT distance="150" swimtime="00:01:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="426" reactiontime="+66" swimtime="00:01:06.17" resultid="8942" heatid="9577" lane="2" entrytime="00:01:04.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-01" firstname="Natalia" gender="F" lastname="Wiśniewska" nation="POL" athleteid="8988">
              <RESULTS>
                <RESULT eventid="1133" points="445" reactiontime="+85" swimtime="00:00:30.99" resultid="8989" heatid="9314" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1212" points="466" reactiontime="+80" swimtime="00:02:42.65" resultid="8990" heatid="9340" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:02:02.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="473" reactiontime="+80" swimtime="00:02:58.49" resultid="8991" heatid="9461" lane="3" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:25.11" />
                    <SPLIT distance="150" swimtime="00:02:11.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="404" reactiontime="+76" swimtime="00:01:09.91" resultid="8992" heatid="9475" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="460" swimtime="00:01:23.07" resultid="8993" heatid="9504" lane="6" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="456" reactiontime="+76" swimtime="00:05:45.83" resultid="8994" heatid="9563" lane="5" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:02:02.27" />
                    <SPLIT distance="200" swimtime="00:02:47.63" />
                    <SPLIT distance="250" swimtime="00:03:33.97" />
                    <SPLIT distance="300" swimtime="00:04:22.10" />
                    <SPLIT distance="350" swimtime="00:05:05.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" license="500115600525" athleteid="8836">
              <RESULTS>
                <RESULT eventid="1133" points="71" reactiontime="+101" swimtime="00:00:57.12" resultid="8837" heatid="9309" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1493" points="126" reactiontime="+101" swimtime="00:04:36.99" resultid="8838" heatid="9458" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.86" />
                    <SPLIT distance="100" swimtime="00:02:12.64" />
                    <SPLIT distance="150" swimtime="00:03:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="132" reactiontime="+108" swimtime="00:02:05.82" resultid="8839" heatid="9501" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="134" reactiontime="+101" swimtime="00:00:57.33" resultid="8840" heatid="9592" lane="5" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" license="500115700493" athleteid="8831">
              <RESULTS>
                <RESULT eventid="1133" points="262" reactiontime="+70" swimtime="00:00:36.97" resultid="8832" heatid="9311" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1493" points="293" reactiontime="+87" swimtime="00:03:29.21" resultid="8833" heatid="9460" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:41.50" />
                    <SPLIT distance="150" swimtime="00:02:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="301" swimtime="00:01:35.66" resultid="8834" heatid="9503" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="294" reactiontime="+84" swimtime="00:00:44.21" resultid="8835" heatid="9593" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="8824">
              <RESULTS>
                <RESULT eventid="1280" points="160" reactiontime="+93" swimtime="00:13:51.63" resultid="8825" heatid="9361" lane="0" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:31.40" />
                    <SPLIT distance="150" swimtime="00:02:22.51" />
                    <SPLIT distance="200" swimtime="00:03:12.80" />
                    <SPLIT distance="250" swimtime="00:04:04.21" />
                    <SPLIT distance="300" swimtime="00:04:56.56" />
                    <SPLIT distance="350" swimtime="00:05:48.62" />
                    <SPLIT distance="400" swimtime="00:06:42.20" />
                    <SPLIT distance="450" swimtime="00:07:35.51" />
                    <SPLIT distance="500" swimtime="00:08:29.08" />
                    <SPLIT distance="550" swimtime="00:09:23.16" />
                    <SPLIT distance="600" swimtime="00:10:18.32" />
                    <SPLIT distance="650" swimtime="00:11:12.30" />
                    <SPLIT distance="700" swimtime="00:12:05.88" />
                    <SPLIT distance="750" swimtime="00:13:00.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="173" reactiontime="+96" swimtime="00:03:20.05" resultid="8826" heatid="9494" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="100" swimtime="00:01:35.00" />
                    <SPLIT distance="150" swimtime="00:02:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="193" reactiontime="+96" swimtime="00:00:38.77" resultid="8827" heatid="9520" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="5399" points="181" reactiontime="+91" swimtime="00:03:00.06" resultid="8828" heatid="9552" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="150" swimtime="00:02:16.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="183" reactiontime="+83" swimtime="00:01:27.62" resultid="8829" heatid="9574" lane="0" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="171" reactiontime="+107" swimtime="00:06:36.22" resultid="8830" heatid="9617" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:34.99" />
                    <SPLIT distance="150" swimtime="00:02:26.45" />
                    <SPLIT distance="200" swimtime="00:03:17.90" />
                    <SPLIT distance="250" swimtime="00:04:08.59" />
                    <SPLIT distance="300" swimtime="00:04:59.76" />
                    <SPLIT distance="350" swimtime="00:05:49.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-08" firstname="Katarzyna" gender="F" lastname="Mendowska" nation="POL" athleteid="8968">
              <RESULTS>
                <RESULT eventid="1133" points="495" reactiontime="+81" swimtime="00:00:29.92" resultid="8969" heatid="9314" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1458" points="475" reactiontime="+76" swimtime="00:00:34.66" resultid="8970" heatid="9445" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1527" points="427" reactiontime="+71" swimtime="00:01:08.66" resultid="8971" heatid="9475" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="429" reactiontime="+77" swimtime="00:00:32.38" resultid="8972" heatid="9516" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="5348" points="445" reactiontime="+71" swimtime="00:01:16.09" resultid="8973" heatid="9533" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="8974" heatid="9582" lane="3" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Szymon" gender="M" lastname="Wieja" nation="POL" license="500115700467" athleteid="8922">
              <RESULTS>
                <RESULT eventid="1195" points="445" reactiontime="+79" swimtime="00:00:27.37" resultid="8923" heatid="9322" lane="9" entrytime="00:00:32.99" />
                <RESULT eventid="1229" points="438" swimtime="00:02:30.03" resultid="8924" heatid="9348" lane="1" entrytime="00:02:33.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="432" swimtime="00:00:31.78" resultid="8925" heatid="9455" lane="6" entrytime="00:00:32.13" />
                <RESULT eventid="1544" points="489" reactiontime="+72" swimtime="00:00:59.51" resultid="8926" heatid="9487" lane="4" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="400" reactiontime="+61" swimtime="00:01:10.32" resultid="8927" heatid="9540" lane="2" entrytime="00:01:09.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="376" reactiontime="+71" swimtime="00:02:35.01" resultid="8928" heatid="9589" lane="2" entrytime="00:02:37.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:01:56.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="380" reactiontime="+81" swimtime="00:00:35.80" resultid="8929" heatid="9602" lane="3" entrytime="00:00:35.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="8868">
              <RESULTS>
                <RESULT eventid="1195" points="381" reactiontime="+85" swimtime="00:00:28.82" resultid="8869" heatid="9326" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1544" points="429" reactiontime="+77" swimtime="00:01:02.19" resultid="8870" heatid="9486" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="374" swimtime="00:02:21.52" resultid="8871" heatid="9556" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:46.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-07-11" firstname="Waldemar" gender="M" lastname="Krakowiak" nation="POL" license="100115700335" athleteid="8857">
              <RESULTS>
                <RESULT eventid="1229" points="434" reactiontime="+59" swimtime="00:02:30.57" resultid="8858" heatid="9349" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:50.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="391" reactiontime="+78" swimtime="00:02:32.95" resultid="8859" heatid="9590" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:50.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" license="100115600353" athleteid="8908">
              <RESULTS>
                <RESULT eventid="1263" points="84" reactiontime="+112" swimtime="00:18:26.87" resultid="8909" heatid="9357" lane="2" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                    <SPLIT distance="100" swimtime="00:01:59.43" />
                    <SPLIT distance="150" swimtime="00:03:07.85" />
                    <SPLIT distance="200" swimtime="00:04:19.19" />
                    <SPLIT distance="250" swimtime="00:05:31.07" />
                    <SPLIT distance="300" swimtime="00:06:42.15" />
                    <SPLIT distance="350" swimtime="00:07:54.40" />
                    <SPLIT distance="400" swimtime="00:16:08.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="138" reactiontime="+124" swimtime="00:04:28.61" resultid="8910" heatid="9458" lane="4" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                    <SPLIT distance="100" swimtime="00:02:10.08" />
                    <SPLIT distance="150" swimtime="00:03:20.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="95" reactiontime="+118" swimtime="00:01:53.01" resultid="8911" heatid="9470" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="119" swimtime="00:02:10.31" resultid="8912" heatid="9501" lane="7" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="68" reactiontime="+91" swimtime="00:02:21.89" resultid="8913" heatid="9530" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="132" reactiontime="+109" swimtime="00:00:57.64" resultid="8914" heatid="9592" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="5619" points="83" swimtime="00:09:00.10" resultid="8915" heatid="9612" lane="1" entrytime="00:09:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.24" />
                    <SPLIT distance="100" swimtime="00:02:01.67" />
                    <SPLIT distance="150" swimtime="00:03:10.66" />
                    <SPLIT distance="200" swimtime="00:04:20.50" />
                    <SPLIT distance="250" swimtime="00:05:31.76" />
                    <SPLIT distance="300" swimtime="00:06:42.40" />
                    <SPLIT distance="350" swimtime="00:07:54.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-02" firstname="Daniel" gender="M" lastname="Osik" nation="POL" license="500115700521" athleteid="8950">
              <RESULTS>
                <RESULT eventid="1476" points="375" reactiontime="+72" swimtime="00:00:33.32" resultid="8952" heatid="9455" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="5365" points="380" reactiontime="+77" swimtime="00:01:11.53" resultid="8953" heatid="9540" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="406" swimtime="00:02:17.72" resultid="8954" heatid="9557" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="371" reactiontime="+81" swimtime="00:02:35.63" resultid="8955" heatid="9589" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:17.86" />
                    <SPLIT distance="150" swimtime="00:01:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="444" reactiontime="+86" swimtime="00:04:48.37" resultid="8956" heatid="9613" lane="8" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                    <SPLIT distance="200" swimtime="00:02:21.71" />
                    <SPLIT distance="250" swimtime="00:02:58.48" />
                    <SPLIT distance="300" swimtime="00:03:36.04" />
                    <SPLIT distance="350" swimtime="00:04:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="414" reactiontime="+99" swimtime="00:19:28.30" resultid="9439" heatid="9367" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                    <SPLIT distance="200" swimtime="00:02:26.91" />
                    <SPLIT distance="250" swimtime="00:03:05.25" />
                    <SPLIT distance="300" swimtime="00:03:44.06" />
                    <SPLIT distance="350" swimtime="00:04:23.03" />
                    <SPLIT distance="400" swimtime="00:05:03.09" />
                    <SPLIT distance="450" swimtime="00:05:42.17" />
                    <SPLIT distance="500" swimtime="00:06:21.75" />
                    <SPLIT distance="550" swimtime="00:07:00.96" />
                    <SPLIT distance="600" swimtime="00:07:40.56" />
                    <SPLIT distance="650" swimtime="00:08:19.81" />
                    <SPLIT distance="700" swimtime="00:08:58.99" />
                    <SPLIT distance="750" swimtime="00:09:38.47" />
                    <SPLIT distance="800" swimtime="00:10:18.58" />
                    <SPLIT distance="850" swimtime="00:10:57.63" />
                    <SPLIT distance="900" swimtime="00:11:37.55" />
                    <SPLIT distance="950" swimtime="00:12:17.28" />
                    <SPLIT distance="1000" swimtime="00:12:57.30" />
                    <SPLIT distance="1050" swimtime="00:13:36.97" />
                    <SPLIT distance="1100" swimtime="00:14:16.73" />
                    <SPLIT distance="1150" swimtime="00:14:55.72" />
                    <SPLIT distance="1200" swimtime="00:15:35.52" />
                    <SPLIT distance="1250" swimtime="00:16:14.87" />
                    <SPLIT distance="1300" swimtime="00:16:54.34" />
                    <SPLIT distance="1350" swimtime="00:17:32.49" />
                    <SPLIT distance="1400" swimtime="00:18:12.08" />
                    <SPLIT distance="1450" swimtime="00:18:50.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-12" firstname="Marcin" gender="M" lastname="Szymkowiak" nation="POL" license="500115700523" athleteid="8916">
              <RESULTS>
                <RESULT eventid="1195" points="494" reactiontime="+83" swimtime="00:00:26.45" resultid="8917" heatid="9331" lane="8" entrytime="00:00:25.48" />
                <RESULT eventid="1544" points="514" reactiontime="+71" swimtime="00:00:58.56" resultid="8918" heatid="9488" lane="5" entrytime="00:00:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5297" points="567" reactiontime="+69" swimtime="00:01:09.01" resultid="8919" heatid="9513" lane="8" entrytime="00:01:09.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="491" reactiontime="+75" swimtime="00:00:28.43" resultid="8920" heatid="9527" lane="2" entrytime="00:00:27.50" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5585" points="578" reactiontime="+67" swimtime="00:00:31.14" resultid="8921" heatid="9605" lane="0" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WARTA 4" number="4">
              <RESULTS>
                <RESULT eventid="1612" points="498" reactiontime="+70" swimtime="00:01:57.87" resultid="9002" heatid="9499" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="150" swimtime="00:01:30.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8995" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="8916" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="8936" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="8943" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 5" number="5">
              <RESULTS>
                <RESULT eventid="1612" points="405" reactiontime="+76" swimtime="00:02:06.19" resultid="9003" heatid="9499" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:37.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8841" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="8848" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="8922" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="8868" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 8" number="8">
              <RESULTS>
                <RESULT eventid="5433" points="415" reactiontime="+69" swimtime="00:01:53.69" resultid="9010" heatid="9561" lane="8" entrytime="00:01:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                    <SPLIT distance="100" swimtime="00:00:54.33" />
                    <SPLIT distance="150" swimtime="00:01:24.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8943" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="8922" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="8841" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="8930" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 9" number="9">
              <RESULTS>
                <RESULT eventid="5433" points="480" reactiontime="+71" swimtime="00:01:48.34" resultid="9005" heatid="9561" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="100" swimtime="00:00:52.34" />
                    <SPLIT distance="150" swimtime="00:01:19.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8916" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8936" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="8848" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="8868" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="WARTA 3" number="3">
              <RESULTS>
                <RESULT eventid="1595" points="213" reactiontime="+123" swimtime="00:02:57.64" resultid="9001" heatid="9497" lane="6" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                    <SPLIT distance="150" swimtime="00:02:08.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8860" number="1" reactiontime="+123" />
                    <RELAYPOSITION athleteid="8831" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8975" number="3" />
                    <RELAYPOSITION athleteid="8908" number="4" reactiontime="+93" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="WARTA 6" number="6">
              <RESULTS>
                <RESULT eventid="5416" points="171" swimtime="00:02:53.96" resultid="9004" heatid="9559" lane="6" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                    <SPLIT distance="150" swimtime="00:02:03.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8860" number="1" />
                    <RELAYPOSITION athleteid="8831" number="2" />
                    <RELAYPOSITION athleteid="8879" number="3" />
                    <RELAYPOSITION athleteid="8908" number="4" reactiontime="+99" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="WARTA 7" number="7">
              <RESULTS>
                <RESULT eventid="5416" points="141" swimtime="00:03:05.44" resultid="9006" heatid="9559" lane="7" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.46" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:25.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8981" number="1" />
                    <RELAYPOSITION athleteid="8975" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="8836" number="3" reactiontime="+99" />
                    <RELAYPOSITION athleteid="8899" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" name="WARTA 1" number="1">
              <RESULTS>
                <RESULT eventid="1246" swimtime="00:01:50.48" resultid="8999" heatid="9354" lane="6" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:00:56.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8968" number="1" />
                    <RELAYPOSITION athleteid="8857" number="2" reactiontime="-2" />
                    <RELAYPOSITION athleteid="8894" number="3" />
                    <RELAYPOSITION athleteid="8885" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="WARTA 2" number="2">
              <RESULTS>
                <RESULT eventid="1246" swimtime="00:02:12.37" resultid="9000" heatid="9353" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:43.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8860" number="1" />
                    <RELAYPOSITION athleteid="8831" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="8916" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="8868" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="WARTA 10" number="10">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+125" swimtime="00:02:40.18" resultid="9009" heatid="9607" lane="7" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                    <SPLIT distance="150" swimtime="00:02:11.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8860" number="1" reactiontime="+125" />
                    <RELAYPOSITION athleteid="8831" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="8824" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="8841" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WARTA 11" number="11">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+71" swimtime="00:02:29.54" resultid="9008" heatid="9607" lane="5" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:56.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8943" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="8916" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="8899" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="8975" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" name="WARTA 12" number="12">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+64" swimtime="00:02:02.25" resultid="9007" heatid="9608" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:38.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8968" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="8857" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="8894" number="3" />
                    <RELAYPOSITION athleteid="8885" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA" nation="POL" region="KR" clubid="6417" name="Korona Kraków Masters">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="6490">
              <RESULTS>
                <RESULT eventid="1133" points="225" reactiontime="+102" swimtime="00:00:38.86" resultid="6491" heatid="9308" lane="3" />
                <RESULT eventid="1212" points="155" reactiontime="+87" swimtime="00:03:54.64" resultid="6492" heatid="9338" lane="7" entrytime="00:03:39.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:50.96" />
                    <SPLIT distance="150" swimtime="00:02:59.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="134" reactiontime="+104" swimtime="00:00:52.80" resultid="6493" heatid="9442" lane="0" entrytime="00:00:49.67" />
                <RESULT eventid="1527" points="152" reactiontime="+104" swimtime="00:01:36.86" resultid="6494" heatid="9471" lane="3" entrytime="00:01:26.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="146" reactiontime="+101" swimtime="00:00:46.32" resultid="6495" heatid="9514" lane="4" entrytime="00:00:43.63" />
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="6496" heatid="9544" lane="0" entrytime="00:03:29.24" />
                <RESULT eventid="5499" points="127" swimtime="00:01:50.25" resultid="6497" heatid="9570" lane="1" entrytime="00:01:43.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="150" reactiontime="+100" swimtime="00:00:55.26" resultid="6498" heatid="9591" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz-Musiał" nation="POL" athleteid="6474">
              <RESULTS>
                <RESULT eventid="1212" points="70" reactiontime="+117" swimtime="00:05:05.36" resultid="6475" heatid="9337" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.93" />
                    <SPLIT distance="100" swimtime="00:02:27.51" />
                    <SPLIT distance="150" swimtime="00:03:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="86" reactiontime="+95" swimtime="00:18:15.55" resultid="6476" heatid="9357" lane="5" entrytime="00:16:24.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.97" />
                    <SPLIT distance="100" swimtime="00:01:59.31" />
                    <SPLIT distance="150" swimtime="00:03:07.22" />
                    <SPLIT distance="200" swimtime="00:04:16.81" />
                    <SPLIT distance="250" swimtime="00:07:48.56" />
                    <SPLIT distance="300" swimtime="00:06:36.33" />
                    <SPLIT distance="350" swimtime="00:10:05.77" />
                    <SPLIT distance="400" swimtime="00:08:56.83" />
                    <SPLIT distance="450" swimtime="00:12:27.31" />
                    <SPLIT distance="500" swimtime="00:11:15.77" />
                    <SPLIT distance="550" swimtime="00:14:49.85" />
                    <SPLIT distance="600" swimtime="00:13:38.37" />
                    <SPLIT distance="650" swimtime="00:17:01.13" />
                    <SPLIT distance="700" swimtime="00:16:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="92" reactiontime="+89" swimtime="00:01:54.45" resultid="6477" heatid="9470" lane="3" entrytime="00:01:47.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="41" reactiontime="+107" swimtime="00:05:50.89" resultid="6478" heatid="9491" lane="3" entrytime="00:04:49.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.01" />
                    <SPLIT distance="100" swimtime="00:02:38.53" />
                    <SPLIT distance="150" swimtime="00:04:18.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="68" swimtime="00:02:36.75" resultid="6479" heatid="9500" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="70" reactiontime="+100" swimtime="00:10:43.31" resultid="6480" heatid="9562" lane="0" entrytime="00:09:51.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.31" />
                    <SPLIT distance="100" swimtime="00:02:34.54" />
                    <SPLIT distance="150" swimtime="00:03:59.23" />
                    <SPLIT distance="200" swimtime="00:05:26.39" />
                    <SPLIT distance="250" swimtime="00:06:54.58" />
                    <SPLIT distance="300" swimtime="00:08:26.72" />
                    <SPLIT distance="350" swimtime="00:09:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="54" reactiontime="+100" swimtime="00:02:25.97" resultid="6481" heatid="9569" lane="3" entrytime="00:02:13.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="95" reactiontime="+116" swimtime="00:08:36.81" resultid="6482" heatid="9612" lane="3" entrytime="00:08:16.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                    <SPLIT distance="100" swimtime="00:01:59.05" />
                    <SPLIT distance="150" swimtime="00:03:06.48" />
                    <SPLIT distance="200" swimtime="00:04:12.92" />
                    <SPLIT distance="250" swimtime="00:05:19.45" />
                    <SPLIT distance="300" swimtime="00:06:25.39" />
                    <SPLIT distance="350" swimtime="00:07:32.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="6483">
              <RESULTS>
                <RESULT eventid="1195" points="297" reactiontime="+99" swimtime="00:00:31.31" resultid="6484" heatid="9323" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1476" points="282" reactiontime="+81" swimtime="00:00:36.62" resultid="6485" heatid="9453" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="5331" points="355" reactiontime="+93" swimtime="00:00:31.66" resultid="6486" heatid="9523" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="5365" points="289" reactiontime="+78" swimtime="00:01:18.41" resultid="6487" heatid="9538" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="279" reactiontime="+98" swimtime="00:01:16.19" resultid="6488" heatid="9575" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="302" reactiontime="+97" swimtime="00:00:38.67" resultid="6489" heatid="9602" lane="9" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="6425">
              <RESULTS>
                <RESULT eventid="1195" points="319" reactiontime="+81" swimtime="00:00:30.60" resultid="6426" heatid="9324" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1229" points="337" reactiontime="+74" swimtime="00:02:43.71" resultid="6427" heatid="9346" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:04.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="6428" heatid="9454" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1510" points="350" reactiontime="+90" swimtime="00:02:59.66" resultid="6429" heatid="9467" lane="0" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="306" swimtime="00:01:24.73" resultid="6430" heatid="9510" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6431" heatid="9538" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6432" heatid="9587" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="5585" points="310" reactiontime="+84" swimtime="00:00:38.32" resultid="6433" heatid="9601" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="6447">
              <RESULTS>
                <RESULT eventid="1133" points="315" reactiontime="+93" swimtime="00:00:34.76" resultid="6448" heatid="9312" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1263" points="268" reactiontime="+77" swimtime="00:12:31.80" resultid="6449" heatid="9356" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                    <SPLIT distance="200" swimtime="00:02:58.89" />
                    <SPLIT distance="250" swimtime="00:03:46.89" />
                    <SPLIT distance="300" swimtime="00:04:35.45" />
                    <SPLIT distance="350" swimtime="00:05:24.03" />
                    <SPLIT distance="400" swimtime="00:06:12.82" />
                    <SPLIT distance="450" swimtime="00:07:01.03" />
                    <SPLIT distance="500" swimtime="00:07:49.49" />
                    <SPLIT distance="550" swimtime="00:08:37.06" />
                    <SPLIT distance="600" swimtime="00:09:25.32" />
                    <SPLIT distance="650" swimtime="00:10:12.99" />
                    <SPLIT distance="700" swimtime="00:11:00.96" />
                    <SPLIT distance="750" swimtime="00:11:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="309" reactiontime="+91" swimtime="00:01:16.42" resultid="6450" heatid="9473" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="213" swimtime="00:03:23.66" resultid="6451" heatid="9492" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:35.52" />
                    <SPLIT distance="150" swimtime="00:02:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="243" reactiontime="+89" swimtime="00:00:39.14" resultid="6452" heatid="9515" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="5382" points="285" swimtime="00:02:51.55" resultid="6453" heatid="9546" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="150" swimtime="00:02:10.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="235" reactiontime="+90" swimtime="00:01:29.83" resultid="6454" heatid="9570" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="279" reactiontime="+94" swimtime="00:06:01.74" resultid="6455" heatid="9610" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:11.65" />
                    <SPLIT distance="200" swimtime="00:02:57.85" />
                    <SPLIT distance="250" swimtime="00:03:44.52" />
                    <SPLIT distance="300" swimtime="00:04:30.67" />
                    <SPLIT distance="350" swimtime="00:05:17.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="6514">
              <RESULTS>
                <RESULT eventid="1212" points="301" swimtime="00:03:08.09" resultid="6515" heatid="9339" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:30.09" />
                    <SPLIT distance="150" swimtime="00:02:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="277" reactiontime="+73" swimtime="00:00:41.48" resultid="6516" heatid="9443" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="6517" heatid="9473" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="5279" points="245" reactiontime="+94" swimtime="00:01:42.38" resultid="6518" heatid="9503" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="282" swimtime="00:06:45.88" resultid="6519" heatid="9562" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="150" swimtime="00:02:21.78" />
                    <SPLIT distance="200" swimtime="00:03:14.51" />
                    <SPLIT distance="250" swimtime="00:04:13.54" />
                    <SPLIT distance="300" swimtime="00:05:13.18" />
                    <SPLIT distance="350" swimtime="00:06:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="277" swimtime="00:01:25.07" resultid="6520" heatid="9570" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="6521" heatid="9593" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="6465">
              <RESULTS>
                <RESULT eventid="1133" points="44" reactiontime="+112" swimtime="00:01:07.04" resultid="6466" heatid="9308" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1212" points="36" reactiontime="+108" swimtime="00:06:20.01" resultid="6467" heatid="9337" lane="3" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.71" />
                    <SPLIT distance="100" swimtime="00:03:14.80" />
                    <SPLIT distance="150" swimtime="00:04:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="49" swimtime="00:06:19.62" resultid="6468" heatid="9458" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.99" />
                    <SPLIT distance="100" swimtime="00:03:05.04" />
                    <SPLIT distance="150" swimtime="00:04:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="45" reactiontime="+108" swimtime="00:02:24.64" resultid="6469" heatid="9469" lane="5" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="49" swimtime="00:02:54.22" resultid="6470" heatid="9500" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="16" reactiontime="+117" swimtime="00:01:36.51" resultid="6471" heatid="9514" lane="0" entrytime="00:01:25.00" />
                <RESULT eventid="5568" points="61" reactiontime="+111" swimtime="00:01:14.65" resultid="6472" heatid="9592" lane="9" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="6456">
              <RESULTS>
                <RESULT eventid="1195" points="206" reactiontime="+122" swimtime="00:00:35.39" resultid="6457" heatid="9321" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1280" points="123" swimtime="00:15:08.27" resultid="6458" heatid="9362" lane="6" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                    <SPLIT distance="100" swimtime="00:01:40.06" />
                    <SPLIT distance="150" swimtime="00:02:35.10" />
                    <SPLIT distance="200" swimtime="00:03:31.23" />
                    <SPLIT distance="250" swimtime="00:04:29.01" />
                    <SPLIT distance="300" swimtime="00:05:26.17" />
                    <SPLIT distance="350" swimtime="00:06:24.51" />
                    <SPLIT distance="400" swimtime="00:07:22.57" />
                    <SPLIT distance="450" swimtime="00:08:20.70" />
                    <SPLIT distance="500" swimtime="00:09:19.61" />
                    <SPLIT distance="550" swimtime="00:10:19.48" />
                    <SPLIT distance="600" swimtime="00:11:19.77" />
                    <SPLIT distance="650" swimtime="00:12:19.46" />
                    <SPLIT distance="700" swimtime="00:13:19.26" />
                    <SPLIT distance="750" swimtime="00:14:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="190" swimtime="00:01:21.51" resultid="6459" heatid="9481" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="6460" heatid="9493" lane="5" entrytime="00:04:20.00" />
                <RESULT eventid="5331" points="100" reactiontime="+124" swimtime="00:00:48.32" resultid="6461" heatid="9520" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="5399" points="147" swimtime="00:03:12.96" resultid="6462" heatid="9551" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:02:24.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="71" reactiontime="+129" swimtime="00:01:59.93" resultid="6463" heatid="9573" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="143" swimtime="00:07:00.40" resultid="9620" heatid="9621" lane="5" late="yes" entrytime="00:06:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="6434">
              <RESULTS>
                <RESULT eventid="1133" points="464" reactiontime="+81" swimtime="00:00:30.56" resultid="6435" heatid="9315" lane="9" entrytime="00:00:29.20" />
                <RESULT eventid="1458" points="318" reactiontime="+69" swimtime="00:00:39.61" resultid="6436" heatid="9444" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1527" points="441" swimtime="00:01:07.91" resultid="6437" heatid="9475" lane="6" entrytime="00:01:06.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="382" reactiontime="+83" swimtime="00:00:33.66" resultid="6438" heatid="9517" lane="9" entrytime="00:00:32.50" />
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="6439" heatid="9532" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="5499" points="355" reactiontime="+71" swimtime="00:01:18.30" resultid="6440" heatid="9571" lane="7" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="6418">
              <RESULTS>
                <RESULT eventid="1133" points="461" reactiontime="+72" swimtime="00:00:30.63" resultid="6419" heatid="9314" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1458" points="404" reactiontime="+72" swimtime="00:00:36.60" resultid="6420" heatid="9445" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1527" points="402" reactiontime="+72" swimtime="00:01:10.04" resultid="6421" heatid="9475" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="400" reactiontime="+80" swimtime="00:00:33.14" resultid="6422" heatid="9516" lane="8" entrytime="00:00:35.38" />
                <RESULT eventid="5348" points="360" reactiontime="+65" swimtime="00:01:21.67" resultid="6423" heatid="9533" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="450" reactiontime="+72" swimtime="00:00:38.35" resultid="6424" heatid="9596" lane="0" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="6508">
              <RESULTS>
                <RESULT eventid="1212" points="123" reactiontime="+91" swimtime="00:04:13.54" resultid="6509" heatid="9338" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.58" />
                    <SPLIT distance="100" swimtime="00:02:09.41" />
                    <SPLIT distance="150" swimtime="00:03:18.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="138" reactiontime="+109" swimtime="00:04:28.86" resultid="6511" heatid="9459" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.43" />
                    <SPLIT distance="100" swimtime="00:02:13.27" />
                    <SPLIT distance="150" swimtime="00:03:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="75" swimtime="00:00:57.85" resultid="6512" heatid="9514" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="5382" points="148" reactiontime="+100" swimtime="00:03:33.49" resultid="6513" heatid="9543" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                    <SPLIT distance="100" swimtime="00:01:46.73" />
                    <SPLIT distance="150" swimtime="00:02:40.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="6441">
              <RESULTS>
                <RESULT eventid="1458" status="DNS" swimtime="00:00:00.00" resultid="6442" heatid="9442" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="5314" points="281" swimtime="00:00:37.29" resultid="6443" heatid="9515" lane="1" entrytime="00:00:39.98" />
                <RESULT eventid="5450" points="193" swimtime="00:07:40.68" resultid="6444" heatid="9562" lane="2" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.92" />
                    <SPLIT distance="100" swimtime="00:01:52.89" />
                    <SPLIT distance="150" swimtime="00:02:55.08" />
                    <SPLIT distance="200" swimtime="00:03:55.53" />
                    <SPLIT distance="250" swimtime="00:05:00.64" />
                    <SPLIT distance="300" swimtime="00:06:01.68" />
                    <SPLIT distance="350" swimtime="00:06:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="160" reactiontime="+97" swimtime="00:01:42.01" resultid="6445" heatid="9570" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="202" reactiontime="+89" swimtime="00:03:31.25" resultid="6446" heatid="9580" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                    <SPLIT distance="100" swimtime="00:01:48.20" />
                    <SPLIT distance="150" swimtime="00:02:44.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="6499">
              <RESULTS>
                <RESULT eventid="1133" points="229" reactiontime="+103" swimtime="00:00:38.64" resultid="6500" heatid="9311" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1263" points="157" reactiontime="+102" swimtime="00:14:58.03" resultid="6501" heatid="9357" lane="4" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:39.28" />
                    <SPLIT distance="150" swimtime="00:02:36.10" />
                    <SPLIT distance="200" swimtime="00:03:33.31" />
                    <SPLIT distance="250" swimtime="00:10:17.05" />
                    <SPLIT distance="300" swimtime="00:05:27.84" />
                    <SPLIT distance="350" swimtime="00:12:11.19" />
                    <SPLIT distance="400" swimtime="00:07:24.33" />
                    <SPLIT distance="500" swimtime="00:09:19.30" />
                    <SPLIT distance="600" swimtime="00:11:13.50" />
                    <SPLIT distance="700" swimtime="00:13:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="193" reactiontime="+85" swimtime="00:00:46.78" resultid="6502" heatid="9442" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1561" points="110" swimtime="00:04:14.02" resultid="6503" heatid="9492" lane="9" entrytime="00:04:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                    <SPLIT distance="100" swimtime="00:01:59.84" />
                    <SPLIT distance="150" swimtime="00:03:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="156" reactiontime="+98" swimtime="00:01:47.74" resultid="6504" heatid="9529" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="143" swimtime="00:08:28.62" resultid="6505" heatid="9562" lane="1" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.78" />
                    <SPLIT distance="100" swimtime="00:02:04.96" />
                    <SPLIT distance="150" swimtime="00:03:12.09" />
                    <SPLIT distance="200" swimtime="00:04:20.07" />
                    <SPLIT distance="250" swimtime="00:05:28.33" />
                    <SPLIT distance="300" swimtime="00:06:37.11" />
                    <SPLIT distance="350" swimtime="00:07:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="118" swimtime="00:01:53.08" resultid="6506" heatid="9570" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="147" reactiontime="+109" swimtime="00:07:27.95" resultid="6507" heatid="9612" lane="5" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:40.47" />
                    <SPLIT distance="150" swimtime="00:02:40.20" />
                    <SPLIT distance="200" swimtime="00:03:38.65" />
                    <SPLIT distance="250" swimtime="00:04:37.48" />
                    <SPLIT distance="300" swimtime="00:05:35.45" />
                    <SPLIT distance="350" swimtime="00:06:33.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1595" points="381" reactiontime="+79" swimtime="00:02:26.39" resultid="6522" heatid="9497" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:20.21" />
                    <SPLIT distance="150" swimtime="00:01:56.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6447" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6418" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="6514" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6434" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5416" points="419" reactiontime="+76" swimtime="00:02:09.05" resultid="6523" heatid="9559" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6418" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6441" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="6447" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="6434" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+80" swimtime="00:02:02.46" resultid="6524" heatid="9354" lane="8" entrytime="00:02:00.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:00.50" />
                    <SPLIT distance="150" swimtime="00:01:31.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6434" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6418" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6483" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="6425" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5602" reactiontime="+65" swimtime="00:02:17.06" resultid="6525" heatid="9608" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6425" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="6418" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="6483" number="3" />
                    <RELAYPOSITION athleteid="6434" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STIL" nation="POL" region="LBS" clubid="5942" name="Kp Stilon Gorzów Wlkp">
          <CONTACT city="Gorzów Wlkp" email="pstilon@hotmail.com" internet="http://www.kpstilon.gorzow.eu/index.php?p=1_5_kontakt" name="K. Świderski" phone="512 428 265" state="LUBUS" street="UL. Słowiańska 1/ 42" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="5943">
              <RESULTS>
                <RESULT eventid="1314" points="151" swimtime="00:27:12.61" resultid="5944" heatid="9367" lane="7" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:40.05" />
                    <SPLIT distance="150" swimtime="00:02:35.17" />
                    <SPLIT distance="200" swimtime="00:03:30.16" />
                    <SPLIT distance="250" swimtime="00:04:24.97" />
                    <SPLIT distance="300" swimtime="00:05:19.86" />
                    <SPLIT distance="350" swimtime="00:06:14.82" />
                    <SPLIT distance="400" swimtime="00:07:09.75" />
                    <SPLIT distance="450" swimtime="00:08:04.67" />
                    <SPLIT distance="500" swimtime="00:08:59.79" />
                    <SPLIT distance="550" swimtime="00:09:54.71" />
                    <SPLIT distance="600" swimtime="00:10:50.14" />
                    <SPLIT distance="650" swimtime="00:11:45.28" />
                    <SPLIT distance="700" swimtime="00:12:40.37" />
                    <SPLIT distance="750" swimtime="00:13:35.76" />
                    <SPLIT distance="800" swimtime="00:14:30.85" />
                    <SPLIT distance="850" swimtime="00:15:25.57" />
                    <SPLIT distance="900" swimtime="00:16:20.88" />
                    <SPLIT distance="950" swimtime="00:17:15.92" />
                    <SPLIT distance="1000" swimtime="00:18:10.57" />
                    <SPLIT distance="1050" swimtime="00:19:05.69" />
                    <SPLIT distance="1100" swimtime="00:20:00.13" />
                    <SPLIT distance="1150" swimtime="00:20:54.89" />
                    <SPLIT distance="1200" swimtime="00:21:50.25" />
                    <SPLIT distance="1250" swimtime="00:22:45.28" />
                    <SPLIT distance="1300" swimtime="00:23:40.48" />
                    <SPLIT distance="1350" swimtime="00:24:35.25" />
                    <SPLIT distance="1400" swimtime="00:25:29.84" />
                    <SPLIT distance="1450" swimtime="00:26:23.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="131" swimtime="00:01:32.14" resultid="5945" heatid="9479" lane="9" entrytime="00:01:33.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="126" reactiontime="+120" swimtime="00:03:23.26" resultid="5946" heatid="9550" lane="3" entrytime="00:03:26.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:38.98" />
                    <SPLIT distance="150" swimtime="00:02:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="73" reactiontime="+91" swimtime="00:04:26.72" resultid="5947" heatid="9584" lane="5" entrytime="00:04:08.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.27" />
                    <SPLIT distance="100" swimtime="00:02:12.77" />
                    <SPLIT distance="150" swimtime="00:03:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="133" reactiontime="+110" swimtime="00:07:10.95" resultid="5948" heatid="9618" lane="0" entrytime="00:06:52.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:40.85" />
                    <SPLIT distance="150" swimtime="00:02:37.46" />
                    <SPLIT distance="200" swimtime="00:03:33.51" />
                    <SPLIT distance="250" swimtime="00:04:28.92" />
                    <SPLIT distance="300" swimtime="00:05:25.84" />
                    <SPLIT distance="350" swimtime="00:06:20.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PŁYWAK" nation="POL" region="WAR" clubid="8302" name="KPiRS PŁYWAK Płock">
          <CONTACT city="Płock" email="pawel.powichrowski@wp.pl" name="Powichrowski Paweł" phone="603694397" state="MAZ" street="Wiatraki 11 B" zip="09-402" />
          <ATHLETES>
            <ATHLETE birthdate="1997-06-02" firstname="Katarzyna" gender="F" lastname="Janiszkiewicz" nation="POL" athleteid="8303">
              <RESULTS>
                <RESULT eventid="1133" points="411" reactiontime="+80" swimtime="00:00:31.82" resultid="8304" heatid="9312" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1493" points="312" swimtime="00:03:25.00" resultid="8305" heatid="9459" lane="6" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:38.52" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="338" reactiontime="+89" swimtime="00:01:14.20" resultid="8306" heatid="9474" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="329" swimtime="00:01:32.89" resultid="8307" heatid="9502" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="8308" heatid="9545" lane="9" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-05-02" firstname="Jakub" gender="M" lastname="Cichocki" nation="POL" athleteid="8309">
              <RESULTS>
                <RESULT eventid="1195" points="428" reactiontime="+77" swimtime="00:00:27.74" resultid="8310" heatid="9327" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1229" points="316" swimtime="00:02:47.34" resultid="8311" heatid="9348" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="150" swimtime="00:02:00.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="289" swimtime="00:03:11.39" resultid="8312" heatid="9467" lane="9" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="150" swimtime="00:02:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="370" reactiontime="+75" swimtime="00:01:05.29" resultid="8313" heatid="9486" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="295" swimtime="00:01:25.80" resultid="8314" heatid="9512" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-02-06" firstname="Dominik" gender="M" lastname="Bruchajzer" nation="POL" athleteid="8315">
              <RESULTS>
                <RESULT eventid="1195" points="412" reactiontime="+69" swimtime="00:00:28.08" resultid="8316" heatid="9329" lane="0" entrytime="00:00:27.00" />
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie." eventid="1476" reactiontime="+71" status="DSQ" swimtime="00:00:32.33" resultid="8317" heatid="9453" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1544" points="453" swimtime="00:01:01.07" resultid="8318" heatid="9488" lane="6" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="330" reactiontime="+76" swimtime="00:01:15.01" resultid="8319" heatid="9540" lane="0" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="8320" heatid="9557" lane="9" entrytime="00:02:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KM" nation="UKR" clubid="7785" name="Kryvbas Masters">
          <CONTACT city="Krivoy Rog" email="elmartienko@ukr.net" name="Martienko Evgeniy Leonidovich" phone="+38 067 564 2476" street="Prospect Pivdennyi b.25, kv.37" zip="50026" />
          <ATHLETES>
            <ATHLETE birthdate="1948-10-30" firstname="Lukash" gender="M" lastname="Kotseba" nation="UKR" athleteid="7786">
              <RESULTS>
                <RESULT eventid="1510" status="DNS" swimtime="00:00:00.00" resultid="7788" heatid="9462" lane="4" entrytime="00:04:50.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="7789" heatid="9535" lane="6" entrytime="00:01:58.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="7790" heatid="9584" lane="8" entrytime="00:04:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02203" nation="POL" region="LU" clubid="6706" name="Ks Azs Awf Biała Podlaska">
          <CONTACT city="Biała Podlaska" email="mielnik_pawel@wpl.pl" name="Mielnik" phone="697552772" state="LUB" street="Akademicka 2" zip="21-500" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-30" firstname="Wojciech" gender="M" lastname="Suszek" nation="POL" license="102203700023" athleteid="6707">
              <RESULTS>
                <RESULT eventid="1195" points="622" reactiontime="+61" swimtime="00:00:24.49" resultid="6708" heatid="9332" lane="3" entrytime="00:00:23.86" entrycourse="LCM" />
                <RESULT eventid="1229" points="439" reactiontime="+64" swimtime="00:02:29.94" resultid="6709" heatid="9342" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                    <SPLIT distance="150" swimtime="00:01:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="524" reactiontime="+61" swimtime="00:00:29.80" resultid="6710" heatid="9457" lane="7" entrytime="00:00:29.29" entrycourse="LCM" />
                <RESULT eventid="1544" points="663" reactiontime="+64" swimtime="00:00:53.78" resultid="6711" heatid="9490" lane="5" entrytime="00:00:53.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="598" reactiontime="+65" swimtime="00:00:26.62" resultid="6712" heatid="9528" lane="1" entrytime="00:00:26.16" entrycourse="LCM" />
                <RESULT eventid="5365" points="427" reactiontime="+61" swimtime="00:01:08.85" resultid="6713" heatid="9541" lane="8" entrytime="00:01:05.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="557" swimtime="00:01:00.54" resultid="6714" heatid="9572" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="350" reactiontime="+60" swimtime="00:02:38.75" resultid="6715" heatid="9583" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:16.33" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="6051" name="Ks Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANOWOL@POCZTA.ONET.PL" name="WOLNIEWICZ JANUSZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="6052">
              <RESULTS>
                <RESULT eventid="1195" points="182" reactiontime="+100" swimtime="00:00:36.87" resultid="6053" heatid="9320" lane="2" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1314" points="99" swimtime="00:31:17.69" resultid="6054" heatid="9367" lane="1" entrytime="00:29:10.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:45.80" />
                    <SPLIT distance="150" swimtime="00:02:45.90" />
                    <SPLIT distance="200" swimtime="00:03:47.27" />
                    <SPLIT distance="250" swimtime="00:04:48.77" />
                    <SPLIT distance="300" swimtime="00:05:50.39" />
                    <SPLIT distance="350" swimtime="00:06:52.40" />
                    <SPLIT distance="400" swimtime="00:07:54.72" />
                    <SPLIT distance="450" swimtime="00:08:57.62" />
                    <SPLIT distance="500" swimtime="00:10:00.48" />
                    <SPLIT distance="550" swimtime="00:11:03.94" />
                    <SPLIT distance="600" swimtime="00:12:07.53" />
                    <SPLIT distance="650" swimtime="00:13:10.49" />
                    <SPLIT distance="700" swimtime="00:14:13.70" />
                    <SPLIT distance="750" swimtime="00:15:17.52" />
                    <SPLIT distance="800" swimtime="00:16:22.32" />
                    <SPLIT distance="850" swimtime="00:17:26.62" />
                    <SPLIT distance="900" swimtime="00:18:30.42" />
                    <SPLIT distance="950" swimtime="00:19:34.51" />
                    <SPLIT distance="1000" swimtime="00:20:38.48" />
                    <SPLIT distance="1050" swimtime="00:21:43.69" />
                    <SPLIT distance="1100" swimtime="00:22:48.05" />
                    <SPLIT distance="1150" swimtime="00:23:52.40" />
                    <SPLIT distance="1200" swimtime="00:24:56.74" />
                    <SPLIT distance="1250" swimtime="00:26:01.62" />
                    <SPLIT distance="1300" swimtime="00:27:05.21" />
                    <SPLIT distance="1350" swimtime="00:28:09.50" />
                    <SPLIT distance="1400" swimtime="00:29:14.04" />
                    <SPLIT distance="1450" swimtime="00:30:17.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6055" heatid="9479" lane="1" entrytime="00:01:30.80" entrycourse="SCM" />
                <RESULT eventid="5399" points="115" swimtime="00:03:29.15" resultid="6056" heatid="9550" lane="6" entrytime="00:03:28.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="102" reactiontime="+114" swimtime="00:07:49.64" resultid="6057" heatid="9619" lane="3" entrytime="00:07:41.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                    <SPLIT distance="100" swimtime="00:01:45.09" />
                    <SPLIT distance="150" swimtime="00:02:46.22" />
                    <SPLIT distance="200" swimtime="00:03:48.01" />
                    <SPLIT distance="250" swimtime="00:04:50.07" />
                    <SPLIT distance="300" swimtime="00:05:51.81" />
                    <SPLIT distance="350" swimtime="00:06:53.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="5984" name="KS Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="5985">
              <RESULTS>
                <RESULT eventid="1229" points="298" reactiontime="+90" swimtime="00:02:50.65" resultid="5986" heatid="9346" lane="8" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="329" swimtime="00:03:03.45" resultid="5987" heatid="9466" lane="1" entrytime="00:03:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:28.83" />
                    <SPLIT distance="150" swimtime="00:02:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="322" swimtime="00:01:23.35" resultid="5988" heatid="9510" lane="1" entrytime="00:01:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="291" reactiontime="+81" swimtime="00:01:18.21" resultid="5989" heatid="9539" lane="8" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="273" reactiontime="+90" swimtime="00:02:52.32" resultid="5990" heatid="9588" lane="2" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                    <SPLIT distance="150" swimtime="00:02:10.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KS PŁETWAL" nation="POL" region="KR" clubid="6285" name="KS Płetwal Zakopane">
          <CONTACT city="Zakopane" email="mdylag@op.pl" name="Dyląg" phone="605075837" state="MAL" zip="34-500" />
          <ATHLETES>
            <ATHLETE birthdate="1968-04-22" firstname="Maciej" gender="M" lastname="Haras" nation="POL" license="104206700018" athleteid="6306">
              <RESULTS>
                <RESULT eventid="5297" points="369" reactiontime="+66" swimtime="00:01:19.62" resultid="6307" heatid="9511" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="399" reactiontime="+81" swimtime="00:00:35.22" resultid="6308" heatid="9603" lane="9" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="7185" name="Ks Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1992-02-23" firstname="Tomasz" gender="M" lastname="Janczyk" nation="POL" athleteid="8379">
              <RESULTS>
                <RESULT eventid="1195" points="306" reactiontime="+72" swimtime="00:00:31.02" resultid="8380" heatid="9326" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="8381" heatid="9453" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="5365" reactiontime="+82" status="DNS" swimtime="00:00:00.00" resultid="8382" heatid="9541" lane="0" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="8373">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="8374" heatid="9314" lane="3" entrytime="00:00:29.90" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="8375" heatid="9461" lane="6" entrytime="00:02:59.90" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="8376" heatid="9475" lane="4" entrytime="00:01:04.90" />
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="8377" heatid="9504" lane="8" entrytime="00:01:25.90" />
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="8378" heatid="9595" lane="4" entrytime="00:00:38.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-10" firstname="Piotr" gender="M" lastname="Tatarynowicz" nation="POL" athleteid="7192">
              <RESULTS>
                <RESULT comment="O8 - Pływak uczestniczył w wyścigu z naklejonym plastrem, który nie został wcześniej zatwierdzony." eventid="1476" reactiontime="+64" status="DSQ" swimtime="00:00:29.86" resultid="7193" heatid="9457" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="5365" points="515" reactiontime="+65" swimtime="00:01:04.67" resultid="7194" heatid="9541" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="462" reactiontime="+69" swimtime="00:02:24.68" resultid="7195" heatid="9590" lane="6" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                    <SPLIT distance="150" swimtime="00:01:47.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-10" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="8364">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="8365" heatid="9329" lane="7" entrytime="00:00:26.90" />
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="8366" heatid="9348" lane="3" entrytime="00:02:29.90" />
                <RESULT eventid="1476" points="521" reactiontime="+66" swimtime="00:00:29.87" resultid="8367" heatid="9457" lane="8" entrytime="00:00:29.90" />
                <RESULT eventid="1578" points="324" reactiontime="+79" swimtime="00:02:42.27" resultid="8368" heatid="9496" lane="0" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="501" reactiontime="+76" swimtime="00:00:28.24" resultid="8369" heatid="9526" lane="5" entrytime="00:00:28.90" />
                <RESULT eventid="5365" points="492" reactiontime="+60" swimtime="00:01:05.66" resultid="8370" heatid="9541" lane="2" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="482" swimtime="00:01:03.54" resultid="8371" heatid="9577" lane="6" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="413" reactiontime="+60" swimtime="00:02:30.18" resultid="8372" heatid="9590" lane="8" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:50.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="7196">
              <RESULTS>
                <RESULT eventid="1195" points="496" reactiontime="+73" swimtime="00:00:26.41" resultid="7197" heatid="9331" lane="2" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1229" points="388" reactiontime="+85" swimtime="00:02:36.17" resultid="7198" heatid="9348" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:11.86" />
                    <SPLIT distance="150" swimtime="00:01:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="464" reactiontime="+73" swimtime="00:00:31.04" resultid="7199" heatid="9456" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1544" points="495" reactiontime="+74" swimtime="00:00:59.30" resultid="7200" heatid="9487" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="484" reactiontime="+78" swimtime="00:00:28.55" resultid="7201" heatid="9527" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="5365" points="395" reactiontime="+97" swimtime="00:01:10.63" resultid="7202" heatid="9541" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="398" reactiontime="+79" swimtime="00:00:35.26" resultid="7203" heatid="9602" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="7204">
              <RESULTS>
                <RESULT eventid="1195" points="506" reactiontime="+71" swimtime="00:00:26.24" resultid="7205" heatid="9331" lane="3" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1544" points="523" reactiontime="+64" swimtime="00:00:58.22" resultid="7206" heatid="9489" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1229" points="355" swimtime="00:02:40.99" resultid="8361" heatid="9348" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:02:03.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="310" reactiontime="+72" swimtime="00:01:13.59" resultid="8362" heatid="9576" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="389" reactiontime="+77" swimtime="00:00:35.53" resultid="8363" heatid="9602" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-22" firstname="Jacek" gender="M" lastname="Hankus" nation="POL" athleteid="8383">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="8384" heatid="9328" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="5331" points="245" reactiontime="+92" swimtime="00:00:35.81" resultid="8385" heatid="9526" lane="9" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="7186">
              <RESULTS>
                <RESULT eventid="1133" points="344" reactiontime="+85" swimtime="00:00:33.75" resultid="7187" heatid="9312" lane="3" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1493" points="209" reactiontime="+104" swimtime="00:03:54.40" resultid="7188" heatid="9458" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:51.74" />
                    <SPLIT distance="150" swimtime="00:02:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="241" reactiontime="+101" swimtime="00:01:33.33" resultid="7189" heatid="9529" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="284" swimtime="00:02:51.72" resultid="7190" heatid="9545" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:22.19" />
                    <SPLIT distance="150" swimtime="00:02:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="235" reactiontime="+104" swimtime="00:03:21.03" resultid="7191" heatid="9581" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                    <SPLIT distance="100" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:02:30.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="REKIN Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="434" reactiontime="+69" swimtime="00:02:03.38" resultid="8386" heatid="9499" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:33.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8383" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="7196" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="7204" number="3" reactiontime="+7" />
                    <RELAYPOSITION athleteid="7192" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5433" points="471" swimtime="00:01:48.98" resultid="8387" heatid="9561" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:00:57.10" />
                    <SPLIT distance="150" swimtime="00:01:23.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8383" number="1" />
                    <RELAYPOSITION athleteid="8379" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="7192" number="3" />
                    <RELAYPOSITION athleteid="7196" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="REKIN Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="1246" status="DNS" swimtime="00:00:00.00" resultid="8388" heatid="9354" lane="7" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8373" number="1" />
                    <RELAYPOSITION athleteid="8364" number="2" />
                    <RELAYPOSITION athleteid="7186" number="3" />
                    <RELAYPOSITION athleteid="7196" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5602" reactiontime="+68" swimtime="00:02:14.64" resultid="8389" heatid="9608" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:42.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8364" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="8373" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="7196" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="7186" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="SLA" clubid="6350" name="KS. Górnik Radlin">
          <ATHLETES>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="6351">
              <RESULTS>
                <RESULT eventid="1133" points="482" reactiontime="+88" swimtime="00:00:30.17" resultid="6352" heatid="9313" lane="5" entrytime="00:00:31.90" />
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /O2" eventid="1212" status="DSQ" swimtime="00:02:54.72" resultid="6353" heatid="9340" lane="9" entrytime="00:02:48.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="150" swimtime="00:02:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="476" reactiontime="+81" swimtime="00:01:06.21" resultid="6354" heatid="9475" lane="2" entrytime="00:01:06.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="404" reactiontime="+87" swimtime="00:00:33.03" resultid="6355" heatid="9516" lane="4" entrytime="00:00:32.59" />
                <RESULT eventid="5568" points="395" swimtime="00:00:40.06" resultid="6356" heatid="9596" lane="9" entrytime="00:00:38.89" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="WIE" clubid="7908" name="KU AZS UAM Poznań">
          <CONTACT email="swimteamuam@gmail.com" name="Sterczyński" phone="693840114" />
          <ATHLETES>
            <ATHLETE birthdate="1979-04-05" firstname="Anna" gender="F" lastname="Walkowiak" nation="POL" athleteid="7967">
              <RESULTS>
                <RESULT eventid="1133" points="388" swimtime="00:00:32.44" resultid="7968" heatid="9313" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="5314" points="323" reactiontime="+90" swimtime="00:00:35.60" resultid="7969" heatid="9515" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="7970" heatid="9582" lane="9" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="7947">
              <RESULTS>
                <RESULT eventid="1195" points="334" reactiontime="+91" swimtime="00:00:30.13" resultid="7948" heatid="9326" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1280" points="250" reactiontime="+99" swimtime="00:11:57.37" resultid="7949" heatid="9361" lane="4" entrytime="00:11:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:03.03" />
                    <SPLIT distance="200" swimtime="00:02:47.89" />
                    <SPLIT distance="250" swimtime="00:05:05.55" />
                    <SPLIT distance="300" swimtime="00:04:19.57" />
                    <SPLIT distance="350" swimtime="00:06:36.98" />
                    <SPLIT distance="400" swimtime="00:05:51.35" />
                    <SPLIT distance="450" swimtime="00:08:09.44" />
                    <SPLIT distance="500" swimtime="00:07:23.21" />
                    <SPLIT distance="550" swimtime="00:09:42.37" />
                    <SPLIT distance="600" swimtime="00:08:55.91" />
                    <SPLIT distance="700" swimtime="00:10:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="308" reactiontime="+84" swimtime="00:01:09.40" resultid="7950" heatid="9483" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="268" swimtime="00:02:38.10" resultid="7951" heatid="9555" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:57.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-13" firstname="Kamil" gender="M" lastname="Bernaś" nation="POL" athleteid="7972">
              <RESULTS>
                <RESULT eventid="1195" points="401" reactiontime="+94" swimtime="00:00:28.34" resultid="7973" heatid="9329" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="1544" points="389" reactiontime="+66" swimtime="00:01:04.26" resultid="7974" heatid="9484" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="352" reactiontime="+78" swimtime="00:00:31.74" resultid="7975" heatid="9525" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-18" firstname="Marek" gender="M" lastname="Michałkowski" nation="POL" athleteid="7963">
              <RESULTS>
                <RESULT eventid="1544" points="532" reactiontime="+65" swimtime="00:00:57.88" resultid="7964" heatid="9489" lane="3" entrytime="00:00:56.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="495" swimtime="00:01:12.21" resultid="7965" heatid="9513" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="545" reactiontime="+72" swimtime="00:00:31.76" resultid="7966" heatid="9605" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="7921">
              <RESULTS>
                <RESULT eventid="1195" points="464" reactiontime="+72" swimtime="00:00:27.00" resultid="7922" heatid="9330" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1229" points="429" reactiontime="+73" swimtime="00:02:31.09" resultid="7923" heatid="9349" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="458" reactiontime="+76" swimtime="00:00:31.17" resultid="7924" heatid="9457" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="5331" points="493" reactiontime="+64" swimtime="00:00:28.39" resultid="7925" heatid="9526" lane="1" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-27" firstname="Maciej" gender="M" lastname="Waliński" nation="POL" athleteid="7937">
              <RESULTS>
                <RESULT eventid="1195" points="368" reactiontime="+65" swimtime="00:00:29.17" resultid="7938" heatid="9324" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1544" points="347" reactiontime="+63" swimtime="00:01:06.74" resultid="7939" heatid="9482" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="236" reactiontime="+72" swimtime="00:00:36.29" resultid="7940" heatid="9521" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="5399" points="267" reactiontime="+70" swimtime="00:02:38.30" resultid="7941" heatid="9555" lane="0" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-09-22" firstname="Bartosz" gender="M" lastname="Ziemniarski" nation="POL" athleteid="7930">
              <RESULTS>
                <RESULT eventid="1195" points="543" reactiontime="+72" swimtime="00:00:25.62" resultid="7931" heatid="9331" lane="1" entrytime="00:00:25.39" />
                <RESULT eventid="1544" points="552" reactiontime="+74" swimtime="00:00:57.17" resultid="7932" heatid="9489" lane="2" entrytime="00:00:57.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="487" reactiontime="+73" swimtime="00:02:09.62" resultid="7933" heatid="9558" lane="0" entrytime="00:02:09.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="100" swimtime="00:01:00.23" />
                    <SPLIT distance="150" swimtime="00:01:34.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-24" firstname="Helena" gender="F" lastname="Rachwał" nation="POL" athleteid="7971" />
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Sterczyńska" nation="POL" athleteid="7915">
              <RESULTS>
                <RESULT eventid="1133" points="599" reactiontime="+81" swimtime="00:00:28.07" resultid="7916" heatid="9315" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1458" points="485" reactiontime="+73" swimtime="00:00:34.43" resultid="7917" heatid="9446" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1527" points="594" swimtime="00:01:01.51" resultid="7918" heatid="9476" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="437" reactiontime="+78" swimtime="00:00:32.17" resultid="7919" heatid="9517" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="5568" points="507" reactiontime="+81" swimtime="00:00:36.86" resultid="7920" heatid="9596" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-05" firstname="Marek" gender="M" lastname="Serafin" nation="POL" athleteid="7926">
              <RESULTS>
                <RESULT eventid="1195" points="281" reactiontime="+64" swimtime="00:00:31.92" resultid="7927" heatid="9321" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="5331" points="166" reactiontime="+92" swimtime="00:00:40.77" resultid="7928" heatid="9520" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="5399" points="213" reactiontime="+90" swimtime="00:02:50.72" resultid="7929" heatid="9551" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:09.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-20" firstname="Krzysztof" gender="M" lastname="Strzelczyk" nation="POL" athleteid="7909">
              <RESULTS>
                <RESULT eventid="1195" points="201" reactiontime="+92" swimtime="00:00:35.64" resultid="7910" heatid="9321" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1544" points="190" reactiontime="+84" swimtime="00:01:21.59" resultid="7911" heatid="9480" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="163" reactiontime="+86" swimtime="00:00:40.99" resultid="7912" heatid="9520" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="5399" points="150" reactiontime="+97" swimtime="00:03:11.55" resultid="7913" heatid="9551" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="150" swimtime="00:02:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" status="DNS" swimtime="00:00:00.00" resultid="7914" heatid="9618" lane="5" entrytime="00:06:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" license="103315200006" athleteid="7952">
              <RESULTS>
                <RESULT eventid="1195" points="581" reactiontime="+70" swimtime="00:00:25.05" resultid="7953" heatid="9332" lane="8" entrytime="00:00:24.50" />
                <RESULT eventid="1476" points="607" reactiontime="+79" swimtime="00:00:28.39" resultid="7954" heatid="9457" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="5331" points="660" reactiontime="+67" swimtime="00:00:25.75" resultid="7955" heatid="9528" lane="4" entrytime="00:00:24.90" />
                <RESULT eventid="5365" points="602" reactiontime="+65" swimtime="00:01:01.38" resultid="7956" heatid="9541" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="643" reactiontime="+67" swimtime="00:00:57.71" resultid="7957" heatid="9578" lane="3" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarosław" gender="M" lastname="Bystry" nation="POL" athleteid="7942">
              <RESULTS>
                <RESULT eventid="1195" points="392" reactiontime="+79" swimtime="00:00:28.55" resultid="7943" heatid="9327" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1544" points="381" reactiontime="+73" swimtime="00:01:04.70" resultid="7944" heatid="9484" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="380" reactiontime="+75" swimtime="00:00:30.95" resultid="7945" heatid="9523" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="7946" heatid="9556" lane="0" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-19" firstname="Damian" gender="M" lastname="Kowalik" nation="POL" license="103315200009" athleteid="7958">
              <RESULTS>
                <RESULT eventid="1195" points="578" reactiontime="+66" swimtime="00:00:25.09" resultid="7959" heatid="9332" lane="2" entrytime="00:00:24.21" />
                <RESULT eventid="1544" points="584" reactiontime="+62" swimtime="00:00:56.10" resultid="7960" heatid="9490" lane="8" entrytime="00:00:54.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="634" reactiontime="+66" swimtime="00:00:26.10" resultid="7961" heatid="9528" lane="2" entrytime="00:00:25.36" />
                <RESULT eventid="5517" points="590" reactiontime="+66" swimtime="00:00:59.38" resultid="7962" heatid="9578" lane="5" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-12" firstname="Joanna" gender="F" lastname="Chomicz" nation="POL" athleteid="7934">
              <RESULTS>
                <RESULT eventid="1133" points="336" reactiontime="+68" swimtime="00:00:34.03" resultid="7935" heatid="9313" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1458" points="272" reactiontime="+81" swimtime="00:00:41.73" resultid="7936" heatid="9445" lane="9" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="5433" points="564" reactiontime="+70" swimtime="00:01:42.68" resultid="7981" heatid="9561" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                    <SPLIT distance="100" swimtime="00:00:51.89" />
                    <SPLIT distance="150" swimtime="00:01:16.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7921" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="7963" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="7952" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="7930" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="520" reactiontime="+61" swimtime="00:01:56.14" resultid="7984" heatid="9499" lane="4" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:00:59.47" />
                    <SPLIT distance="150" swimtime="00:01:31.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7952" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="7963" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="7972" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="7930" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="5433" points="382" reactiontime="+79" swimtime="00:01:56.85" resultid="7982" heatid="9561" lane="2" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:00.82" />
                    <SPLIT distance="150" swimtime="00:01:28.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7947" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="7937" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="7972" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="7942" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1612" points="356" reactiontime="+72" swimtime="00:02:11.72" resultid="7983" heatid="9499" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:42.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7921" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7947" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="7942" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7937" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5416" points="487" reactiontime="+87" swimtime="00:02:02.77" resultid="7979" heatid="9559" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="150" swimtime="00:01:35.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7967" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="7971" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7934" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="7915" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1595" points="397" reactiontime="+66" swimtime="00:02:24.48" resultid="7980" heatid="9497" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:01:54.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7934" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="7915" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="7967" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="7971" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1246" reactiontime="+77" swimtime="00:01:50.73" resultid="7976" heatid="9354" lane="3" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:00:57.57" />
                    <SPLIT distance="150" swimtime="00:01:25.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7934" number="1" reactiontime="+77" status="DSQ" />
                    <RELAYPOSITION athleteid="7952" number="2" reactiontime="+20" status="DSQ" />
                    <RELAYPOSITION athleteid="7915" number="3" reactiontime="+15" status="DSQ" />
                    <RELAYPOSITION athleteid="7930" number="4" reactiontime="+20" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+70" swimtime="00:02:04.08" resultid="7977" heatid="9608" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                    <SPLIT distance="150" swimtime="00:01:36.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7967" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="7963" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7952" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="7915" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="5602" status="DNS" swimtime="00:00:00.00" resultid="7978" heatid="9608" lane="3" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7934" number="1" />
                    <RELAYPOSITION athleteid="7921" number="2" />
                    <RELAYPOSITION athleteid="7930" number="3" />
                    <RELAYPOSITION athleteid="7971" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZS WUM" nation="POL" region="WAR" clubid="6327" name="Ku Azs Wum Warszawa">
          <CONTACT email="joogr@hotmail.com" name="Joanna Grzeszczuk" phone="668499613" />
          <ATHLETES>
            <ATHLETE birthdate="1991-02-25" firstname="Joanna" gender="F" lastname="Grzeszczuk" nation="POL" athleteid="6328">
              <RESULTS>
                <RESULT eventid="1458" points="336" reactiontime="+75" swimtime="00:00:38.90" resultid="6329" heatid="9445" lane="0" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="5279" points="518" reactiontime="+72" swimtime="00:01:19.81" resultid="6330" heatid="9504" lane="5" entrytime="00:01:18.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="457" reactiontime="+73" swimtime="00:00:31.71" resultid="6331" heatid="9517" lane="1" entrytime="00:00:31.41" entrycourse="LCM" />
                <RESULT eventid="5568" points="569" reactiontime="+76" swimtime="00:00:35.47" resultid="6332" heatid="9596" lane="5" entrytime="00:00:35.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEG" nation="POL" clubid="7753" name="Legia Warszawa">
          <CONTACT email="agnieszka.kaczmarek85@gmail.vo" name="Kaczmarek" phone="531799855" />
          <ATHLETES>
            <ATHLETE birthdate="1963-05-11" firstname="Maciej" gender="M" lastname="Rybicki" nation="POL" athleteid="7767">
              <RESULTS>
                <RESULT eventid="1195" points="303" reactiontime="+68" swimtime="00:00:31.13" resultid="7768" heatid="9323" lane="0" entrytime="00:00:31.05" />
                <RESULT eventid="1476" points="188" reactiontime="+65" swimtime="00:00:41.90" resultid="7769" heatid="9451" lane="0" entrytime="00:00:42.70" />
                <RESULT eventid="5585" points="239" reactiontime="+73" swimtime="00:00:41.79" resultid="7770" heatid="9599" lane="0" entrytime="00:00:42.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-16" firstname="Adrian" gender="M" lastname="Kulisz" nation="POL" athleteid="7764">
              <RESULTS>
                <RESULT eventid="1544" points="226" swimtime="00:01:16.94" resultid="7765" heatid="9480" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="209" reactiontime="+98" swimtime="00:01:36.17" resultid="7766" heatid="9505" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-04" firstname="Hubert" gender="M" lastname="Markowski" nation="POL" athleteid="7758">
              <RESULTS>
                <RESULT eventid="1229" points="350" swimtime="00:02:41.65" resultid="7759" heatid="9347" lane="1" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="330" reactiontime="+71" swimtime="00:00:34.77" resultid="7760" heatid="9454" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="5365" points="323" reactiontime="+61" swimtime="00:01:15.56" resultid="7761" heatid="9539" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="329" reactiontime="+92" swimtime="00:05:52.86" resultid="7762" heatid="9568" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:01:57.21" />
                    <SPLIT distance="200" swimtime="00:02:45.14" />
                    <SPLIT distance="250" swimtime="00:03:36.38" />
                    <SPLIT distance="300" swimtime="00:04:28.22" />
                    <SPLIT distance="350" swimtime="00:05:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="379" reactiontime="+83" swimtime="00:01:08.84" resultid="7763" heatid="9576" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="7754">
              <RESULTS>
                <RESULT eventid="5297" points="561" reactiontime="+66" swimtime="00:01:09.24" resultid="7755" heatid="9513" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="7756" heatid="9528" lane="9" entrytime="00:00:26.99" />
                <RESULT eventid="5585" points="604" reactiontime="+71" swimtime="00:00:30.69" resultid="7757" heatid="9605" lane="6" entrytime="00:00:29.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MB" nation="POL" clubid="6309" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="DM" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="6314">
              <RESULTS>
                <RESULT eventid="1133" points="233" reactiontime="+77" swimtime="00:00:38.45" resultid="6315" heatid="9311" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1527" points="194" swimtime="00:01:29.27" resultid="6316" heatid="9471" lane="7" entrytime="00:01:27.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="114" reactiontime="+82" swimtime="00:01:59.58" resultid="6317" heatid="9531" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="6318" heatid="9544" lane="8" entrytime="00:03:25.00" />
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="6319" heatid="9580" lane="8" entrytime="00:04:10.00" />
                <RESULT eventid="5619" points="160" swimtime="00:07:15.48" resultid="6320" heatid="9611" lane="7" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:41.55" />
                    <SPLIT distance="150" swimtime="00:02:37.08" />
                    <SPLIT distance="200" swimtime="00:03:33.56" />
                    <SPLIT distance="250" swimtime="00:04:30.32" />
                    <SPLIT distance="300" swimtime="00:05:26.05" />
                    <SPLIT distance="350" swimtime="00:06:22.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="6310">
              <RESULTS>
                <RESULT eventid="1263" points="423" reactiontime="+77" swimtime="00:10:45.56" resultid="6311" heatid="9355" lane="5" entrytime="00:10:24.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:53.80" />
                    <SPLIT distance="200" swimtime="00:02:34.34" />
                    <SPLIT distance="250" swimtime="00:03:14.46" />
                    <SPLIT distance="300" swimtime="00:03:54.95" />
                    <SPLIT distance="350" swimtime="00:04:35.14" />
                    <SPLIT distance="400" swimtime="00:05:15.74" />
                    <SPLIT distance="450" swimtime="00:05:56.47" />
                    <SPLIT distance="500" swimtime="00:06:37.45" />
                    <SPLIT distance="550" swimtime="00:07:18.57" />
                    <SPLIT distance="600" swimtime="00:07:59.97" />
                    <SPLIT distance="650" swimtime="00:08:41.61" />
                    <SPLIT distance="700" swimtime="00:09:23.72" />
                    <SPLIT distance="750" swimtime="00:10:05.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="469" swimtime="00:02:25.40" resultid="6312" heatid="9547" lane="7" entrytime="00:02:22.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="452" reactiontime="+79" swimtime="00:05:08.04" resultid="6313" heatid="9609" lane="3" entrytime="00:05:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                    <SPLIT distance="150" swimtime="00:01:54.30" />
                    <SPLIT distance="200" swimtime="00:02:33.95" />
                    <SPLIT distance="250" swimtime="00:03:12.91" />
                    <SPLIT distance="300" swimtime="00:03:52.07" />
                    <SPLIT distance="350" swimtime="00:04:30.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="6321">
              <RESULTS>
                <RESULT eventid="1510" status="DNS" swimtime="00:00:00.00" resultid="6323" heatid="9464" lane="0" entrytime="00:03:35.00" />
                <RESULT eventid="5297" points="208" swimtime="00:01:36.42" resultid="6324" heatid="9507" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="253" reactiontime="+97" swimtime="00:00:41.02" resultid="6325" heatid="9600" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="5636" points="185" reactiontime="+95" swimtime="00:06:25.58" resultid="6326" heatid="9617" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:16.91" />
                    <SPLIT distance="200" swimtime="00:03:06.30" />
                    <SPLIT distance="250" swimtime="00:03:56.69" />
                    <SPLIT distance="300" swimtime="00:04:47.23" />
                    <SPLIT distance="350" swimtime="00:05:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="199" reactiontime="+98" swimtime="00:00:38.41" resultid="9300" heatid="9521" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKAR" nation="POL" region="RZ" clubid="5853" name="Masters Ikar Mielec">
          <CONTACT email="sebastianboicetta@gmail.com" name="BOICETTA SEBASTIAN" phone="501072284" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-24" firstname="Bartek" gender="M" lastname="Kowalik" nation="POL" license="503208700001" athleteid="5854">
              <RESULTS>
                <RESULT eventid="1229" points="443" reactiontime="+69" swimtime="00:02:29.44" resultid="5855" heatid="9348" lane="5" entrytime="00:02:29.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="150" swimtime="00:01:51.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="5856" heatid="9567" lane="5" entrytime="00:05:30.00" />
                <RESULT eventid="5551" points="376" reactiontime="+83" swimtime="00:02:34.94" resultid="5857" heatid="9590" lane="1" entrytime="00:02:28.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" status="OTL" swimtime="00:11:05.72" resultid="5865" heatid="9359" lane="6" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:49.94" />
                    <SPLIT distance="200" swimtime="00:02:30.77" />
                    <SPLIT distance="250" swimtime="00:03:12.53" />
                    <SPLIT distance="300" swimtime="00:03:54.39" />
                    <SPLIT distance="350" swimtime="00:04:37.02" />
                    <SPLIT distance="400" swimtime="00:05:20.45" />
                    <SPLIT distance="450" swimtime="00:06:04.03" />
                    <SPLIT distance="500" swimtime="00:06:47.91" />
                    <SPLIT distance="550" swimtime="00:07:31.81" />
                    <SPLIT distance="600" swimtime="00:08:15.14" />
                    <SPLIT distance="650" swimtime="00:08:58.36" />
                    <SPLIT distance="700" swimtime="00:09:41.85" />
                    <SPLIT distance="750" swimtime="00:10:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1510" reactiontime="+46" status="DSQ" swimtime="00:02:37.31" resultid="5866" heatid="9468" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="551" reactiontime="+72" swimtime="00:01:09.68" resultid="5867" heatid="9513" lane="2" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="525" reactiontime="+78" swimtime="00:00:32.16" resultid="5868" heatid="9605" lane="9" entrytime="00:00:31.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" license="503208700002" athleteid="5858">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1314" points="471" reactiontime="+76" swimtime="00:18:38.97" resultid="5859" heatid="9365" lane="3" entrytime="00:18:44.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.98" />
                    <SPLIT distance="200" swimtime="00:02:19.45" />
                    <SPLIT distance="250" swimtime="00:02:55.90" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                    <SPLIT distance="350" swimtime="00:04:10.36" />
                    <SPLIT distance="400" swimtime="00:04:48.23" />
                    <SPLIT distance="450" swimtime="00:05:25.85" />
                    <SPLIT distance="500" swimtime="00:06:04.33" />
                    <SPLIT distance="550" swimtime="00:06:41.99" />
                    <SPLIT distance="600" swimtime="00:07:20.22" />
                    <SPLIT distance="650" swimtime="00:07:58.23" />
                    <SPLIT distance="700" swimtime="00:08:36.59" />
                    <SPLIT distance="750" swimtime="00:09:14.13" />
                    <SPLIT distance="800" swimtime="00:09:52.33" />
                    <SPLIT distance="850" swimtime="00:10:29.76" />
                    <SPLIT distance="900" swimtime="00:11:08.38" />
                    <SPLIT distance="950" swimtime="00:11:45.50" />
                    <SPLIT distance="1000" swimtime="00:12:23.73" />
                    <SPLIT distance="1050" swimtime="00:13:01.35" />
                    <SPLIT distance="1100" swimtime="00:13:39.53" />
                    <SPLIT distance="1150" swimtime="00:14:17.64" />
                    <SPLIT distance="1200" swimtime="00:14:55.50" />
                    <SPLIT distance="1250" swimtime="00:15:33.05" />
                    <SPLIT distance="1300" swimtime="00:16:11.31" />
                    <SPLIT distance="1350" swimtime="00:16:48.71" />
                    <SPLIT distance="1400" swimtime="00:17:26.81" />
                    <SPLIT distance="1450" swimtime="00:17:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="498" reactiontime="+79" swimtime="00:02:20.64" resultid="5860" heatid="9496" lane="3" entrytime="00:02:16.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="5861" heatid="9557" lane="1" entrytime="00:02:14.22" />
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="5862" heatid="9567" lane="3" entrytime="00:05:30.44" />
                <RESULT eventid="5517" points="459" reactiontime="+75" swimtime="00:01:04.57" resultid="5863" heatid="9577" lane="7" entrytime="00:01:04.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ML" nation="POL" region="LBL" clubid="7874" name="MASTERS Lublin">
          <CONTACT city="Lublin" email="masters_lublion@wp.pl" name="Wójcicki" phone="+48501794954" state="LUBEL" street="Stanisława Lema 18" zip="20-445" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-28" firstname="Anna" gender="F" lastname="Michalska" nation="POL" license="103503600002" athleteid="7886">
              <RESULTS>
                <RESULT eventid="1212" points="292" swimtime="00:03:10.00" resultid="7887" heatid="9338" lane="6" entrytime="00:03:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                    <SPLIT distance="100" swimtime="00:01:28.52" />
                    <SPLIT distance="150" swimtime="00:02:23.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="358" reactiontime="+75" swimtime="00:00:38.09" resultid="7888" heatid="9445" lane="1" entrytime="00:00:36.60" entrycourse="LCM" />
                <RESULT eventid="5348" points="355" reactiontime="+74" swimtime="00:01:22.01" resultid="7889" heatid="9532" lane="4" entrytime="00:01:21.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="318" reactiontime="+84" swimtime="00:03:01.66" resultid="7890" heatid="9581" lane="6" entrytime="00:03:02.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:01:27.09" />
                    <SPLIT distance="150" swimtime="00:02:15.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-07" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" license="103503700005" athleteid="7899">
              <RESULTS>
                <RESULT eventid="1544" points="385" swimtime="00:01:04.43" resultid="7900" heatid="9485" lane="1" entrytime="00:01:04.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="294" reactiontime="+92" swimtime="00:02:33.32" resultid="7901" heatid="9554" lane="7" entrytime="00:02:30.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="282" reactiontime="+86" swimtime="00:05:35.59" resultid="7902" heatid="9616" lane="3" entrytime="00:05:30.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:02:02.35" />
                    <SPLIT distance="200" swimtime="00:02:45.89" />
                    <SPLIT distance="250" swimtime="00:03:29.76" />
                    <SPLIT distance="300" swimtime="00:04:13.99" />
                    <SPLIT distance="350" swimtime="00:04:57.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-26" firstname="Rafał" gender="M" lastname="Zielonka" nation="POL" license="103503700008" athleteid="7891">
              <RESULTS>
                <RESULT eventid="1195" points="525" reactiontime="+80" swimtime="00:00:25.91" resultid="7892" heatid="9331" lane="5" entrytime="00:00:24.94" entrycourse="LCM" />
                <RESULT eventid="1280" points="414" reactiontime="+77" swimtime="00:10:06.21" resultid="7893" heatid="9359" lane="2" entrytime="00:10:05.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:44.68" />
                    <SPLIT distance="200" swimtime="00:02:22.14" />
                    <SPLIT distance="250" swimtime="00:02:59.95" />
                    <SPLIT distance="300" swimtime="00:03:38.30" />
                    <SPLIT distance="350" swimtime="00:04:16.75" />
                    <SPLIT distance="400" swimtime="00:04:55.27" />
                    <SPLIT distance="450" swimtime="00:05:33.86" />
                    <SPLIT distance="500" swimtime="00:06:12.95" />
                    <SPLIT distance="550" swimtime="00:06:51.94" />
                    <SPLIT distance="600" swimtime="00:07:31.01" />
                    <SPLIT distance="650" swimtime="00:08:10.19" />
                    <SPLIT distance="700" swimtime="00:08:49.02" />
                    <SPLIT distance="750" swimtime="00:09:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="563" reactiontime="+69" swimtime="00:00:56.79" resultid="7894" heatid="9489" lane="7" entrytime="00:00:57.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="532" reactiontime="+76" swimtime="00:00:27.67" resultid="7895" heatid="9527" lane="4" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="5399" points="496" reactiontime="+65" swimtime="00:02:08.84" resultid="7896" heatid="9558" lane="7" entrytime="00:02:07.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                    <SPLIT distance="150" swimtime="00:01:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="494" reactiontime="+76" swimtime="00:01:02.99" resultid="7897" heatid="9577" lane="3" entrytime="00:01:03.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="478" reactiontime="+69" swimtime="00:04:41.34" resultid="7898" heatid="9613" lane="7" entrytime="00:04:37.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:40.10" />
                    <SPLIT distance="200" swimtime="00:02:16.51" />
                    <SPLIT distance="250" swimtime="00:02:52.95" />
                    <SPLIT distance="300" swimtime="00:03:29.75" />
                    <SPLIT distance="350" swimtime="00:04:05.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-06" firstname="Marek" gender="M" lastname="Walencik" nation="POL" license="103503700010" athleteid="7903">
              <RESULTS>
                <RESULT eventid="1476" points="392" reactiontime="+81" swimtime="00:00:32.82" resultid="7904" heatid="9454" lane="3" entrytime="00:00:33.70" entrycourse="LCM" />
                <RESULT eventid="5297" points="394" reactiontime="+86" swimtime="00:01:17.90" resultid="7905" heatid="9511" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="361" reactiontime="+80" swimtime="00:01:12.76" resultid="7906" heatid="9540" lane="8" entrytime="00:01:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="443" reactiontime="+82" swimtime="00:00:34.03" resultid="7907" heatid="9603" lane="1" entrytime="00:00:34.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MO" nation="POL" region="MAL" clubid="6650" name="Masters Oświęcim">
          <CONTACT city="Oświęcim" email="js.formasy@interia.pl" name="Masters Oświęcim" phone="793691105" state="MAL" street="Tysiąclecia" zip="32-600" />
          <ATHLETES>
            <ATHLETE birthdate="1969-11-05" firstname="Sławomir" gender="M" lastname="Formas" nation="POL" athleteid="6655">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1510" points="522" swimtime="00:02:37.24" resultid="6656" heatid="9468" lane="6" entrytime="00:02:38.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5297" points="520" reactiontime="+73" swimtime="00:01:11.04" resultid="6657" heatid="9512" lane="4" entrytime="00:01:11.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="431" reactiontime="+80" swimtime="00:00:29.68" resultid="6658" heatid="9526" lane="3" entrytime="00:00:28.90" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5585" points="536" reactiontime="+72" swimtime="00:00:31.93" resultid="6659" heatid="9604" lane="2" entrytime="00:00:32.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-27" firstname="Robert" gender="M" lastname="Krulikowski" nation="POL" athleteid="6660">
              <RESULTS>
                <RESULT eventid="1476" points="304" reactiontime="+83" swimtime="00:00:35.72" resultid="6661" heatid="9453" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="5331" points="363" reactiontime="+94" swimtime="00:00:31.43" resultid="6662" heatid="9522" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="5365" points="286" reactiontime="+79" swimtime="00:01:18.69" resultid="6663" heatid="9539" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="250" reactiontime="+83" swimtime="00:02:57.62" resultid="6664" heatid="9587" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="150" swimtime="00:02:10.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="6651">
              <RESULTS>
                <RESULT eventid="1476" points="243" reactiontime="+78" swimtime="00:00:38.51" resultid="6652" heatid="9451" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="5365" points="233" reactiontime="+75" swimtime="00:01:24.25" resultid="6653" heatid="9537" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="212" reactiontime="+72" swimtime="00:03:07.59" resultid="6654" heatid="9586" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:28.46" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" athleteid="6671">
              <RESULTS>
                <RESULT eventid="1458" points="370" reactiontime="+83" swimtime="00:00:37.68" resultid="6672" heatid="9444" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="5348" points="310" reactiontime="+86" swimtime="00:01:25.83" resultid="6673" heatid="9531" lane="7" entrytime="00:01:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="277" reactiontime="+93" swimtime="00:03:10.19" resultid="6674" heatid="9581" lane="9" entrytime="00:03:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="100" swimtime="00:01:32.04" />
                    <SPLIT distance="150" swimtime="00:02:21.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" nation="POL" athleteid="6665">
              <RESULTS>
                <RESULT eventid="1458" points="209" reactiontime="+76" swimtime="00:00:45.54" resultid="6666" heatid="9442" lane="4" entrytime="00:00:43.30" />
                <RESULT eventid="1527" points="252" swimtime="00:01:21.82" resultid="6667" heatid="9473" lane="9" entrytime="00:01:18.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="248" reactiontime="+91" swimtime="00:01:41.96" resultid="6668" heatid="9502" lane="5" entrytime="00:01:38.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="233" reactiontime="+79" swimtime="00:03:03.56" resultid="6669" heatid="9545" lane="2" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                    <SPLIT distance="150" swimtime="00:02:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="253" reactiontime="+93" swimtime="00:00:46.43" resultid="6670" heatid="9594" lane="8" entrytime="00:00:44.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+82" swimtime="00:02:16.12" resultid="6675" heatid="9607" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:40.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6671" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="6655" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="6660" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="6665" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="5880" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="5901">
              <RESULTS>
                <RESULT eventid="1195" points="86" reactiontime="+130" swimtime="00:00:47.21" resultid="5902" heatid="9318" lane="8" entrytime="00:00:55.00" entrycourse="LCM" />
                <RESULT eventid="1229" points="51" reactiontime="+129" swimtime="00:05:05.87" resultid="5903" heatid="9342" lane="4" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="65" reactiontime="+99" swimtime="00:00:59.62" resultid="5904" heatid="9448" lane="7" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="78" reactiontime="+126" swimtime="00:01:49.67" resultid="5905" heatid="9478" lane="8" entrytime="00:01:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="67" reactiontime="+118" swimtime="00:02:20.53" resultid="5906" heatid="9506" lane="8" entrytime="00:02:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="5907" heatid="9549" lane="1" entrytime="00:04:10.00" entrycourse="LCM" />
                <RESULT eventid="5585" points="70" reactiontime="+130" swimtime="00:01:02.78" resultid="5908" heatid="9597" lane="2" entrytime="00:01:02.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-12" firstname="Janusz" gender="M" lastname="Mrozik" nation="POL" athleteid="5897">
              <RESULTS>
                <RESULT eventid="1510" points="55" reactiontime="+112" swimtime="00:05:31.73" resultid="5898" heatid="9462" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.92" />
                    <SPLIT distance="100" swimtime="00:02:43.41" />
                    <SPLIT distance="150" swimtime="00:04:10.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="45" reactiontime="+109" swimtime="00:02:40.08" resultid="5899" heatid="9505" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="52" reactiontime="+127" swimtime="00:04:32.86" resultid="5900" heatid="9548" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.44" />
                    <SPLIT distance="100" swimtime="00:02:11.03" />
                    <SPLIT distance="150" swimtime="00:03:21.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" license="501806600049" athleteid="5923">
              <RESULTS>
                <RESULT eventid="1133" points="556" reactiontime="+81" swimtime="00:00:28.78" resultid="5924" heatid="9315" lane="7" entrytime="00:00:28.21" entrycourse="LCM" />
                <RESULT eventid="1212" points="598" reactiontime="+81" swimtime="00:02:29.63" resultid="5925" heatid="9340" lane="5" entrytime="00:02:26.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                    <SPLIT distance="150" swimtime="00:01:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="506" reactiontime="+80" swimtime="00:02:54.52" resultid="5926" heatid="9461" lane="5" entrytime="00:02:46.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                    <SPLIT distance="150" swimtime="00:02:08.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="586" reactiontime="+77" swimtime="00:01:01.79" resultid="5927" heatid="9476" lane="3" entrytime="00:01:00.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="608" reactiontime="+74" swimtime="00:02:13.36" resultid="5928" heatid="9547" lane="4" entrytime="00:02:10.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="582" reactiontime="+79" swimtime="00:05:18.94" resultid="5929" heatid="9563" lane="4" entrytime="00:05:10.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:55.07" />
                    <SPLIT distance="200" swimtime="00:02:36.20" />
                    <SPLIT distance="250" swimtime="00:03:21.14" />
                    <SPLIT distance="300" swimtime="00:04:06.38" />
                    <SPLIT distance="350" swimtime="00:04:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="480" swimtime="00:01:10.84" resultid="5930" heatid="9571" lane="6" entrytime="00:01:10.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="550" reactiontime="+78" swimtime="00:00:35.88" resultid="5931" heatid="9596" lane="4" entrytime="00:00:35.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="5881">
              <RESULTS>
                <RESULT eventid="1212" points="89" reactiontime="+108" swimtime="00:04:42.43" resultid="5882" heatid="9337" lane="4" entrytime="00:04:34.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.63" />
                    <SPLIT distance="100" swimtime="00:02:13.99" />
                    <SPLIT distance="150" swimtime="00:03:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="102" swimtime="00:17:15.38" resultid="5883" heatid="9357" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.31" />
                    <SPLIT distance="100" swimtime="00:01:58.05" />
                    <SPLIT distance="150" swimtime="00:03:06.26" />
                    <SPLIT distance="200" swimtime="00:04:13.11" />
                    <SPLIT distance="250" swimtime="00:05:22.32" />
                    <SPLIT distance="300" swimtime="00:06:28.70" />
                    <SPLIT distance="350" swimtime="00:09:45.26" />
                    <SPLIT distance="400" swimtime="00:08:40.03" />
                    <SPLIT distance="450" swimtime="00:11:56.19" />
                    <SPLIT distance="500" swimtime="00:10:50.85" />
                    <SPLIT distance="550" swimtime="00:14:05.57" />
                    <SPLIT distance="600" swimtime="00:12:59.61" />
                    <SPLIT distance="650" swimtime="00:16:13.83" />
                    <SPLIT distance="700" swimtime="00:15:09.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="101" reactiontime="+78" swimtime="00:00:58.00" resultid="5884" heatid="9441" lane="6" entrytime="00:00:57.50" entrycourse="LCM" />
                <RESULT eventid="1527" points="108" swimtime="00:01:48.27" resultid="5885" heatid="9470" lane="6" entrytime="00:01:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="62" reactiontime="+103" swimtime="00:01:01.54" resultid="5886" heatid="9514" lane="1" entrytime="00:01:02.00" entrycourse="LCM" />
                <RESULT eventid="5348" points="90" reactiontime="+81" swimtime="00:02:09.26" resultid="5887" heatid="9530" lane="6" entrytime="00:02:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="69" swimtime="00:02:14.64" resultid="5888" heatid="9569" lane="6" entrytime="00:02:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="91" reactiontime="+85" swimtime="00:04:35.03" resultid="5889" heatid="9579" lane="4" entrytime="00:04:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.61" />
                    <SPLIT distance="100" swimtime="00:02:14.06" />
                    <SPLIT distance="150" swimtime="00:03:24.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzata" gender="F" lastname="Wach" nation="POL" athleteid="5918">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="5919" heatid="9311" lane="7" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1458" points="268" reactiontime="+61" swimtime="00:00:41.92" resultid="5920" heatid="9443" lane="1" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1527" points="256" swimtime="00:01:21.43" resultid="5921" heatid="9472" lane="6" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="240" reactiontime="+89" swimtime="00:03:01.59" resultid="5922" heatid="9545" lane="0" entrytime="00:02:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:14.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="5890">
              <RESULTS>
                <RESULT eventid="1476" points="74" reactiontime="+67" swimtime="00:00:57.23" resultid="5891" heatid="9448" lane="6" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="65" reactiontime="+104" swimtime="00:01:56.39" resultid="5892" heatid="9477" lane="5" entrytime="00:02:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="70" reactiontime="+74" swimtime="00:02:05.59" resultid="5893" heatid="9535" lane="0" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="61" reactiontime="+111" swimtime="00:04:17.72" resultid="5894" heatid="9549" lane="8" entrytime="00:04:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.18" />
                    <SPLIT distance="100" swimtime="00:02:04.62" />
                    <SPLIT distance="150" swimtime="00:03:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="5895" heatid="9584" lane="0" entrytime="00:04:58.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" license="501806600060" athleteid="5909">
              <RESULTS>
                <RESULT eventid="1133" points="91" reactiontime="+101" swimtime="00:00:52.53" resultid="5910" heatid="9309" lane="5" entrytime="00:00:49.06" entrycourse="LCM" />
                <RESULT eventid="1263" points="85" reactiontime="+118" swimtime="00:18:19.60" resultid="5911" heatid="9357" lane="3" entrytime="00:18:09.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.15" />
                    <SPLIT distance="100" swimtime="00:01:57.94" />
                    <SPLIT distance="150" swimtime="00:03:05.61" />
                    <SPLIT distance="200" swimtime="00:04:15.06" />
                    <SPLIT distance="250" swimtime="00:05:25.09" />
                    <SPLIT distance="300" swimtime="00:06:34.21" />
                    <SPLIT distance="350" swimtime="00:07:45.44" />
                    <SPLIT distance="400" swimtime="00:08:56.41" />
                    <SPLIT distance="450" swimtime="00:10:06.43" />
                    <SPLIT distance="500" swimtime="00:11:17.13" />
                    <SPLIT distance="550" swimtime="00:12:28.43" />
                    <SPLIT distance="600" swimtime="00:13:39.37" />
                    <SPLIT distance="650" swimtime="00:14:49.59" />
                    <SPLIT distance="700" swimtime="00:15:59.69" />
                    <SPLIT distance="750" swimtime="00:17:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="84" reactiontime="+98" swimtime="00:01:01.76" resultid="5912" heatid="9441" lane="9" entrytime="00:01:04.00" entrycourse="LCM" />
                <RESULT eventid="1527" points="83" reactiontime="+107" swimtime="00:01:58.29" resultid="5913" heatid="9470" lane="7" entrytime="00:01:54.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="56" swimtime="00:01:03.51" resultid="5914" heatid="9514" lane="8" entrytime="00:01:03.23" entrycourse="LCM" />
                <RESULT eventid="5382" points="91" reactiontime="+129" swimtime="00:04:11.03" resultid="5915" heatid="9542" lane="5" entrytime="00:04:04.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:02:00.89" />
                    <SPLIT distance="150" swimtime="00:03:07.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="49" reactiontime="+121" swimtime="00:02:31.26" resultid="5916" heatid="9569" lane="2" entrytime="00:02:23.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="94" swimtime="00:08:38.70" resultid="5917" heatid="9612" lane="7" entrytime="00:08:53.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                    <SPLIT distance="100" swimtime="00:01:56.41" />
                    <SPLIT distance="150" swimtime="00:03:02.64" />
                    <SPLIT distance="200" swimtime="00:04:09.50" />
                    <SPLIT distance="250" swimtime="00:05:16.66" />
                    <SPLIT distance="300" swimtime="00:06:25.62" />
                    <SPLIT distance="350" swimtime="00:07:32.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MZ" nation="POL" clubid="8321" name="MASTERS Zdzieszowice">
          <CONTACT email="dejot.swim@gmail.com" name="Jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1988-03-21" firstname="Szymon" gender="M" lastname="Paciej" nation="POL" athleteid="8322">
              <RESULTS>
                <RESULT eventid="1476" points="404" reactiontime="+91" swimtime="00:00:32.50" resultid="8323" heatid="9455" lane="9" entrytime="00:00:33.20" />
                <RESULT eventid="1510" points="379" swimtime="00:02:54.92" resultid="8324" heatid="9467" lane="1" entrytime="00:02:55.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="399" reactiontime="+81" swimtime="00:01:10.41" resultid="8325" heatid="9540" lane="1" entrytime="00:01:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="323" reactiontime="+84" swimtime="00:05:55.10" resultid="8326" heatid="9567" lane="7" entrytime="00:05:45.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:09.97" />
                    <SPLIT distance="200" swimtime="00:02:54.55" />
                    <SPLIT distance="250" swimtime="00:03:44.29" />
                    <SPLIT distance="300" swimtime="00:04:34.22" />
                    <SPLIT distance="350" swimtime="00:05:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="382" reactiontime="+96" swimtime="00:02:34.15" resultid="8327" heatid="9589" lane="6" entrytime="00:02:35.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-08" firstname="Sasha" gender="M" lastname="Broshevan" nation="POL" athleteid="8337">
              <RESULTS>
                <RESULT eventid="1195" points="396" reactiontime="+92" swimtime="00:00:28.47" resultid="8338" heatid="9317" lane="6" />
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /G8" eventid="1229" status="DSQ" swimtime="00:02:53.69" resultid="8339" heatid="9346" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:02:15.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="315" reactiontime="+72" swimtime="00:00:35.31" resultid="8340" heatid="9452" lane="3" entrytime="00:00:37.65" />
                <RESULT eventid="1544" points="382" reactiontime="+78" swimtime="00:01:04.65" resultid="8341" heatid="9485" lane="8" entrytime="00:01:04.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="376" reactiontime="+78" swimtime="00:00:31.06" resultid="8342" heatid="9518" lane="2" />
                <RESULT eventid="5365" points="276" reactiontime="+75" swimtime="00:01:19.59" resultid="8343" heatid="9537" lane="4" entrytime="00:01:20.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="231" reactiontime="+98" swimtime="00:03:02.26" resultid="8344" heatid="9583" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="321" reactiontime="+85" swimtime="00:00:37.89" resultid="8345" heatid="9600" lane="4" entrytime="00:00:38.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-04" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="8346">
              <RESULTS>
                <RESULT eventid="1493" points="248" reactiontime="+97" swimtime="00:03:41.39" resultid="8347" heatid="9459" lane="4" entrytime="00:03:33.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                    <SPLIT distance="100" swimtime="00:01:42.51" />
                    <SPLIT distance="150" swimtime="00:02:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="261" reactiontime="+82" swimtime="00:01:20.86" resultid="8348" heatid="9472" lane="7" entrytime="00:01:22.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="278" swimtime="00:01:38.22" resultid="8349" heatid="9502" lane="7" entrytime="00:01:41.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" reactiontime="+88" status="DNS" swimtime="00:00:00.00" resultid="8350" heatid="9563" lane="0" entrytime="00:06:55.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="272" reactiontime="+92" swimtime="00:00:45.36" resultid="8351" heatid="9593" lane="3" entrytime="00:00:45.65" />
                <RESULT eventid="5619" points="209" reactiontime="+99" swimtime="00:06:38.35" resultid="8352" heatid="9611" lane="5" entrytime="00:06:40.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                    <SPLIT distance="200" swimtime="00:03:12.53" />
                    <SPLIT distance="250" swimtime="00:04:04.54" />
                    <SPLIT distance="300" swimtime="00:04:56.77" />
                    <SPLIT distance="350" swimtime="00:05:49.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-05" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="8353">
              <RESULTS>
                <RESULT eventid="1458" points="300" reactiontime="+75" swimtime="00:00:40.38" resultid="8354" heatid="9444" lane="1" entrytime="00:00:39.65" />
                <RESULT eventid="1561" points="220" reactiontime="+104" swimtime="00:03:21.76" resultid="8355" heatid="9492" lane="2" entrytime="00:03:14.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                    <SPLIT distance="150" swimtime="00:02:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="317" reactiontime="+82" swimtime="00:01:25.18" resultid="8356" heatid="9532" lane="7" entrytime="00:01:25.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="274" swimtime="00:06:49.72" resultid="8357" heatid="9563" lane="7" entrytime="00:06:20.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:34.66" />
                    <SPLIT distance="150" swimtime="00:02:28.48" />
                    <SPLIT distance="200" swimtime="00:03:20.65" />
                    <SPLIT distance="250" swimtime="00:04:19.51" />
                    <SPLIT distance="300" swimtime="00:05:18.23" />
                    <SPLIT distance="350" swimtime="00:06:02.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="299" reactiontime="+75" swimtime="00:03:05.39" resultid="8358" heatid="9581" lane="3" entrytime="00:03:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                    <SPLIT distance="150" swimtime="00:02:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="255" reactiontime="+97" swimtime="00:06:12.76" resultid="8359" heatid="9610" lane="7" entrytime="00:06:05.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                    <SPLIT distance="200" swimtime="00:03:01.91" />
                    <SPLIT distance="250" swimtime="00:03:49.77" />
                    <SPLIT distance="300" swimtime="00:04:37.79" />
                    <SPLIT distance="350" swimtime="00:05:25.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="8328">
              <RESULTS>
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="8329" heatid="9349" lane="1" entrytime="00:02:24.34" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="8331" heatid="9490" lane="9" entrytime="00:00:56.02" />
                <RESULT eventid="1578" points="440" reactiontime="+76" swimtime="00:02:26.59" resultid="8332" heatid="9496" lane="8" entrytime="00:02:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="150" swimtime="00:01:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="470" reactiontime="+73" swimtime="00:01:13.43" resultid="8333" heatid="9512" lane="5" entrytime="00:01:12.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="434" swimtime="00:05:21.93" resultid="8334" heatid="9568" lane="9" entrytime="00:05:15.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                    <SPLIT distance="200" swimtime="00:02:35.97" />
                    <SPLIT distance="250" swimtime="00:03:20.48" />
                    <SPLIT distance="300" swimtime="00:04:06.86" />
                    <SPLIT distance="350" swimtime="00:04:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="514" swimtime="00:01:02.18" resultid="8335" heatid="9578" lane="9" entrytime="00:01:02.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="517" reactiontime="+79" swimtime="00:00:32.33" resultid="8336" heatid="9604" lane="6" entrytime="00:00:32.23" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+79" swimtime="00:02:19.83" resultid="8360" heatid="9608" lane="9" entrytime="00:02:20.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8353" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="8322" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="8346" number="3" />
                    <RELAYPOSITION athleteid="8328" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ML" nation="POL" clubid="6676" name="MASTERS Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" license="103605700004" athleteid="6677">
              <RESULTS>
                <RESULT eventid="1195" points="364" reactiontime="+101" swimtime="00:00:29.26" resultid="6678" heatid="9319" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1229" points="254" reactiontime="+93" swimtime="00:02:59.91" resultid="6679" heatid="9344" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:16.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="276" reactiontime="+90" swimtime="00:00:36.92" resultid="6680" heatid="9450" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1510" points="264" reactiontime="+97" swimtime="00:03:17.32" resultid="6681" heatid="9463" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="100" swimtime="00:01:31.74" />
                    <SPLIT distance="150" swimtime="00:02:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="224" reactiontime="+91" swimtime="00:01:25.27" resultid="6682" heatid="9536" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="168" reactiontime="+107" swimtime="00:07:21.28" resultid="6683" heatid="9564" lane="3" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:31.34" />
                    <SPLIT distance="150" swimtime="00:02:33.18" />
                    <SPLIT distance="200" swimtime="00:03:32.05" />
                    <SPLIT distance="250" swimtime="00:04:35.24" />
                    <SPLIT distance="300" swimtime="00:05:38.69" />
                    <SPLIT distance="350" swimtime="00:06:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="206" reactiontime="+85" swimtime="00:03:09.43" resultid="6684" heatid="9585" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="150" swimtime="00:02:18.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="285" reactiontime="+96" swimtime="00:00:39.43" resultid="6685" heatid="9598" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASTKRAS" nation="POL" region="LBL" clubid="6582" name="Masterskrasnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" name="Michalczyk Jerzy" phone="601 69 89 77" state="LUB" street="Żwirki i Wigury 2" zip="23-204" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-04" firstname="Mirisław" gender="M" lastname="Leszczyński" nation="POL" athleteid="6597">
              <RESULTS>
                <RESULT eventid="1510" points="285" swimtime="00:03:12.34" resultid="6598" heatid="9465" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                    <SPLIT distance="150" swimtime="00:02:23.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="275" reactiontime="+94" swimtime="00:01:27.83" resultid="6599" heatid="9508" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="289" reactiontime="+101" swimtime="00:00:39.24" resultid="6600" heatid="9600" lane="8" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="6583">
              <RESULTS>
                <RESULT eventid="1314" reactiontime="+127" status="OTL" swimtime="00:00:00.00" resultid="6584" heatid="9368" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.87" />
                    <SPLIT distance="100" swimtime="00:02:08.68" />
                    <SPLIT distance="150" swimtime="00:03:19.62" />
                    <SPLIT distance="200" swimtime="00:04:29.81" />
                    <SPLIT distance="250" swimtime="00:05:45.80" />
                    <SPLIT distance="300" swimtime="00:06:56.09" />
                    <SPLIT distance="350" swimtime="00:08:11.54" />
                    <SPLIT distance="400" swimtime="00:09:22.35" />
                    <SPLIT distance="450" swimtime="00:10:37.91" />
                    <SPLIT distance="500" swimtime="00:11:47.75" />
                    <SPLIT distance="550" swimtime="00:13:03.03" />
                    <SPLIT distance="600" swimtime="00:14:15.04" />
                    <SPLIT distance="650" swimtime="00:15:28.81" />
                    <SPLIT distance="700" swimtime="00:16:42.66" />
                    <SPLIT distance="750" swimtime="00:17:56.30" />
                    <SPLIT distance="800" swimtime="00:19:05.64" />
                    <SPLIT distance="850" swimtime="00:20:17.92" />
                    <SPLIT distance="900" swimtime="00:21:27.84" />
                    <SPLIT distance="950" swimtime="00:22:39.84" />
                    <SPLIT distance="1000" swimtime="00:23:51.24" />
                    <SPLIT distance="1050" swimtime="00:24:58.83" />
                    <SPLIT distance="1100" swimtime="00:26:06.91" />
                    <SPLIT distance="1150" swimtime="00:27:18.55" />
                    <SPLIT distance="1200" swimtime="00:28:29.61" />
                    <SPLIT distance="1250" swimtime="00:29:40.85" />
                    <SPLIT distance="1300" swimtime="00:30:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="126" swimtime="00:04:12.58" resultid="6585" heatid="9463" lane="1" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.63" />
                    <SPLIT distance="100" swimtime="00:02:00.21" />
                    <SPLIT distance="150" swimtime="00:03:09.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="53" swimtime="00:04:56.82" resultid="6586" heatid="9493" lane="6" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.45" />
                    <SPLIT distance="100" swimtime="00:02:10.12" />
                    <SPLIT distance="150" swimtime="00:03:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="116" reactiontime="+162" swimtime="00:01:56.83" resultid="6587" heatid="9506" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="6591">
              <RESULTS>
                <RESULT eventid="1195" points="120" reactiontime="+101" swimtime="00:00:42.35" resultid="6592" heatid="9318" lane="7" entrytime="00:00:49.30" />
                <RESULT eventid="1476" points="86" reactiontime="+84" swimtime="00:00:54.28" resultid="6593" heatid="9448" lane="1" entrytime="00:01:02.25" />
                <RESULT eventid="1544" points="97" reactiontime="+94" swimtime="00:01:41.85" resultid="6594" heatid="9478" lane="0" entrytime="00:01:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="67" reactiontime="+93" swimtime="00:00:55.20" resultid="6595" heatid="9519" lane="0" entrytime="00:00:55.25" />
                <RESULT eventid="5517" points="56" reactiontime="+94" swimtime="00:02:09.98" resultid="6596" heatid="9572" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="6607">
              <RESULTS>
                <RESULT eventid="1229" points="163" reactiontime="+79" swimtime="00:03:28.41" resultid="6608" heatid="9345" lane="8" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="100" swimtime="00:01:36.85" />
                    <SPLIT distance="150" swimtime="00:02:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="6610" heatid="9452" lane="8" entrytime="00:00:39.10" />
                <RESULT eventid="1578" points="71" reactiontime="+88" swimtime="00:04:28.63" resultid="6611" heatid="9493" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.88" />
                    <SPLIT distance="100" swimtime="00:02:01.06" />
                    <SPLIT distance="150" swimtime="00:03:14.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6612" heatid="9536" lane="2" entrytime="00:01:36.10" />
                <RESULT eventid="5467" points="125" swimtime="00:08:07.60" resultid="6613" heatid="9565" lane="7" entrytime="00:07:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.71" />
                    <SPLIT distance="100" swimtime="00:02:13.73" />
                    <SPLIT distance="150" swimtime="00:03:18.53" />
                    <SPLIT distance="200" swimtime="00:04:24.26" />
                    <SPLIT distance="250" swimtime="00:05:31.79" />
                    <SPLIT distance="300" swimtime="00:06:36.31" />
                    <SPLIT distance="350" swimtime="00:07:26.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6614" heatid="9586" lane="0" entrytime="00:03:21.10" />
                <RESULT eventid="5636" points="157" reactiontime="+74" swimtime="00:06:47.60" resultid="6615" heatid="9617" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:34.50" />
                    <SPLIT distance="150" swimtime="00:02:26.80" />
                    <SPLIT distance="200" swimtime="00:03:22.24" />
                    <SPLIT distance="250" swimtime="00:04:15.65" />
                    <SPLIT distance="300" swimtime="00:05:09.60" />
                    <SPLIT distance="350" swimtime="00:06:01.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-17" firstname="Jacek" gender="M" lastname="Janik" nation="POL" athleteid="6601">
              <RESULTS>
                <RESULT eventid="1195" points="174" reactiontime="+102" swimtime="00:00:37.39" resultid="6602" heatid="9320" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1544" points="153" reactiontime="+98" swimtime="00:01:27.70" resultid="6603" heatid="9480" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="146" reactiontime="+102" swimtime="00:01:48.37" resultid="6604" heatid="9506" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="6605" heatid="9551" lane="9" entrytime="00:03:15.00" />
                <RESULT eventid="5585" points="173" reactiontime="+98" swimtime="00:00:46.55" resultid="6606" heatid="9598" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MUK" nation="EST" clubid="8214" name="Meisterujumise U-Klubi">
          <CONTACT email="a_kristiina@hotmail.com" name="Kristiina Arusoo" phone="+37256656831" />
          <ATHLETES>
            <ATHLETE birthdate="1954-08-05" firstname="Ossi Albin" gender="M" lastname="Vallemaa" nation="FIN" athleteid="8240">
              <RESULTS>
                <RESULT eventid="1510" status="DNS" swimtime="00:00:00.00" resultid="8241" heatid="9463" lane="3" entrytime="00:03:42.99" entrycourse="LCM" />
                <RESULT eventid="5297" points="186" reactiontime="+70" swimtime="00:01:39.92" resultid="8242" heatid="9507" lane="3" entrytime="00:01:36.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" status="DNS" swimtime="00:00:00.00" resultid="8243" heatid="9599" lane="6" entrytime="00:00:41.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="SZ" clubid="6786" name="MKP Szczecin">
          <CONTACT name="Kowalczyk" />
          <ATHLETES>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="6800">
              <RESULTS>
                <RESULT eventid="1314" points="356" swimtime="00:20:28.11" resultid="6801" heatid="9365" lane="1" entrytime="00:20:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                    <SPLIT distance="200" swimtime="00:02:34.29" />
                    <SPLIT distance="250" swimtime="00:03:14.11" />
                    <SPLIT distance="300" swimtime="00:03:55.14" />
                    <SPLIT distance="350" swimtime="00:04:35.57" />
                    <SPLIT distance="400" swimtime="00:05:16.38" />
                    <SPLIT distance="450" swimtime="00:05:57.08" />
                    <SPLIT distance="500" swimtime="00:06:37.99" />
                    <SPLIT distance="550" swimtime="00:07:18.96" />
                    <SPLIT distance="600" swimtime="00:08:00.47" />
                    <SPLIT distance="650" swimtime="00:08:41.95" />
                    <SPLIT distance="700" swimtime="00:09:24.01" />
                    <SPLIT distance="750" swimtime="00:10:05.73" />
                    <SPLIT distance="800" swimtime="00:10:47.67" />
                    <SPLIT distance="850" swimtime="00:11:29.36" />
                    <SPLIT distance="900" swimtime="00:12:11.22" />
                    <SPLIT distance="950" swimtime="00:12:53.60" />
                    <SPLIT distance="1000" swimtime="00:13:34.53" />
                    <SPLIT distance="1050" swimtime="00:14:16.83" />
                    <SPLIT distance="1100" swimtime="00:14:58.57" />
                    <SPLIT distance="1150" swimtime="00:15:40.40" />
                    <SPLIT distance="1200" swimtime="00:16:21.94" />
                    <SPLIT distance="1250" swimtime="00:17:03.83" />
                    <SPLIT distance="1300" swimtime="00:17:45.30" />
                    <SPLIT distance="1350" swimtime="00:18:26.84" />
                    <SPLIT distance="1400" swimtime="00:19:09.03" />
                    <SPLIT distance="1450" swimtime="00:19:50.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="279" reactiontime="+82" swimtime="00:00:36.77" resultid="6802" heatid="9453" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1544" points="395" reactiontime="+83" swimtime="00:01:03.89" resultid="6803" heatid="9485" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6804" heatid="9538" lane="2" entrytime="00:01:18.00" />
                <RESULT eventid="5399" points="352" reactiontime="+83" swimtime="00:02:24.34" resultid="6805" heatid="9556" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="307" reactiontime="+79" swimtime="00:02:45.86" resultid="6806" heatid="9589" lane="9" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="6838">
              <RESULTS>
                <RESULT eventid="1458" points="37" reactiontime="+101" swimtime="00:01:21.07" resultid="6839" heatid="9440" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1493" points="76" swimtime="00:05:27.22" resultid="6840" heatid="9458" lane="2" entrytime="00:05:06.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.60" />
                    <SPLIT distance="100" swimtime="00:02:40.88" />
                    <SPLIT distance="150" swimtime="00:04:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="73" swimtime="00:02:33.23" resultid="6841" heatid="9500" lane="5" entrytime="00:02:25.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="68" swimtime="00:01:11.83" resultid="6842" heatid="9592" lane="0" entrytime="00:01:09.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-31" firstname="Konrad" gender="M" lastname="Tekiel" nation="POL" athleteid="6849">
              <RESULTS>
                <RESULT eventid="1280" status="OTL" swimtime="00:13:41.15" resultid="6850" heatid="9361" lane="9" entrytime="00:13:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:21.76" />
                    <SPLIT distance="200" swimtime="00:03:14.14" />
                    <SPLIT distance="250" swimtime="00:04:07.17" />
                    <SPLIT distance="300" swimtime="00:04:59.93" />
                    <SPLIT distance="350" swimtime="00:05:51.67" />
                    <SPLIT distance="400" swimtime="00:06:44.24" />
                    <SPLIT distance="450" swimtime="00:07:36.49" />
                    <SPLIT distance="500" swimtime="00:08:28.99" />
                    <SPLIT distance="550" swimtime="00:09:21.25" />
                    <SPLIT distance="600" swimtime="00:10:14.87" />
                    <SPLIT distance="650" swimtime="00:11:07.66" />
                    <SPLIT distance="700" swimtime="00:12:00.09" />
                    <SPLIT distance="750" swimtime="00:12:52.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="175" reactiontime="+81" swimtime="00:01:23.83" resultid="6851" heatid="9479" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="6843">
              <RESULTS>
                <RESULT comment="Czas Lepszy od rekordu Polski Kat F" eventid="1263" points="434" reactiontime="+80" swimtime="00:10:40.15" resultid="6844" heatid="9355" lane="2" entrytime="00:10:50.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:53.84" />
                    <SPLIT distance="200" swimtime="00:02:33.92" />
                    <SPLIT distance="250" swimtime="00:03:14.07" />
                    <SPLIT distance="300" swimtime="00:03:54.42" />
                    <SPLIT distance="350" swimtime="00:04:34.92" />
                    <SPLIT distance="400" swimtime="00:05:15.51" />
                    <SPLIT distance="450" swimtime="00:05:56.06" />
                    <SPLIT distance="500" swimtime="00:06:36.72" />
                    <SPLIT distance="550" swimtime="00:07:17.32" />
                    <SPLIT distance="600" swimtime="00:07:58.02" />
                    <SPLIT distance="650" swimtime="00:08:38.99" />
                    <SPLIT distance="700" swimtime="00:09:20.01" />
                    <SPLIT distance="750" swimtime="00:10:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="405" reactiontime="+83" swimtime="00:01:09.84" resultid="6845" heatid="9474" lane="3" entrytime="00:01:11.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="426" reactiontime="+82" swimtime="00:02:30.08" resultid="6846" heatid="9547" lane="0" entrytime="00:02:30.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="302" reactiontime="+79" swimtime="00:03:04.83" resultid="6847" heatid="9582" lane="8" entrytime="00:02:58.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5619" points="422" reactiontime="+82" swimtime="00:05:15.11" resultid="6848" heatid="9609" lane="7" entrytime="00:05:23.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:55.27" />
                    <SPLIT distance="200" swimtime="00:02:35.61" />
                    <SPLIT distance="250" swimtime="00:03:15.41" />
                    <SPLIT distance="300" swimtime="00:03:55.73" />
                    <SPLIT distance="350" swimtime="00:04:35.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="6829">
              <RESULTS>
                <RESULT eventid="1195" points="270" reactiontime="+69" swimtime="00:00:32.34" resultid="6830" heatid="9322" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1314" points="234" swimtime="00:23:31.54" resultid="6831" heatid="9366" lane="1" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:02:15.62" />
                    <SPLIT distance="200" swimtime="00:03:04.11" />
                    <SPLIT distance="250" swimtime="00:03:53.72" />
                    <SPLIT distance="300" swimtime="00:04:42.82" />
                    <SPLIT distance="350" swimtime="00:05:31.69" />
                    <SPLIT distance="400" swimtime="00:06:19.83" />
                    <SPLIT distance="450" swimtime="00:07:06.51" />
                    <SPLIT distance="500" swimtime="00:07:54.88" />
                    <SPLIT distance="550" swimtime="00:08:43.62" />
                    <SPLIT distance="600" swimtime="00:09:30.83" />
                    <SPLIT distance="650" swimtime="00:10:18.77" />
                    <SPLIT distance="700" swimtime="00:11:05.76" />
                    <SPLIT distance="750" swimtime="00:11:53.26" />
                    <SPLIT distance="800" swimtime="00:12:41.45" />
                    <SPLIT distance="850" swimtime="00:13:29.97" />
                    <SPLIT distance="900" swimtime="00:14:17.25" />
                    <SPLIT distance="950" swimtime="00:15:05.26" />
                    <SPLIT distance="1000" swimtime="00:15:52.90" />
                    <SPLIT distance="1050" swimtime="00:16:39.80" />
                    <SPLIT distance="1100" swimtime="00:17:26.33" />
                    <SPLIT distance="1150" swimtime="00:18:12.24" />
                    <SPLIT distance="1200" swimtime="00:18:58.76" />
                    <SPLIT distance="1250" swimtime="00:19:44.72" />
                    <SPLIT distance="1300" swimtime="00:20:31.07" />
                    <SPLIT distance="1350" swimtime="00:21:17.14" />
                    <SPLIT distance="1400" swimtime="00:22:02.54" />
                    <SPLIT distance="1450" swimtime="00:22:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="6832" heatid="9452" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1544" points="295" reactiontime="+87" swimtime="00:01:10.44" resultid="6833" heatid="9483" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6834" heatid="9537" lane="7" entrytime="00:01:25.00" />
                <RESULT eventid="5399" points="271" reactiontime="+87" swimtime="00:02:37.54" resultid="6835" heatid="9553" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:01:58.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6836" heatid="9586" lane="3" entrytime="00:03:10.00" />
                <RESULT eventid="5636" points="251" reactiontime="+97" swimtime="00:05:48.75" resultid="6837" heatid="9616" lane="8" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:07.59" />
                    <SPLIT distance="200" swimtime="00:02:53.71" />
                    <SPLIT distance="250" swimtime="00:03:38.96" />
                    <SPLIT distance="300" swimtime="00:04:23.75" />
                    <SPLIT distance="350" swimtime="00:05:08.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="6813">
              <RESULTS>
                <RESULT eventid="1458" points="271" reactiontime="+101" swimtime="00:00:41.81" resultid="6814" heatid="9443" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1527" points="251" reactiontime="+109" swimtime="00:01:21.93" resultid="6815" heatid="9472" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="274" reactiontime="+88" swimtime="00:01:29.40" resultid="6816" heatid="9531" lane="5" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5382" points="260" reactiontime="+110" swimtime="00:02:56.98" resultid="6817" heatid="9544" lane="3" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:02:10.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5534" points="273" reactiontime="+90" swimtime="00:03:11.01" resultid="6818" heatid="9581" lane="8" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                    <SPLIT distance="150" swimtime="00:02:20.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="242" reactiontime="+112" swimtime="00:06:19.32" resultid="6819" heatid="9611" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:01:27.19" />
                    <SPLIT distance="150" swimtime="00:02:14.46" />
                    <SPLIT distance="200" swimtime="00:03:03.19" />
                    <SPLIT distance="250" swimtime="00:03:52.03" />
                    <SPLIT distance="300" swimtime="00:04:42.13" />
                    <SPLIT distance="350" swimtime="00:05:31.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="6808">
              <RESULTS>
                <RESULT eventid="1229" points="179" reactiontime="+75" swimtime="00:03:22.14" resultid="6809" heatid="9343" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:36.08" />
                    <SPLIT distance="150" swimtime="00:02:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="201" reactiontime="+79" swimtime="00:03:36.10" resultid="6810" heatid="9463" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="100" swimtime="00:01:44.75" />
                    <SPLIT distance="150" swimtime="00:02:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="202" reactiontime="+75" swimtime="00:01:37.24" resultid="6811" heatid="9507" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="260" reactiontime="+83" swimtime="00:00:40.62" resultid="6812" heatid="9599" lane="8" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="6820">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1229" reactiontime="+65" status="DSQ" swimtime="00:03:07.25" resultid="6821" heatid="9344" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="150" swimtime="00:02:20.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="174" reactiontime="+96" swimtime="00:13:29.72" resultid="6822" heatid="9361" lane="2" entrytime="00:12:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:28.94" />
                    <SPLIT distance="150" swimtime="00:02:19.11" />
                    <SPLIT distance="200" swimtime="00:03:09.62" />
                    <SPLIT distance="250" swimtime="00:04:01.13" />
                    <SPLIT distance="300" swimtime="00:04:52.64" />
                    <SPLIT distance="350" swimtime="00:05:43.30" />
                    <SPLIT distance="400" swimtime="00:06:34.09" />
                    <SPLIT distance="450" swimtime="00:07:25.26" />
                    <SPLIT distance="500" swimtime="00:08:16.75" />
                    <SPLIT distance="550" swimtime="00:09:08.88" />
                    <SPLIT distance="600" swimtime="00:10:01.09" />
                    <SPLIT distance="650" swimtime="00:10:53.68" />
                    <SPLIT distance="700" swimtime="00:11:46.78" />
                    <SPLIT distance="750" swimtime="00:12:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="226" reactiontime="+105" swimtime="00:03:27.65" resultid="6824" heatid="9464" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="224" reactiontime="+95" swimtime="00:01:33.99" resultid="6825" heatid="9509" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="192" reactiontime="+103" swimtime="00:01:26.30" resultid="6827" heatid="9574" lane="8" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6828" heatid="9586" lane="1" entrytime="00:03:13.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="ZAC" clubid="7685" name="MKS Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1994-09-30" firstname="Mateusz" gender="M" lastname="Drozd" nation="POL" athleteid="7700">
              <RESULTS>
                <RESULT eventid="1195" points="576" reactiontime="+71" swimtime="00:00:25.13" resultid="7701" heatid="9332" lane="0" entrytime="00:00:24.73" />
                <RESULT eventid="1229" points="507" reactiontime="+70" swimtime="00:02:22.88" resultid="7702" heatid="9349" lane="5" entrytime="00:02:12.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="429" swimtime="00:02:27.80" resultid="7703" heatid="9496" lane="6" entrytime="00:02:18.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:03.51" />
                    <SPLIT distance="150" swimtime="00:01:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="584" reactiontime="+71" swimtime="00:02:02.01" resultid="7704" heatid="9558" lane="4" entrytime="00:01:56.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:00:59.32" />
                    <SPLIT distance="150" swimtime="00:01:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="470" reactiontime="+73" swimtime="00:05:13.58" resultid="7705" heatid="9568" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:48.82" />
                    <SPLIT distance="200" swimtime="00:02:29.29" />
                    <SPLIT distance="250" swimtime="00:03:13.63" />
                    <SPLIT distance="300" swimtime="00:04:00.82" />
                    <SPLIT distance="350" swimtime="00:04:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="514" reactiontime="+68" swimtime="00:01:02.19" resultid="7706" heatid="9578" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="456" reactiontime="+76" swimtime="00:00:33.70" resultid="7707" heatid="9604" lane="9" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-20" firstname="Mariusz" gender="M" lastname="Chrzan" nation="POL" athleteid="7693">
              <RESULTS>
                <RESULT eventid="1229" points="424" swimtime="00:02:31.74" resultid="7694" heatid="9349" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:09.14" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="463" reactiontime="+86" swimtime="00:00:31.06" resultid="7695" heatid="9456" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1544" points="487" reactiontime="+70" swimtime="00:00:59.61" resultid="7696" heatid="9489" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="456" reactiontime="+76" swimtime="00:01:07.33" resultid="7697" heatid="9541" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="391" reactiontime="+68" swimtime="00:05:33.32" resultid="7698" heatid="9568" lane="7" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                    <SPLIT distance="200" swimtime="00:02:35.99" />
                    <SPLIT distance="250" swimtime="00:03:25.29" />
                    <SPLIT distance="300" swimtime="00:04:16.52" />
                    <SPLIT distance="350" swimtime="00:04:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="422" reactiontime="+75" swimtime="00:02:29.12" resultid="7699" heatid="9590" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:50.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSIR" nation="POL" clubid="6072" name="MOSiR Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="6073">
              <RESULTS>
                <RESULT eventid="1195" points="249" reactiontime="+92" swimtime="00:00:33.21" resultid="6074" heatid="9321" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1229" points="143" reactiontime="+97" swimtime="00:03:37.78" resultid="6075" heatid="9343" lane="3" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:43.16" />
                    <SPLIT distance="150" swimtime="00:02:49.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="210" swimtime="00:01:18.82" resultid="6076" heatid="9481" lane="1" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="82" reactiontime="+99" swimtime="00:04:16.38" resultid="6077" heatid="9493" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.14" />
                    <SPLIT distance="150" swimtime="00:03:12.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="220" reactiontime="+101" swimtime="00:00:37.13" resultid="6078" heatid="9521" lane="8" entrytime="00:00:36.90" />
                <RESULT eventid="5467" points="116" reactiontime="+98" swimtime="00:08:19.88" resultid="6079" heatid="9565" lane="8" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.98" />
                    <SPLIT distance="100" swimtime="00:02:07.17" />
                    <SPLIT distance="150" swimtime="00:03:16.80" />
                    <SPLIT distance="200" swimtime="00:04:23.50" />
                    <SPLIT distance="250" swimtime="00:05:33.28" />
                    <SPLIT distance="300" swimtime="00:06:41.38" />
                    <SPLIT distance="350" swimtime="00:07:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="120" swimtime="00:01:40.79" resultid="6080" heatid="9573" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="132" reactiontime="+95" swimtime="00:07:11.27" resultid="6081" heatid="9618" lane="8" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:36.62" />
                    <SPLIT distance="150" swimtime="00:02:31.51" />
                    <SPLIT distance="200" swimtime="00:03:29.12" />
                    <SPLIT distance="250" swimtime="00:04:25.18" />
                    <SPLIT distance="300" swimtime="00:05:22.20" />
                    <SPLIT distance="350" swimtime="00:06:18.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" clubid="6532" name="MOTYL Senior MOSiR Stalowa Wola" shortname="MOTYL Senior MOSiR Stalowa Wol">
          <CONTACT name="Berwecki" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="6533">
              <RESULTS>
                <RESULT eventid="1229" points="509" reactiontime="+68" swimtime="00:02:22.72" resultid="6534" heatid="9349" lane="7" entrytime="00:02:23.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1578" points="459" swimtime="00:02:24.55" resultid="6535" heatid="9496" lane="1" entrytime="00:02:23.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="513" swimtime="00:02:07.36" resultid="6536" heatid="9558" lane="1" entrytime="00:02:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="150" swimtime="00:01:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5467" points="460" reactiontime="+92" swimtime="00:05:15.71" resultid="6537" heatid="9568" lane="0" entrytime="00:05:14.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:52.89" />
                    <SPLIT distance="200" swimtime="00:02:33.92" />
                    <SPLIT distance="250" swimtime="00:03:19.03" />
                    <SPLIT distance="300" swimtime="00:04:04.52" />
                    <SPLIT distance="350" swimtime="00:04:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5517" points="537" swimtime="00:01:01.27" resultid="6538" heatid="9578" lane="1" entrytime="00:01:01.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5636" points="501" reactiontime="+79" swimtime="00:04:37.07" resultid="6539" heatid="9613" lane="2" entrytime="00:04:36.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="150" swimtime="00:01:41.81" />
                    <SPLIT distance="200" swimtime="00:02:17.47" />
                    <SPLIT distance="250" swimtime="00:02:53.32" />
                    <SPLIT distance="300" swimtime="00:03:29.26" />
                    <SPLIT distance="350" swimtime="00:04:04.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MSC" nation="UKR" clubid="7778" name="MSC Euro-Lviv">
          <CONTACT city="Lviv" email="riff.lviv@gmail.com, eurolviv.masters@gmail.com" fax="+38 067 371 2151" internet="www.mastersswim.com.ua" name="Lyudmyla Khiresh" phone="+38 067 673 4796" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1969-11-03" firstname="Volodymyr" gender="M" lastname="Ivat" nation="UKR" athleteid="7782">
              <RESULTS>
                <RESULT eventid="1510" points="409" reactiontime="+89" swimtime="00:02:50.52" resultid="7783" heatid="9467" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="413" swimtime="00:01:16.71" resultid="7784" heatid="9511" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="7779">
              <RESULTS>
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="7780" heatid="9451" lane="3" entrytime="00:00:40.30" />
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="7781" heatid="9509" lane="8" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NABAIJI" nation="POL" clubid="7535" name="Nabaiji Team Decathlon">
          <CONTACT city="Warszawa" email="filip.wojciechowski@decathlon.com" name="Filip Wojciechowski" phone="731981998" street="Ostrobramska 97" zip="04-118" />
          <ATHLETES>
            <ATHLETE birthdate="1976-01-01" firstname="Agnieszka" gender="F" lastname="Dusza-Sabadasz" nation="POL" athleteid="7569">
              <RESULTS>
                <RESULT eventid="1133" points="210" reactiontime="+99" swimtime="00:00:39.76" resultid="7570" heatid="9310" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1458" points="179" reactiontime="+84" swimtime="00:00:47.96" resultid="7571" heatid="9443" lane="0" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Jacek" gender="M" lastname="Sokulski" nation="POL" athleteid="7587">
              <RESULTS>
                <RESULT eventid="1195" points="649" reactiontime="+73" swimtime="00:00:24.14" resultid="7588" heatid="9330" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="5331" points="722" reactiontime="+71" swimtime="00:00:25.00" resultid="7589" heatid="9527" lane="6" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Maciej" gender="M" lastname="Jekiełek" nation="POL" athleteid="7541">
              <RESULTS>
                <RESULT eventid="1195" points="434" reactiontime="+86" swimtime="00:00:27.60" resultid="7542" heatid="9330" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1476" points="376" reactiontime="+72" swimtime="00:00:33.30" resultid="7543" heatid="9455" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="7544" heatid="9510" lane="5" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Agnieszka" gender="F" lastname="Kos" nation="POL" athleteid="7552">
              <RESULTS>
                <RESULT eventid="1133" points="217" reactiontime="+94" swimtime="00:00:39.33" resultid="7553" heatid="9312" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1527" points="194" swimtime="00:01:29.29" resultid="7554" heatid="9471" lane="9" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="115" reactiontime="+97" swimtime="00:01:00.36" resultid="7555" heatid="9594" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="7536">
              <RESULTS>
                <RESULT eventid="1195" points="421" reactiontime="+75" swimtime="00:00:27.89" resultid="7537" heatid="9329" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="1476" points="370" reactiontime="+83" swimtime="00:00:33.48" resultid="7538" heatid="9455" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="5297" points="386" reactiontime="+70" swimtime="00:01:18.45" resultid="7539" heatid="9511" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="501" reactiontime="+78" swimtime="00:00:32.67" resultid="7540" heatid="9603" lane="3" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Izabella" gender="F" lastname="Grzegorczyk" nation="POL" athleteid="7578">
              <RESULTS>
                <RESULT eventid="1133" points="591" reactiontime="+75" swimtime="00:00:28.19" resultid="7579" heatid="9315" lane="5" entrytime="00:00:27.27" />
                <RESULT eventid="1212" points="627" reactiontime="+68" swimtime="00:02:27.35" resultid="7580" heatid="9340" lane="4" entrytime="00:02:23.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas równy Rekordowi Polski" eventid="1527" points="630" reactiontime="+71" swimtime="00:01:00.31" resultid="7581" heatid="9476" lane="5" entrytime="00:00:59.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="7545">
              <RESULTS>
                <RESULT eventid="1195" points="605" reactiontime="+78" swimtime="00:00:24.71" resultid="7546" heatid="9332" lane="6" entrytime="00:00:24.00" />
                <RESULT eventid="1544" points="609" reactiontime="+73" swimtime="00:00:55.32" resultid="7548" heatid="9490" lane="3" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="636" reactiontime="+73" swimtime="00:00:26.08" resultid="7549" heatid="9528" lane="3" entrytime="00:00:25.00" />
                <RESULT eventid="5399" points="454" reactiontime="+80" swimtime="00:02:12.67" resultid="7550" heatid="9558" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:02.39" />
                    <SPLIT distance="150" swimtime="00:01:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="589" reactiontime="+71" swimtime="00:00:59.41" resultid="7551" heatid="9578" lane="4" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="331" swimtime="00:10:53.19" resultid="9437" heatid="9362" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                    <SPLIT distance="150" swimtime="00:01:46.56" />
                    <SPLIT distance="200" swimtime="00:02:26.54" />
                    <SPLIT distance="250" swimtime="00:03:06.72" />
                    <SPLIT distance="300" swimtime="00:03:47.89" />
                    <SPLIT distance="350" swimtime="00:04:29.67" />
                    <SPLIT distance="400" swimtime="00:05:12.53" />
                    <SPLIT distance="450" swimtime="00:05:54.97" />
                    <SPLIT distance="500" swimtime="00:06:37.86" />
                    <SPLIT distance="550" swimtime="00:07:20.26" />
                    <SPLIT distance="600" swimtime="00:08:03.48" />
                    <SPLIT distance="650" swimtime="00:08:46.28" />
                    <SPLIT distance="700" swimtime="00:09:29.48" />
                    <SPLIT distance="750" swimtime="00:10:12.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="7572">
              <RESULTS>
                <RESULT eventid="1133" points="382" reactiontime="+81" swimtime="00:00:32.62" resultid="7573" heatid="9314" lane="1" entrytime="00:00:30.30" />
                <RESULT eventid="5279" points="320" swimtime="00:01:33.71" resultid="7574" heatid="9504" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="350" reactiontime="+80" swimtime="00:00:41.69" resultid="7575" heatid="9595" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Barbara" gender="F" lastname="Król" nation="POL" athleteid="7582">
              <RESULTS>
                <RESULT eventid="1133" points="159" swimtime="00:00:43.68" resultid="9307" heatid="9310" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Karolina" gender="F" lastname="Mazurek-Świstak" nation="POL" athleteid="7556">
              <RESULTS>
                <RESULT eventid="1133" points="519" reactiontime="+81" swimtime="00:00:29.45" resultid="7557" heatid="9315" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1493" points="455" reactiontime="+82" swimtime="00:03:00.83" resultid="7558" heatid="9461" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                    <SPLIT distance="150" swimtime="00:02:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="456" reactiontime="+79" swimtime="00:01:23.26" resultid="7559" heatid="9504" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="442" reactiontime="+85" swimtime="00:00:32.05" resultid="7560" heatid="9517" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="5568" points="488" reactiontime="+81" swimtime="00:00:37.34" resultid="7561" heatid="9596" lane="1" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Dominika" gender="F" lastname="Sasin" nation="POL" athleteid="7590">
              <RESULTS>
                <RESULT eventid="1458" points="493" reactiontime="+72" swimtime="00:00:34.25" resultid="7591" heatid="9446" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1527" points="577" reactiontime="+72" swimtime="00:01:02.09" resultid="7592" heatid="9476" lane="2" entrytime="00:01:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="568" reactiontime="+76" swimtime="00:00:29.49" resultid="7593" heatid="9517" lane="4" entrytime="00:00:29.13" />
                <RESULT eventid="5382" points="553" swimtime="00:02:17.62" resultid="7594" heatid="9547" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Aleksander" gender="M" lastname="Ziemiński" nation="POL" athleteid="7576">
              <RESULTS>
                <RESULT eventid="1195" points="188" reactiontime="+87" swimtime="00:00:36.49" resultid="7577" heatid="9320" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Mieszko" gender="M" lastname="Palmi-Kukiełko" nation="POL" athleteid="7562">
              <RESULTS>
                <RESULT eventid="1229" points="595" reactiontime="+74" swimtime="00:02:15.47" resultid="7563" heatid="9349" lane="4" entrytime="00:02:07.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="150" swimtime="00:01:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="498" reactiontime="+73" swimtime="00:18:18.33" resultid="7564" heatid="9365" lane="4" entrytime="00:17:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:39.37" />
                    <SPLIT distance="200" swimtime="00:02:15.49" />
                    <SPLIT distance="250" swimtime="00:02:51.93" />
                    <SPLIT distance="300" swimtime="00:03:28.69" />
                    <SPLIT distance="350" swimtime="00:04:05.87" />
                    <SPLIT distance="400" swimtime="00:04:43.57" />
                    <SPLIT distance="450" swimtime="00:05:21.35" />
                    <SPLIT distance="500" swimtime="00:05:58.94" />
                    <SPLIT distance="550" swimtime="00:06:36.00" />
                    <SPLIT distance="600" swimtime="00:07:13.14" />
                    <SPLIT distance="650" swimtime="00:07:50.53" />
                    <SPLIT distance="700" swimtime="00:08:27.67" />
                    <SPLIT distance="750" swimtime="00:09:04.99" />
                    <SPLIT distance="800" swimtime="00:09:42.59" />
                    <SPLIT distance="850" swimtime="00:10:20.13" />
                    <SPLIT distance="900" swimtime="00:10:57.59" />
                    <SPLIT distance="950" swimtime="00:11:35.01" />
                    <SPLIT distance="1000" swimtime="00:12:12.10" />
                    <SPLIT distance="1050" swimtime="00:12:49.34" />
                    <SPLIT distance="1100" swimtime="00:13:26.47" />
                    <SPLIT distance="1150" swimtime="00:14:03.94" />
                    <SPLIT distance="1200" swimtime="00:14:41.35" />
                    <SPLIT distance="1250" swimtime="00:15:18.38" />
                    <SPLIT distance="1300" swimtime="00:15:55.27" />
                    <SPLIT distance="1350" swimtime="00:16:31.91" />
                    <SPLIT distance="1400" swimtime="00:17:08.58" />
                    <SPLIT distance="1450" swimtime="00:17:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="574" reactiontime="+73" swimtime="00:00:28.92" resultid="7565" heatid="9457" lane="4" entrytime="00:00:27.21" />
                <RESULT eventid="1578" points="393" reactiontime="+74" swimtime="00:02:32.21" resultid="7566" heatid="9496" lane="4" entrytime="00:02:09.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="7567" heatid="9541" lane="4" entrytime="00:00:59.88" />
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="7568" heatid="9568" lane="4" entrytime="00:04:34.92" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="5433" status="DNS" swimtime="00:00:00.00" resultid="7599" heatid="9560" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7545" number="1" />
                    <RELAYPOSITION athleteid="7541" number="2" />
                    <RELAYPOSITION athleteid="7536" number="3" />
                    <RELAYPOSITION athleteid="7562" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1612" points="489" reactiontime="+67" swimtime="00:01:58.55" resultid="7600" heatid="9498" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="100" swimtime="00:01:01.39" />
                    <SPLIT distance="150" swimtime="00:01:31.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7541" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="7536" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="7587" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="7562" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="5416" points="416" reactiontime="+87" swimtime="00:02:09.37" resultid="7601" heatid="9559" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:40.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7590" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="7556" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="7552" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="7572" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="7602" heatid="9497" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7590" number="1" />
                    <RELAYPOSITION athleteid="7556" number="2" />
                    <RELAYPOSITION athleteid="7582" number="3" />
                    <RELAYPOSITION athleteid="7578" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" status="DNS" swimtime="00:00:00.00" resultid="7595" heatid="9608" lane="7" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7556" number="1" />
                    <RELAYPOSITION athleteid="7536" number="2" />
                    <RELAYPOSITION athleteid="7545" number="3" />
                    <RELAYPOSITION athleteid="7572" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1246" swimtime="00:01:51.63" resultid="7596" heatid="9353" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                    <SPLIT distance="150" swimtime="00:01:24.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7556" number="1" />
                    <RELAYPOSITION athleteid="7541" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="7578" number="3" />
                    <RELAYPOSITION athleteid="7536" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="5602" status="DNS" swimtime="00:00:00.00" resultid="7597" heatid="9608" lane="5" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7562" number="1" />
                    <RELAYPOSITION athleteid="7572" number="2" />
                    <RELAYPOSITION athleteid="7545" number="3" />
                    <RELAYPOSITION athleteid="7578" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1246" status="DNS" swimtime="00:00:00.00" resultid="7598" heatid="9353" lane="9">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7545" number="1" />
                    <RELAYPOSITION athleteid="7562" number="2" />
                    <RELAYPOSITION athleteid="7590" number="3" />
                    <RELAYPOSITION athleteid="7578" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+72" swimtime="00:01:59.54" resultid="7603" heatid="9353" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.78" />
                    <SPLIT distance="100" swimtime="00:00:56.52" />
                    <SPLIT distance="150" swimtime="00:01:32.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7572" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7552" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="7587" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="7576" number="4" reactiontime="-14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NMP" nation="CZE" clubid="6163" name="Neptun Masters Praha">
          <ATHLETES>
            <ATHLETE birthdate="1968-05-18" firstname="Hana" gender="F" lastname="Bohuslávková" nation="CZE" athleteid="6162">
              <RESULTS>
                <RESULT eventid="1212" points="424" reactiontime="+80" swimtime="00:02:47.78" resultid="6164" heatid="9339" lane="3" entrytime="00:02:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:02:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="451" reactiontime="+71" swimtime="00:03:01.27" resultid="6165" heatid="9461" lane="2" entrytime="00:03:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:27.77" />
                    <SPLIT distance="150" swimtime="00:02:14.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="470" reactiontime="+82" swimtime="00:01:22.48" resultid="6166" heatid="9504" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="458" reactiontime="+81" swimtime="00:00:38.14" resultid="6167" heatid="9596" lane="8" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-31" firstname="Šárka" gender="F" lastname="Landsmannová " nation="CZE" athleteid="6168">
              <RESULTS>
                <RESULT eventid="1263" points="559" reactiontime="+85" swimtime="00:09:48.42" resultid="6169" heatid="9355" lane="4" entrytime="00:09:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                    <SPLIT distance="200" swimtime="00:02:19.92" />
                    <SPLIT distance="250" swimtime="00:02:57.28" />
                    <SPLIT distance="300" swimtime="00:03:34.12" />
                    <SPLIT distance="350" swimtime="00:04:11.40" />
                    <SPLIT distance="400" swimtime="00:04:48.67" />
                    <SPLIT distance="450" swimtime="00:05:26.33" />
                    <SPLIT distance="500" swimtime="00:06:04.03" />
                    <SPLIT distance="550" swimtime="00:06:41.76" />
                    <SPLIT distance="600" swimtime="00:07:19.64" />
                    <SPLIT distance="650" swimtime="00:07:57.87" />
                    <SPLIT distance="700" swimtime="00:08:35.57" />
                    <SPLIT distance="750" swimtime="00:09:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="549" reactiontime="+82" swimtime="00:01:03.13" resultid="6170" heatid="9476" lane="0" entrytime="00:01:03.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="581" reactiontime="+83" swimtime="00:02:15.37" resultid="6171" heatid="9547" lane="2" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="576" reactiontime="+82" swimtime="00:04:44.15" resultid="6172" heatid="9609" lane="4" entrytime="00:04:52.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:43.75" />
                    <SPLIT distance="200" swimtime="00:02:20.15" />
                    <SPLIT distance="250" swimtime="00:02:56.54" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                    <SPLIT distance="350" swimtime="00:04:10.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="UKR" clubid="6042" name="nierzeszony UKR">
          <ATHLETES>
            <ATHLETE birthdate="1963-11-11" firstname="Mykhaylo" gender="M" lastname="Zakharchevskiy" nation="UKR" athleteid="6041">
              <RESULTS>
                <RESULT eventid="5365" points="174" reactiontime="+90" swimtime="00:01:32.82" resultid="6043" heatid="9537" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="164" reactiontime="+111" swimtime="00:07:25.42" resultid="6044" heatid="9565" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                    <SPLIT distance="100" swimtime="00:01:47.88" />
                    <SPLIT distance="150" swimtime="00:02:41.54" />
                    <SPLIT distance="200" swimtime="00:03:35.70" />
                    <SPLIT distance="250" swimtime="00:04:38.61" />
                    <SPLIT distance="300" swimtime="00:05:41.08" />
                    <SPLIT distance="350" swimtime="00:06:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6045" heatid="9586" lane="8" entrytime="00:03:15.00" />
                <RESULT eventid="5585" status="DNS" swimtime="00:00:00.00" resultid="6046" heatid="9598" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5773" name="nierzeszony ZD">
          <ATHLETES>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="Ziółkowski" nation="POL" athleteid="5772">
              <RESULTS>
                <RESULT eventid="1195" points="360" reactiontime="+83" swimtime="00:00:29.38" resultid="5774" heatid="9327" lane="1" entrytime="00:00:28.19" />
                <RESULT eventid="5331" points="318" reactiontime="+84" swimtime="00:00:32.86" resultid="5775" heatid="9524" lane="5" entrytime="00:00:30.83" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6387" name="niezrzeszeni">
          <ATHLETES>
            <ATHLETE birthdate="1994-09-14" firstname="Łukasz" gender="M" lastname="Machowski" nation="POL" athleteid="6394">
              <RESULTS>
                <RESULT eventid="1510" points="230" swimtime="00:03:26.57" resultid="6395" heatid="9465" lane="1" entrytime="00:03:16.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:37.74" />
                    <SPLIT distance="150" swimtime="00:02:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="163" swimtime="00:03:24.02" resultid="6396" heatid="9495" lane="9" entrytime="00:03:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="205" reactiontime="+78" swimtime="00:06:53.26" resultid="6397" heatid="9565" lane="4" entrytime="00:06:50.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:32.67" />
                    <SPLIT distance="150" swimtime="00:02:29.86" />
                    <SPLIT distance="200" swimtime="00:03:27.89" />
                    <SPLIT distance="250" swimtime="00:04:20.98" />
                    <SPLIT distance="300" swimtime="00:05:16.80" />
                    <SPLIT distance="350" swimtime="00:06:07.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="163" reactiontime="+80" swimtime="00:03:24.87" resultid="6398" heatid="9587" lane="5" entrytime="00:02:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:40.35" />
                    <SPLIT distance="150" swimtime="00:02:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="227" reactiontime="+86" swimtime="00:01:21.66" resultid="6399" heatid="9574" lane="3" entrytime="00:01:23.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-20" firstname="Aleksandra" gender="F" lastname="Marczewska" nation="POL" athleteid="6386">
              <RESULTS>
                <RESULT eventid="1458" points="305" reactiontime="+85" swimtime="00:00:40.20" resultid="6388" heatid="9445" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="1527" points="321" reactiontime="+87" swimtime="00:01:15.52" resultid="6389" heatid="9474" lane="0" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="266" reactiontime="+87" swimtime="00:00:37.98" resultid="6390" heatid="9516" lane="7" entrytime="00:00:34.80" />
                <RESULT eventid="5348" points="288" reactiontime="+75" swimtime="00:01:27.95" resultid="6391" heatid="9533" lane="0" entrytime="00:01:19.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="217" reactiontime="+89" swimtime="00:01:32.20" resultid="6392" heatid="9571" lane="8" entrytime="00:01:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="288" reactiontime="+84" swimtime="00:03:07.71" resultid="6393" heatid="9582" lane="0" entrytime="00:02:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                    <SPLIT distance="150" swimtime="00:02:19.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7720" name="niezrzeszona">
          <CONTACT city="Głosków" name="Zawadzka Jolanta" state="MAZ" street="Parkowa 2" zip="05-503" />
          <ATHLETES>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="7721">
              <RESULTS>
                <RESULT eventid="1212" points="223" swimtime="00:03:27.85" resultid="7722" heatid="9338" lane="1" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:38.83" />
                    <SPLIT distance="150" swimtime="00:02:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="244" swimtime="00:01:42.56" resultid="7723" heatid="9502" lane="1" entrytime="00:01:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="222" reactiontime="+82" swimtime="00:00:40.31" resultid="7724" heatid="9515" lane="0" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="7725" heatid="9593" lane="4" entrytime="00:00:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7680" name="Niezrzeszona JH">
          <ATHLETES>
            <ATHLETE birthdate="1996-03-07" firstname="Joanna" gender="F" lastname="Halagiera" nation="POL" athleteid="7679">
              <RESULTS>
                <RESULT eventid="1263" points="291" swimtime="00:12:10.88" resultid="7681" heatid="9355" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                    <SPLIT distance="200" swimtime="00:02:49.73" />
                    <SPLIT distance="250" swimtime="00:03:35.23" />
                    <SPLIT distance="300" swimtime="00:04:20.92" />
                    <SPLIT distance="350" swimtime="00:05:07.06" />
                    <SPLIT distance="400" swimtime="00:05:52.73" />
                    <SPLIT distance="450" swimtime="00:06:39.54" />
                    <SPLIT distance="500" swimtime="00:07:26.64" />
                    <SPLIT distance="550" swimtime="00:08:14.22" />
                    <SPLIT distance="600" swimtime="00:09:01.24" />
                    <SPLIT distance="650" swimtime="00:09:49.50" />
                    <SPLIT distance="700" swimtime="00:10:36.76" />
                    <SPLIT distance="750" swimtime="00:11:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="238" swimtime="00:03:16.38" resultid="7682" heatid="9492" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="296" reactiontime="+79" swimtime="00:06:39.30" resultid="7683" heatid="9563" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="200" swimtime="00:03:10.80" />
                    <SPLIT distance="250" swimtime="00:04:08.25" />
                    <SPLIT distance="300" swimtime="00:05:05.02" />
                    <SPLIT distance="350" swimtime="00:05:52.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="311" swimtime="00:05:48.94" resultid="7684" heatid="9609" lane="1" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:21.39" />
                    <SPLIT distance="150" swimtime="00:02:05.93" />
                    <SPLIT distance="200" swimtime="00:02:50.85" />
                    <SPLIT distance="250" swimtime="00:03:36.25" />
                    <SPLIT distance="300" swimtime="00:04:21.67" />
                    <SPLIT distance="350" swimtime="00:05:06.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6376" name="niezrzeszona KM">
          <ATHLETES>
            <ATHLETE birthdate="1975-01-12" firstname="Maja" gender="F" lastname="Klusek" nation="POL" athleteid="6375">
              <RESULTS>
                <RESULT eventid="5450" points="287" reactiontime="+97" swimtime="00:06:43.56" resultid="6378" heatid="9563" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:02:24.62" />
                    <SPLIT distance="200" swimtime="00:03:19.02" />
                    <SPLIT distance="250" swimtime="00:04:13.88" />
                    <SPLIT distance="300" swimtime="00:05:10.19" />
                    <SPLIT distance="350" swimtime="00:05:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="232" swimtime="00:01:30.20" resultid="6379" heatid="9571" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7139" name="niezrzeszona KZ">
          <ATHLETES>
            <ATHLETE birthdate="1995-09-29" firstname="Zuzanna" gender="F" lastname="Kasperczak" nation="POL" athleteid="7138">
              <RESULTS>
                <RESULT eventid="1527" points="118" swimtime="00:01:45.23" resultid="7140" heatid="9469" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7793" name="niezrzeszona LB" />
        <CLUB type="CLUB" code="N" nation="POL" clubid="5982" name="niezrzeszona PA">
          <ATHLETES>
            <ATHLETE birthdate="1947-07-15" firstname="Alina" gender="F" lastname="Piekarska" nation="POL" athleteid="5981">
              <RESULTS>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="5568" status="DSQ" swimtime="00:02:51.48" resultid="5983" heatid="9591" lane="5" entrytime="00:02:13.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6105" name="niezrzeszona RA">
          <ATHLETES>
            <ATHLETE birthdate="1997-05-30" firstname="Adrianna" gender="F" lastname="Rzewuska" nation="POL" athleteid="6104">
              <RESULTS>
                <RESULT eventid="1458" points="460" reactiontime="+70" swimtime="00:00:35.05" resultid="6106" heatid="9446" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="5348" points="413" reactiontime="+68" swimtime="00:01:18.01" resultid="6107" heatid="9533" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6381" name="niezrzeszona SK">
          <ATHLETES>
            <ATHLETE birthdate="1976-03-14" firstname="Katarzyna" gender="F" lastname="Szwagiel" nation="POL" athleteid="6380">
              <RESULTS>
                <RESULT eventid="1212" points="307" swimtime="00:03:06.86" resultid="6382" heatid="9339" lane="1" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:02:23.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="258" reactiontime="+108" swimtime="00:12:40.96" resultid="6383" heatid="9356" lane="0" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:12.83" />
                    <SPLIT distance="200" swimtime="00:03:00.12" />
                    <SPLIT distance="250" swimtime="00:03:48.10" />
                    <SPLIT distance="300" swimtime="00:04:36.70" />
                    <SPLIT distance="350" swimtime="00:05:25.12" />
                    <SPLIT distance="400" swimtime="00:06:14.15" />
                    <SPLIT distance="450" swimtime="00:07:02.79" />
                    <SPLIT distance="500" swimtime="00:07:51.39" />
                    <SPLIT distance="550" swimtime="00:08:39.88" />
                    <SPLIT distance="600" swimtime="00:09:28.76" />
                    <SPLIT distance="650" swimtime="00:10:17.32" />
                    <SPLIT distance="700" swimtime="00:11:05.75" />
                    <SPLIT distance="750" swimtime="00:11:54.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="311" reactiontime="+94" swimtime="00:02:46.61" resultid="6384" heatid="9545" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="284" reactiontime="+106" swimtime="00:05:59.67" resultid="6385" heatid="9610" lane="0" entrytime="00:06:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                    <SPLIT distance="200" swimtime="00:02:54.81" />
                    <SPLIT distance="250" swimtime="00:03:41.26" />
                    <SPLIT distance="300" swimtime="00:04:28.45" />
                    <SPLIT distance="350" swimtime="00:05:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5667" name="niezrzeszona WZ">
          <ATHLETES>
            <ATHLETE birthdate="1952-04-04" firstname="Zdzisława" gender="F" lastname="Wiese" nation="POL" athleteid="5666">
              <RESULTS>
                <RESULT eventid="1493" points="79" swimtime="00:05:23.67" resultid="5669" heatid="9458" lane="6" entrytime="00:05:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.43" />
                    <SPLIT distance="100" swimtime="00:02:32.05" />
                    <SPLIT distance="150" swimtime="00:03:59.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="84" reactiontime="+118" swimtime="00:02:26.03" resultid="5670" heatid="9500" lane="4" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="5671" heatid="9592" lane="8" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9301" name="Niezrzeszony">
          <CONTACT city="Dolaszewo" email="andrzej.harenda@op.pl" name="Harenda Andrzej" phone="608629706" state="WIELK" street="Dębowa 1" zip="64-930" />
          <ATHLETES>
            <ATHLETE birthdate="1968-12-28" firstname="Andrzej" gender="M" lastname="Harenda" nation="POL" athleteid="9302">
              <RESULTS>
                <RESULT eventid="1510" points="225" swimtime="00:03:28.03" resultid="9303" heatid="9465" lane="6" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:02:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="272" reactiontime="+89" swimtime="00:01:12.37" resultid="9304" heatid="9482" lane="5" entrytime="00:01:09.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="9305" heatid="9508" lane="7" entrytime="00:01:33.56" entrycourse="SCM" />
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="9306" heatid="9552" lane="4" entrytime="00:02:45.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6127" name="Niezrzeszony">
          <CONTACT city="BYDGOSZCZ" email="MACIEJLUBAS@GMAIL.COM" name="LUBAS" phone="667905450" state="KUJAW" street="BOCIANOWO" zip="85-042" />
          <ATHLETES>
            <ATHLETE birthdate="1978-01-05" firstname="Maciej" gender="M" lastname="Lubas" nation="POL" athleteid="6128">
              <RESULTS>
                <RESULT eventid="1510" points="329" reactiontime="+89" swimtime="00:03:03.34" resultid="6129" heatid="9467" lane="5" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="344" reactiontime="+81" swimtime="00:01:21.53" resultid="6130" heatid="9511" lane="7" entrytime="00:01:17.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="391" reactiontime="+84" swimtime="00:00:35.48" resultid="6131" heatid="9603" lane="7" entrytime="00:00:34.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" region="POM" clubid="5680" name="Niezrzeszony">
          <CONTACT city="Gdynia" email="januszmasters1@gmail.com" name="Płonka" phone="58 6291045" street="Iwaszkiewicza 2C m.2" zip="81-597" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="5681">
              <RESULTS>
                <RESULT eventid="1229" points="51" swimtime="00:05:06.22" resultid="5682" heatid="9343" lane="9" entrytime="00:04:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.20" />
                    <SPLIT distance="100" swimtime="00:02:28.72" />
                    <SPLIT distance="150" swimtime="00:03:59.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="82" reactiontime="+81" swimtime="00:00:55.15" resultid="5683" heatid="9449" lane="0" entrytime="00:00:57.00" />
                <RESULT eventid="1578" points="34" reactiontime="+108" swimtime="00:05:42.73" resultid="5684" heatid="9493" lane="8" entrytime="00:05:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.52" />
                    <SPLIT distance="100" swimtime="00:02:39.83" />
                    <SPLIT distance="150" swimtime="00:04:12.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="59" reactiontime="+115" swimtime="00:00:57.45" resultid="5685" heatid="9519" lane="9" entrytime="00:00:56.00" />
                <RESULT eventid="5399" points="47" reactiontime="+105" swimtime="00:04:41.92" resultid="5686" heatid="9549" lane="0" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.40" />
                    <SPLIT distance="100" swimtime="00:02:15.99" />
                    <SPLIT distance="150" swimtime="00:03:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="37" reactiontime="+106" swimtime="00:02:29.28" resultid="5687" heatid="9572" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="46" swimtime="00:10:11.49" resultid="9622" heatid="9621" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5991" name="niezrzeszony">
          <CONTACT name="Gogacz" />
          <ATHLETES>
            <ATHLETE birthdate="1960-12-21" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="5997">
              <RESULTS>
                <RESULT eventid="1314" points="179" swimtime="00:25:43.93" resultid="5998" heatid="9367" lane="6" entrytime="00:26:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                    <SPLIT distance="150" swimtime="00:02:18.71" />
                    <SPLIT distance="200" swimtime="00:03:09.44" />
                    <SPLIT distance="250" swimtime="00:04:01.14" />
                    <SPLIT distance="300" swimtime="00:04:52.67" />
                    <SPLIT distance="350" swimtime="00:07:29.79" />
                    <SPLIT distance="400" swimtime="00:06:37.10" />
                    <SPLIT distance="450" swimtime="00:09:14.55" />
                    <SPLIT distance="500" swimtime="00:08:21.34" />
                    <SPLIT distance="550" swimtime="00:12:42.88" />
                    <SPLIT distance="600" swimtime="00:10:04.88" />
                    <SPLIT distance="650" swimtime="00:14:27.44" />
                    <SPLIT distance="700" swimtime="00:11:49.06" />
                    <SPLIT distance="750" swimtime="00:16:11.00" />
                    <SPLIT distance="800" swimtime="00:13:33.62" />
                    <SPLIT distance="850" swimtime="00:17:54.51" />
                    <SPLIT distance="900" swimtime="00:15:17.39" />
                    <SPLIT distance="950" swimtime="00:21:24.30" />
                    <SPLIT distance="1000" swimtime="00:17:01.35" />
                    <SPLIT distance="1050" swimtime="00:23:09.58" />
                    <SPLIT distance="1100" swimtime="00:18:45.80" />
                    <SPLIT distance="1150" swimtime="00:24:54.51" />
                    <SPLIT distance="1200" swimtime="00:20:30.60" />
                    <SPLIT distance="1300" swimtime="00:22:15.54" />
                    <SPLIT distance="1400" swimtime="00:24:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="174" reactiontime="+115" swimtime="00:01:23.91" resultid="5999" heatid="9480" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="120" reactiontime="+118" swimtime="00:08:13.24" resultid="6000" heatid="9565" lane="0" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                    <SPLIT distance="100" swimtime="00:02:00.06" />
                    <SPLIT distance="150" swimtime="00:03:10.86" />
                    <SPLIT distance="200" swimtime="00:04:20.38" />
                    <SPLIT distance="250" swimtime="00:05:30.73" />
                    <SPLIT distance="300" swimtime="00:06:40.80" />
                    <SPLIT distance="350" swimtime="00:07:26.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="196" swimtime="00:06:18.63" resultid="6001" heatid="9618" lane="6" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                    <SPLIT distance="200" swimtime="00:03:02.79" />
                    <SPLIT distance="250" swimtime="00:03:53.83" />
                    <SPLIT distance="300" swimtime="00:04:41.93" />
                    <SPLIT distance="350" swimtime="00:05:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" athleteid="5992">
              <RESULTS>
                <RESULT eventid="1314" points="385" reactiontime="+92" swimtime="00:19:56.53" resultid="5993" heatid="9365" lane="0" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                    <SPLIT distance="200" swimtime="00:02:34.75" />
                    <SPLIT distance="250" swimtime="00:03:14.86" />
                    <SPLIT distance="300" swimtime="00:03:54.78" />
                    <SPLIT distance="350" swimtime="00:04:34.36" />
                    <SPLIT distance="400" swimtime="00:05:14.31" />
                    <SPLIT distance="450" swimtime="00:05:53.57" />
                    <SPLIT distance="500" swimtime="00:06:33.29" />
                    <SPLIT distance="550" swimtime="00:07:12.94" />
                    <SPLIT distance="600" swimtime="00:07:52.72" />
                    <SPLIT distance="650" swimtime="00:08:32.27" />
                    <SPLIT distance="700" swimtime="00:09:12.58" />
                    <SPLIT distance="750" swimtime="00:09:52.22" />
                    <SPLIT distance="800" swimtime="00:10:32.02" />
                    <SPLIT distance="850" swimtime="00:11:11.75" />
                    <SPLIT distance="900" swimtime="00:11:52.45" />
                    <SPLIT distance="950" swimtime="00:12:32.36" />
                    <SPLIT distance="1000" swimtime="00:13:12.73" />
                    <SPLIT distance="1050" swimtime="00:13:52.69" />
                    <SPLIT distance="1100" swimtime="00:14:33.10" />
                    <SPLIT distance="1150" swimtime="00:15:13.48" />
                    <SPLIT distance="1200" swimtime="00:15:54.46" />
                    <SPLIT distance="1250" swimtime="00:16:34.85" />
                    <SPLIT distance="1300" swimtime="00:17:15.21" />
                    <SPLIT distance="1350" swimtime="00:17:55.84" />
                    <SPLIT distance="1400" swimtime="00:18:37.08" />
                    <SPLIT distance="1450" swimtime="00:19:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="348" swimtime="00:02:38.46" resultid="5994" heatid="9496" lane="9" entrytime="00:02:37.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="333" swimtime="00:05:51.73" resultid="5995" heatid="9566" lane="6" entrytime="00:06:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:02:07.44" />
                    <SPLIT distance="200" swimtime="00:02:54.80" />
                    <SPLIT distance="250" swimtime="00:03:44.18" />
                    <SPLIT distance="300" swimtime="00:04:33.93" />
                    <SPLIT distance="350" swimtime="00:05:14.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="371" swimtime="00:05:06.00" resultid="5996" heatid="9618" lane="1" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:13.32" />
                    <SPLIT distance="150" swimtime="00:01:52.65" />
                    <SPLIT distance="200" swimtime="00:02:32.01" />
                    <SPLIT distance="250" swimtime="00:03:11.04" />
                    <SPLIT distance="300" swimtime="00:03:50.08" />
                    <SPLIT distance="350" swimtime="00:04:28.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5700" name="Niezrzeszony">
          <CONTACT city="WARSZAWA" email="zbyszek@paluszak.pl" name="PALUSZAK ZBIGNIEW" phone="601643732" state="MAZ" street="HUCULSKA 3/35" zip="00-730" />
          <ATHLETES>
            <ATHLETE birthdate="1967-02-17" firstname="Zbigniew" gender="M" lastname="Paluszak" nation="POL" athleteid="5701">
              <RESULTS>
                <RESULT eventid="1510" points="134" reactiontime="+79" swimtime="00:04:07.25" resultid="5702" heatid="9463" lane="8" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                    <SPLIT distance="100" swimtime="00:01:55.18" />
                    <SPLIT distance="150" swimtime="00:03:02.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="135" swimtime="00:01:51.18" resultid="5703" heatid="9506" lane="6" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="97" swimtime="00:03:41.28" resultid="5704" heatid="9549" lane="6" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                    <SPLIT distance="100" swimtime="00:01:42.29" />
                    <SPLIT distance="150" swimtime="00:02:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="147" reactiontime="+84" swimtime="00:00:49.13" resultid="5705" heatid="9598" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="5636" points="99" swimtime="00:07:54.69" resultid="5706" heatid="9619" lane="1" entrytime="00:08:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:43.31" />
                    <SPLIT distance="150" swimtime="00:02:44.47" />
                    <SPLIT distance="200" swimtime="00:03:46.53" />
                    <SPLIT distance="250" swimtime="00:04:50.26" />
                    <SPLIT distance="300" swimtime="00:05:53.24" />
                    <SPLIT distance="350" swimtime="00:06:55.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6082" name="Niezrzeszony Białystok">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko" phone="797309140" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="6083">
              <RESULTS>
                <RESULT eventid="1195" points="388" reactiontime="+80" swimtime="00:00:28.65" resultid="6084" heatid="9326" lane="3" entrytime="00:00:28.95" />
                <RESULT eventid="1229" points="337" reactiontime="+79" swimtime="00:02:43.80" resultid="6085" heatid="9346" lane="7" entrytime="00:02:45.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:02:05.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="305" reactiontime="+63" swimtime="00:00:35.68" resultid="6086" heatid="9453" lane="2" entrytime="00:00:35.95" />
                <RESULT eventid="1544" points="402" reactiontime="+80" swimtime="00:01:03.52" resultid="6087" heatid="9484" lane="4" entrytime="00:01:04.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="390" reactiontime="+83" swimtime="00:00:30.69" resultid="6088" heatid="9524" lane="3" entrytime="00:00:30.85" />
                <RESULT eventid="5365" points="286" reactiontime="+77" swimtime="00:01:18.69" resultid="6089" heatid="9538" lane="8" entrytime="00:01:18.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="358" reactiontime="+83" swimtime="00:01:10.14" resultid="6090" heatid="9575" lane="4" entrytime="00:01:12.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="335" reactiontime="+87" swimtime="00:00:37.33" resultid="6091" heatid="9601" lane="5" entrytime="00:00:37.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7122" name="niezrzeszony Białystok">
          <ATHLETES>
            <ATHLETE birthdate="1943-01-01" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="7121">
              <RESULTS>
                <RESULT eventid="1195" points="125" reactiontime="+107" swimtime="00:00:41.77" resultid="7123" heatid="9319" lane="6" entrytime="00:00:40.50" />
                <RESULT eventid="1280" points="105" reactiontime="+117" swimtime="00:15:55.85" resultid="7124" heatid="9362" lane="0" entrytime="00:15:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.94" />
                    <SPLIT distance="100" swimtime="00:01:52.25" />
                    <SPLIT distance="150" swimtime="00:02:52.66" />
                    <SPLIT distance="200" swimtime="00:03:52.61" />
                    <SPLIT distance="250" swimtime="00:04:52.43" />
                    <SPLIT distance="300" swimtime="00:05:52.19" />
                    <SPLIT distance="350" swimtime="00:06:52.88" />
                    <SPLIT distance="400" swimtime="00:07:54.03" />
                    <SPLIT distance="450" swimtime="00:08:54.76" />
                    <SPLIT distance="500" swimtime="00:09:55.82" />
                    <SPLIT distance="550" swimtime="00:10:57.42" />
                    <SPLIT distance="600" swimtime="00:11:58.83" />
                    <SPLIT distance="650" swimtime="00:12:59.52" />
                    <SPLIT distance="700" swimtime="00:13:59.41" />
                    <SPLIT distance="750" swimtime="00:14:59.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="84" reactiontime="+109" swimtime="00:00:54.69" resultid="7125" heatid="9449" lane="6" entrytime="00:00:51.00" />
                <RESULT eventid="1544" points="115" reactiontime="+103" swimtime="00:01:36.20" resultid="7126" heatid="9479" lane="8" entrytime="00:01:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="116" reactiontime="+130" swimtime="00:00:45.90" resultid="7127" heatid="9519" lane="3" entrytime="00:00:45.50" />
                <RESULT eventid="5399" points="108" reactiontime="+106" swimtime="00:03:34.12" resultid="7128" heatid="9550" lane="7" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:44.38" />
                    <SPLIT distance="150" swimtime="00:02:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="63" reactiontime="+114" swimtime="00:02:04.91" resultid="7129" heatid="9572" lane="4" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="60" reactiontime="+117" swimtime="00:04:44.48" resultid="7130" heatid="9584" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.40" />
                    <SPLIT distance="100" swimtime="00:02:23.23" />
                    <SPLIT distance="150" swimtime="00:03:39.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7716" name="niezrzeszony CB">
          <ATHLETES>
            <ATHLETE birthdate="1948-06-28" firstname="Bolesław" gender="M" lastname="Czyż" nation="POL" athleteid="7715">
              <RESULTS>
                <RESULT eventid="1578" points="58" reactiontime="+107" swimtime="00:04:46.76" resultid="7717" heatid="9493" lane="2" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.02" />
                    <SPLIT distance="100" swimtime="00:02:18.42" />
                    <SPLIT distance="150" swimtime="00:03:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="86" swimtime="00:09:11.79" resultid="7718" heatid="9565" lane="9" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.15" />
                    <SPLIT distance="100" swimtime="00:02:13.75" />
                    <SPLIT distance="150" swimtime="00:03:24.94" />
                    <SPLIT distance="200" swimtime="00:04:31.52" />
                    <SPLIT distance="250" swimtime="00:05:45.94" />
                    <SPLIT distance="300" swimtime="00:07:02.48" />
                    <SPLIT distance="350" swimtime="00:08:09.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="7719" heatid="9584" lane="3" entrytime="00:04:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5661" name="niezrzeszony DR">
          <ATHLETES>
            <ATHLETE birthdate="1976-10-28" firstname="Robert" gender="M" lastname="Drzazga" nation="POL" athleteid="5660">
              <RESULTS>
                <RESULT eventid="1544" points="293" swimtime="00:01:10.58" resultid="5662" heatid="9483" lane="1" entrytime="00:01:08.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="279" reactiontime="+87" swimtime="00:00:34.30" resultid="5663" heatid="9522" lane="9" entrytime="00:00:33.86" />
                <RESULT eventid="5399" points="246" reactiontime="+83" swimtime="00:02:42.76" resultid="5664" heatid="9553" lane="3" entrytime="00:02:34.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:01.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7208" name="niezrzeszony GA">
          <ATHLETES>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="7207">
              <RESULTS>
                <RESULT eventid="1133" points="362" reactiontime="+76" swimtime="00:00:33.21" resultid="7209" heatid="9312" lane="4" entrytime="00:00:33.12" />
                <RESULT eventid="1263" points="311" reactiontime="+77" swimtime="00:11:54.98" resultid="7210" heatid="9356" lane="4" entrytime="00:12:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:01:59.36" />
                    <SPLIT distance="200" swimtime="00:02:42.71" />
                    <SPLIT distance="250" swimtime="00:03:27.38" />
                    <SPLIT distance="300" swimtime="00:04:12.71" />
                    <SPLIT distance="350" swimtime="00:04:58.77" />
                    <SPLIT distance="400" swimtime="00:05:45.15" />
                    <SPLIT distance="450" swimtime="00:06:31.66" />
                    <SPLIT distance="500" swimtime="00:07:18.37" />
                    <SPLIT distance="550" swimtime="00:08:05.33" />
                    <SPLIT distance="600" swimtime="00:08:52.39" />
                    <SPLIT distance="650" swimtime="00:09:38.50" />
                    <SPLIT distance="700" swimtime="00:10:24.78" />
                    <SPLIT distance="750" swimtime="00:11:10.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="287" reactiontime="+90" swimtime="00:00:41.01" resultid="7211" heatid="9443" lane="6" entrytime="00:00:41.32" />
                <RESULT eventid="1493" points="306" reactiontime="+81" swimtime="00:03:26.28" resultid="7212" heatid="9459" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:35.96" />
                    <SPLIT distance="150" swimtime="00:02:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="313" reactiontime="+45" swimtime="00:01:34.38" resultid="7213" heatid="9503" lane="7" entrytime="00:01:32.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="354" reactiontime="+64" swimtime="00:02:39.61" resultid="7214" heatid="9546" lane="7" entrytime="00:02:45.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="329" reactiontime="+78" swimtime="00:00:42.56" resultid="7215" heatid="9594" lane="4" entrytime="00:00:42.08" />
                <RESULT eventid="5619" points="328" swimtime="00:05:42.65" resultid="7216" heatid="9610" lane="6" entrytime="00:05:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:02:01.73" />
                    <SPLIT distance="200" swimtime="00:02:46.07" />
                    <SPLIT distance="250" swimtime="00:03:30.24" />
                    <SPLIT distance="300" swimtime="00:04:14.98" />
                    <SPLIT distance="350" swimtime="00:04:59.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7167" name="niezrzeszony JG">
          <ATHLETES>
            <ATHLETE birthdate="1959-02-19" firstname="Grzegorz" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="7166">
              <RESULTS>
                <RESULT eventid="1195" points="188" reactiontime="+119" swimtime="00:00:36.44" resultid="7168" heatid="9321" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1476" points="153" reactiontime="+98" swimtime="00:00:44.85" resultid="7169" heatid="9450" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6037" name="niezrzeszony KJ">
          <ATHLETES>
            <ATHLETE birthdate="1998-05-04" firstname="Jędrzej" gender="M" lastname="Kuczma" nation="POL" athleteid="6036">
              <RESULTS>
                <RESULT eventid="1195" points="484" reactiontime="+75" swimtime="00:00:26.63" resultid="6038" heatid="9325" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1544" points="523" swimtime="00:00:58.22" resultid="6039" heatid="9487" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="456" reactiontime="+76" swimtime="00:00:29.13" resultid="6040" heatid="9525" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6034" name="niezrzeszony KK">
          <ATHLETES>
            <ATHLETE birthdate="1974-12-30" firstname="Krzysztof" gender="M" lastname="Krzak" nation="POL" athleteid="6033">
              <RESULTS>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6047" heatid="9538" lane="6" entrytime="00:01:17.31" />
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="6048" heatid="9566" lane="4" entrytime="00:06:05.90" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="6049" heatid="9588" lane="4" entrytime="00:02:43.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5758" name="niezrzeszony Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1938-04-28" firstname="Andrzej" gender="M" lastname="Wiśniewski" nation="POL" athleteid="5757">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1314" points="71" reactiontime="+133" swimtime="00:34:54.91" resultid="5759" heatid="9368" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.65" />
                    <SPLIT distance="100" swimtime="00:02:05.88" />
                    <SPLIT distance="150" swimtime="00:03:14.20" />
                    <SPLIT distance="200" swimtime="00:04:23.73" />
                    <SPLIT distance="250" swimtime="00:05:33.09" />
                    <SPLIT distance="300" swimtime="00:06:42.29" />
                    <SPLIT distance="350" swimtime="00:07:51.02" />
                    <SPLIT distance="400" swimtime="00:09:00.63" />
                    <SPLIT distance="450" swimtime="00:10:10.13" />
                    <SPLIT distance="500" swimtime="00:11:19.83" />
                    <SPLIT distance="550" swimtime="00:12:29.59" />
                    <SPLIT distance="600" swimtime="00:13:39.69" />
                    <SPLIT distance="650" swimtime="00:14:49.35" />
                    <SPLIT distance="700" swimtime="00:15:59.68" />
                    <SPLIT distance="750" swimtime="00:17:09.33" />
                    <SPLIT distance="800" swimtime="00:18:20.12" />
                    <SPLIT distance="850" swimtime="00:19:30.82" />
                    <SPLIT distance="900" swimtime="00:20:41.15" />
                    <SPLIT distance="950" swimtime="00:21:51.47" />
                    <SPLIT distance="1000" swimtime="00:23:02.29" />
                    <SPLIT distance="1050" swimtime="00:24:12.95" />
                    <SPLIT distance="1100" swimtime="00:25:25.93" />
                    <SPLIT distance="1150" swimtime="00:26:37.85" />
                    <SPLIT distance="1200" swimtime="00:27:49.56" />
                    <SPLIT distance="1250" swimtime="00:29:00.32" />
                    <SPLIT distance="1300" swimtime="00:30:12.58" />
                    <SPLIT distance="1350" swimtime="00:31:24.06" />
                    <SPLIT distance="1400" swimtime="00:32:34.96" />
                    <SPLIT distance="1450" swimtime="00:33:46.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5761" name="niezrzeszony KT">
          <ATHLETES>
            <ATHLETE birthdate="1974-06-11" firstname="Tomasz" gender="M" lastname="Karczewski" nation="POL" athleteid="5760">
              <RESULTS>
                <RESULT eventid="1195" points="327" reactiontime="+86" swimtime="00:00:30.33" resultid="5762" heatid="9323" lane="2" entrytime="00:00:30.90" />
                <RESULT eventid="5331" points="344" reactiontime="+83" swimtime="00:00:32.00" resultid="5763" heatid="9522" lane="4" entrytime="00:00:32.46" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5811" name="niezrzeszony MA">
          <ATHLETES>
            <ATHLETE birthdate="1954-10-24" firstname="Andrzej" gender="M" lastname="Marszałek" nation="POL" athleteid="5810">
              <RESULTS>
                <RESULT eventid="1544" points="125" swimtime="00:01:33.77" resultid="5812" heatid="9478" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="96" reactiontime="+102" swimtime="00:00:48.82" resultid="5813" heatid="9519" lane="8" entrytime="00:00:53.00" />
                <RESULT eventid="5399" points="114" swimtime="00:03:29.90" resultid="5814" heatid="9550" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                    <SPLIT distance="150" swimtime="00:02:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="82" swimtime="00:01:54.53" resultid="5815" heatid="9573" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="118" swimtime="00:07:28.02" resultid="5816" heatid="9619" lane="6" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:45.17" />
                    <SPLIT distance="150" swimtime="00:02:43.59" />
                    <SPLIT distance="200" swimtime="00:03:39.08" />
                    <SPLIT distance="250" swimtime="00:04:36.41" />
                    <SPLIT distance="300" swimtime="00:05:34.25" />
                    <SPLIT distance="350" swimtime="00:06:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5765" name="niezrzeszony NL">
          <ATHLETES>
            <ATHLETE birthdate="1979-04-05" firstname="Bartłomiej" gender="M" lastname="Sieczyński" nation="POL" athleteid="5764">
              <RESULTS>
                <RESULT eventid="1195" points="317" reactiontime="+77" swimtime="00:00:30.64" resultid="5766" heatid="9324" lane="6" entrytime="00:00:29.70" />
                <RESULT eventid="1544" points="339" reactiontime="+73" swimtime="00:01:07.25" resultid="5767" heatid="9484" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="288" reactiontime="+78" swimtime="00:00:33.93" resultid="5768" heatid="9522" lane="7" entrytime="00:00:33.20" />
                <RESULT eventid="5399" points="338" swimtime="00:02:26.33" resultid="5769" heatid="9554" lane="9" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="192" swimtime="00:01:26.35" resultid="5770" heatid="9574" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="329" swimtime="00:05:18.76" resultid="5771" heatid="9615" lane="9" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                    <SPLIT distance="200" swimtime="00:02:31.77" />
                    <SPLIT distance="250" swimtime="00:03:13.21" />
                    <SPLIT distance="300" swimtime="00:03:55.36" />
                    <SPLIT distance="350" swimtime="00:04:38.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6109" name="niezrzeszony Radom">
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Włodzimierz" gender="M" lastname="Zieleziński" nation="POL" athleteid="6108">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="6110" heatid="9321" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1280" points="121" swimtime="00:15:11.71" resultid="6111" heatid="9362" lane="7" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:35.68" />
                    <SPLIT distance="150" swimtime="00:02:32.29" />
                    <SPLIT distance="200" swimtime="00:03:30.28" />
                    <SPLIT distance="250" swimtime="00:04:28.16" />
                    <SPLIT distance="300" swimtime="00:05:26.59" />
                    <SPLIT distance="350" swimtime="00:06:25.37" />
                    <SPLIT distance="400" swimtime="00:07:24.66" />
                    <SPLIT distance="450" swimtime="00:08:24.02" />
                    <SPLIT distance="500" swimtime="00:09:23.07" />
                    <SPLIT distance="550" swimtime="00:10:22.22" />
                    <SPLIT distance="600" swimtime="00:11:21.95" />
                    <SPLIT distance="650" swimtime="00:12:21.96" />
                    <SPLIT distance="700" swimtime="00:13:20.56" />
                    <SPLIT distance="750" swimtime="00:14:17.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="177" reactiontime="+79" swimtime="00:00:42.77" resultid="6112" heatid="9451" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6113" heatid="9481" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="5365" points="147" reactiontime="+82" swimtime="00:01:38.23" resultid="6114" heatid="9536" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="6115" heatid="9551" lane="1" entrytime="00:03:05.00" />
                <RESULT eventid="5551" points="108" reactiontime="+76" swimtime="00:03:54.44" resultid="6116" heatid="9585" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.97" />
                    <SPLIT distance="100" swimtime="00:01:49.94" />
                    <SPLIT distance="150" swimtime="00:02:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="119" swimtime="00:07:27.18" resultid="6117" heatid="9617" lane="9" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:38.94" />
                    <SPLIT distance="150" swimtime="00:02:35.82" />
                    <SPLIT distance="200" swimtime="00:03:34.66" />
                    <SPLIT distance="250" swimtime="00:04:33.27" />
                    <SPLIT distance="300" swimtime="00:05:33.26" />
                    <SPLIT distance="350" swimtime="00:06:31.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7461" name="niezrzeszony SE">
          <ATHLETES>
            <ATHLETE birthdate="1988-05-18" firstname="Emil" gender="M" lastname="Strumiński" nation="POL" athleteid="7460">
              <RESULTS>
                <RESULT eventid="1195" points="467" reactiontime="+72" swimtime="00:00:26.94" resultid="7462" heatid="9328" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1544" points="496" reactiontime="+69" swimtime="00:00:59.24" resultid="7463" heatid="9488" lane="2" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="456" reactiontime="+74" swimtime="00:00:29.13" resultid="7464" heatid="9526" lane="7" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="6344" name="niezrzeszony SL">
          <ATHLETES>
            <ATHLETE birthdate="1965-06-11" firstname="Ludwik" gender="M" lastname="Schwarz" nation="BLR" athleteid="6343">
              <RESULTS>
                <RESULT eventid="1195" points="199" reactiontime="+107" swimtime="00:00:35.81" resultid="6345" heatid="9320" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1280" points="169" reactiontime="+94" swimtime="00:13:36.33" resultid="6346" heatid="9362" lane="4" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:33.78" />
                    <SPLIT distance="150" swimtime="00:02:25.66" />
                    <SPLIT distance="200" swimtime="00:03:19.05" />
                    <SPLIT distance="250" swimtime="00:04:11.48" />
                    <SPLIT distance="300" swimtime="00:05:03.92" />
                    <SPLIT distance="350" swimtime="00:05:56.94" />
                    <SPLIT distance="400" swimtime="00:06:50.42" />
                    <SPLIT distance="450" swimtime="00:07:42.82" />
                    <SPLIT distance="500" swimtime="00:08:35.32" />
                    <SPLIT distance="550" swimtime="00:09:27.34" />
                    <SPLIT distance="600" swimtime="00:10:19.02" />
                    <SPLIT distance="650" swimtime="00:11:10.52" />
                    <SPLIT distance="700" swimtime="00:12:01.45" />
                    <SPLIT distance="750" swimtime="00:12:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6347" heatid="9479" lane="5" entrytime="00:01:28.00" />
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="6348" heatid="9550" lane="2" entrytime="00:03:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="7772" name="niezrzeszony ST">
          <ATHLETES>
            <ATHLETE birthdate="1974-10-05" firstname="Tomasz" gender="M" lastname="Sitkowski" nation="POL" athleteid="7771">
              <RESULTS>
                <RESULT eventid="1195" points="368" reactiontime="+89" swimtime="00:00:29.17" resultid="7773" heatid="9326" lane="2" entrytime="00:00:29.00" />
                <RESULT comment="G3 - Pływak obrócił się na piersi (z wyjątkiem momentu wykonania nawrotu)." eventid="1476" reactiontime="+69" status="DSQ" swimtime="00:00:35.75" resultid="7774" heatid="9452" lane="4" entrytime="00:00:36.60" />
                <RESULT eventid="1544" points="336" reactiontime="+84" swimtime="00:01:07.46" resultid="7775" heatid="9483" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="228" reactiontime="+78" swimtime="00:01:24.82" resultid="7776" heatid="9538" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="217" reactiontime="+68" swimtime="00:03:05.98" resultid="7777" heatid="9588" lane="5" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="8296" name="niezrzeszony SW">
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Witold" gender="M" lastname="Szczechla" nation="POL" athleteid="8295">
              <RESULTS>
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="8297" heatid="9343" lane="5" entrytime="00:03:40.00" />
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="8298" heatid="9507" lane="2" entrytime="00:01:40.00" />
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="8299" heatid="9520" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="8300" heatid="9573" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="5585" status="DNS" swimtime="00:00:00.00" resultid="8301" heatid="9599" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="8705" name="niezrzeszony SW">
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="8704">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="8706" heatid="9322" lane="2" entrytime="00:00:32.30" />
                <RESULT eventid="1314" points="188" reactiontime="+129" swimtime="00:25:19.11" resultid="8707" heatid="9367" lane="5" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:16.70" />
                    <SPLIT distance="200" swimtime="00:04:47.17" />
                    <SPLIT distance="250" swimtime="00:03:55.85" />
                    <SPLIT distance="300" swimtime="00:06:31.60" />
                    <SPLIT distance="350" swimtime="00:05:37.96" />
                    <SPLIT distance="400" swimtime="00:08:15.52" />
                    <SPLIT distance="450" swimtime="00:07:23.44" />
                    <SPLIT distance="500" swimtime="00:11:44.18" />
                    <SPLIT distance="550" swimtime="00:09:07.18" />
                    <SPLIT distance="600" swimtime="00:22:00.71" />
                    <SPLIT distance="650" swimtime="00:10:51.77" />
                    <SPLIT distance="700" swimtime="00:23:42.29" />
                    <SPLIT distance="750" swimtime="00:14:19.68" />
                    <SPLIT distance="850" swimtime="00:16:01.82" />
                    <SPLIT distance="950" swimtime="00:17:43.31" />
                    <SPLIT distance="1050" swimtime="00:21:08.68" />
                    <SPLIT distance="1150" swimtime="00:22:51.79" />
                    <SPLIT distance="1250" swimtime="00:24:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="251" reactiontime="+87" swimtime="00:01:14.29" resultid="8708" heatid="9482" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="201" swimtime="00:06:15.43" resultid="8709" heatid="9617" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:14.11" />
                    <SPLIT distance="200" swimtime="00:03:04.01" />
                    <SPLIT distance="250" swimtime="00:03:53.62" />
                    <SPLIT distance="300" swimtime="00:04:42.92" />
                    <SPLIT distance="350" swimtime="00:05:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="210" reactiontime="+88" swimtime="00:02:51.57" resultid="8710" heatid="9552" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="150" swimtime="00:02:11.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ONE" nation="POL" clubid="6868" name="One Man Team">
          <CONTACT city="Poznań - Daszewice" email="gmo@o2.pl" name="MONCZAK" phone="608639696" zip="61-160" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="6869">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1314" points="463" swimtime="00:18:45.61" resultid="6870" heatid="9365" lane="6" entrytime="00:18:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                    <SPLIT distance="200" swimtime="00:02:25.13" />
                    <SPLIT distance="250" swimtime="00:03:02.33" />
                    <SPLIT distance="300" swimtime="00:03:39.71" />
                    <SPLIT distance="350" swimtime="00:04:17.76" />
                    <SPLIT distance="400" swimtime="00:04:54.99" />
                    <SPLIT distance="450" swimtime="00:05:32.29" />
                    <SPLIT distance="500" swimtime="00:06:10.01" />
                    <SPLIT distance="550" swimtime="00:06:47.67" />
                    <SPLIT distance="600" swimtime="00:07:25.18" />
                    <SPLIT distance="650" swimtime="00:08:03.07" />
                    <SPLIT distance="700" swimtime="00:08:40.67" />
                    <SPLIT distance="750" swimtime="00:09:18.34" />
                    <SPLIT distance="800" swimtime="00:09:56.06" />
                    <SPLIT distance="850" swimtime="00:10:33.73" />
                    <SPLIT distance="900" swimtime="00:11:11.73" />
                    <SPLIT distance="950" swimtime="00:11:49.72" />
                    <SPLIT distance="1000" swimtime="00:12:27.68" />
                    <SPLIT distance="1050" swimtime="00:13:05.64" />
                    <SPLIT distance="1100" swimtime="00:13:43.65" />
                    <SPLIT distance="1150" swimtime="00:14:21.53" />
                    <SPLIT distance="1200" swimtime="00:14:59.65" />
                    <SPLIT distance="1250" swimtime="00:15:37.43" />
                    <SPLIT distance="1300" swimtime="00:16:15.18" />
                    <SPLIT distance="1350" swimtime="00:16:53.12" />
                    <SPLIT distance="1400" swimtime="00:17:31.08" />
                    <SPLIT distance="1450" swimtime="00:18:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6871" heatid="9488" lane="9" entrytime="00:00:59.99" entrycourse="LCM" />
                <RESULT eventid="5399" points="466" reactiontime="+80" swimtime="00:02:11.48" resultid="6872" heatid="9557" lane="2" entrytime="00:02:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:03.79" />
                    <SPLIT distance="150" swimtime="00:01:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="468" reactiontime="+80" swimtime="00:04:43.28" resultid="6873" heatid="9614" lane="5" entrytime="00:04:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:08.90" />
                    <SPLIT distance="150" swimtime="00:01:45.74" />
                    <SPLIT distance="200" swimtime="00:02:21.93" />
                    <SPLIT distance="250" swimtime="00:02:57.97" />
                    <SPLIT distance="300" swimtime="00:03:33.88" />
                    <SPLIT distance="350" swimtime="00:04:09.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PKZA" nation="CZE" clubid="5724" name="Plavecky klub Zabreh">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-26" firstname="David" gender="M" lastname="Kochwasser" nation="CZE" athleteid="5733">
              <RESULTS>
                <RESULT eventid="1195" points="367" reactiontime="+76" swimtime="00:00:29.19" resultid="5734" heatid="9325" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1229" points="285" reactiontime="+76" swimtime="00:02:53.17" resultid="5735" heatid="9345" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="150" swimtime="00:02:11.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="373" reactiontime="+74" swimtime="00:01:05.16" resultid="5736" heatid="9483" lane="4" entrytime="00:01:06.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="322" swimtime="00:01:23.30" resultid="5737" heatid="9510" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="342" reactiontime="+75" swimtime="00:00:32.07" resultid="5738" heatid="9524" lane="0" entrytime="00:00:31.50" />
                <RESULT eventid="5399" points="290" swimtime="00:02:33.95" resultid="5739" heatid="9553" lane="1" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="274" reactiontime="+74" swimtime="00:01:16.62" resultid="5740" heatid="9575" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="375" reactiontime="+70" swimtime="00:00:35.96" resultid="5741" heatid="9602" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-01" firstname="Petr" gender="M" lastname="Horvat" nation="CZE" athleteid="5723">
              <RESULTS>
                <RESULT eventid="1195" points="306" reactiontime="+88" swimtime="00:00:31.02" resultid="5725" heatid="9322" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1476" points="199" reactiontime="+75" swimtime="00:00:41.13" resultid="5727" heatid="9451" lane="7" entrytime="00:00:41.10" />
                <RESULT eventid="1510" points="309" reactiontime="+80" swimtime="00:03:07.26" resultid="5728" heatid="9466" lane="0" entrytime="00:03:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                    <SPLIT distance="150" swimtime="00:02:19.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="274" reactiontime="+81" swimtime="00:00:34.52" resultid="5729" heatid="9521" lane="6" entrytime="00:00:35.20" />
                <RESULT eventid="5399" points="234" reactiontime="+82" swimtime="00:02:45.42" resultid="5730" heatid="9553" lane="8" entrytime="00:02:41.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:03.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="304" reactiontime="+89" swimtime="00:00:38.59" resultid="5731" heatid="9600" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="5636" points="251" reactiontime="+79" swimtime="00:05:48.75" resultid="5732" heatid="9616" lane="0" entrytime="00:05:54.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:07.54" />
                    <SPLIT distance="200" swimtime="00:02:52.23" />
                    <SPLIT distance="250" swimtime="00:03:36.49" />
                    <SPLIT distance="300" swimtime="00:04:21.27" />
                    <SPLIT distance="350" swimtime="00:05:05.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="240" reactiontime="+81" swimtime="00:23:20.21" resultid="9438" heatid="9367" lane="8" late="yes" entrytime="00:23:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:02:10.45" />
                    <SPLIT distance="200" swimtime="00:02:55.86" />
                    <SPLIT distance="250" swimtime="00:03:41.05" />
                    <SPLIT distance="300" swimtime="00:04:26.74" />
                    <SPLIT distance="350" swimtime="00:05:13.03" />
                    <SPLIT distance="400" swimtime="00:05:59.53" />
                    <SPLIT distance="450" swimtime="00:06:45.69" />
                    <SPLIT distance="500" swimtime="00:07:32.32" />
                    <SPLIT distance="550" swimtime="00:08:19.00" />
                    <SPLIT distance="600" swimtime="00:09:06.20" />
                    <SPLIT distance="650" swimtime="00:09:52.65" />
                    <SPLIT distance="700" swimtime="00:10:39.37" />
                    <SPLIT distance="750" swimtime="00:11:25.62" />
                    <SPLIT distance="800" swimtime="00:12:12.80" />
                    <SPLIT distance="850" swimtime="00:12:59.51" />
                    <SPLIT distance="900" swimtime="00:13:47.75" />
                    <SPLIT distance="950" swimtime="00:14:35.79" />
                    <SPLIT distance="1000" swimtime="00:15:23.75" />
                    <SPLIT distance="1050" swimtime="00:16:11.73" />
                    <SPLIT distance="1100" swimtime="00:16:59.77" />
                    <SPLIT distance="1150" swimtime="00:17:47.04" />
                    <SPLIT distance="1200" swimtime="00:18:35.35" />
                    <SPLIT distance="1250" swimtime="00:19:22.98" />
                    <SPLIT distance="1300" swimtime="00:20:11.07" />
                    <SPLIT distance="1350" swimtime="00:20:59.52" />
                    <SPLIT distance="1400" swimtime="00:21:47.32" />
                    <SPLIT distance="1450" swimtime="00:22:34.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-19" firstname="Jiri" gender="M" lastname="Sip" nation="CZE" athleteid="5742">
              <RESULTS>
                <RESULT eventid="1195" points="416" reactiontime="+90" swimtime="00:00:28.01" resultid="5743" heatid="9328" lane="8" entrytime="00:00:27.70" />
                <RESULT eventid="1229" points="383" reactiontime="+93" swimtime="00:02:36.95" resultid="5744" heatid="9347" lane="4" entrytime="00:02:37.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:02:01.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="382" reactiontime="+80" swimtime="00:00:33.12" resultid="5745" heatid="9454" lane="4" entrytime="00:00:33.40" />
                <RESULT eventid="1544" points="473" reactiontime="+87" swimtime="00:01:00.20" resultid="5746" heatid="9487" lane="8" entrytime="00:01:01.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="389" reactiontime="+77" swimtime="00:01:11.02" resultid="5747" heatid="9539" lane="4" entrytime="00:01:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="347" reactiontime="+85" swimtime="00:02:39.18" resultid="5748" heatid="9589" lane="0" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:57.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Jakub" gender="M" lastname="Smid" nation="CZE" athleteid="5749">
              <RESULTS>
                <RESULT eventid="1195" points="473" reactiontime="+84" swimtime="00:00:26.82" resultid="5750" heatid="9328" lane="2" entrytime="00:00:27.40" />
                <RESULT eventid="1229" points="430" reactiontime="+81" swimtime="00:02:30.94" resultid="5751" heatid="9347" lane="5" entrytime="00:02:37.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="495" reactiontime="+77" swimtime="00:00:59.28" resultid="5752" heatid="9486" lane="4" entrytime="00:01:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="494" reactiontime="+80" swimtime="00:01:12.23" resultid="5753" heatid="9512" lane="7" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="420" reactiontime="+80" swimtime="00:00:29.94" resultid="5754" heatid="9526" lane="0" entrytime="00:00:29.40" />
                <RESULT eventid="5585" points="540" reactiontime="+85" swimtime="00:00:31.85" resultid="5755" heatid="9604" lane="7" entrytime="00:00:32.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PREGEL" nation="RUS" clubid="7625" name="Pregel">
          <CONTACT city="Kaliningrad" email="alkonter@gmail.com" name="Pregel" phone="+79062384111" street="Turgeneva 5-9" zip="236008" />
          <ATHLETES>
            <ATHLETE birthdate="1961-10-04" firstname="Dmitriy" gender="M" lastname="Kromskiy" nation="RUS" athleteid="7662">
              <RESULTS>
                <RESULT eventid="1195" points="356" reactiontime="+90" swimtime="00:00:29.50" resultid="7663" heatid="9326" lane="4" entrytime="00:00:28.55" />
                <RESULT eventid="1476" points="290" reactiontime="+83" swimtime="00:00:36.29" resultid="7664" heatid="9454" lane="8" entrytime="00:00:34.60" />
                <RESULT eventid="5365" points="289" reactiontime="+78" swimtime="00:01:18.42" resultid="7665" heatid="9539" lane="9" entrytime="00:01:15.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-04-17" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="7666">
              <RESULTS>
                <RESULT eventid="1229" points="269" swimtime="00:02:56.52" resultid="7667" heatid="9345" lane="6" entrytime="00:02:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:27.98" />
                    <SPLIT distance="150" swimtime="00:02:16.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="271" reactiontime="+72" swimtime="00:22:24.46" resultid="7668" heatid="9366" lane="3" entrytime="00:21:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:26.66" />
                    <SPLIT distance="150" swimtime="00:02:12.31" />
                    <SPLIT distance="200" swimtime="00:02:58.66" />
                    <SPLIT distance="250" swimtime="00:03:44.53" />
                    <SPLIT distance="300" swimtime="00:04:30.71" />
                    <SPLIT distance="350" swimtime="00:05:16.95" />
                    <SPLIT distance="400" swimtime="00:06:03.15" />
                    <SPLIT distance="450" swimtime="00:06:49.19" />
                    <SPLIT distance="500" swimtime="00:07:35.98" />
                    <SPLIT distance="550" swimtime="00:08:21.99" />
                    <SPLIT distance="600" swimtime="00:09:08.22" />
                    <SPLIT distance="650" swimtime="00:09:53.81" />
                    <SPLIT distance="700" swimtime="00:10:39.77" />
                    <SPLIT distance="750" swimtime="00:11:25.27" />
                    <SPLIT distance="800" swimtime="00:12:11.41" />
                    <SPLIT distance="850" swimtime="00:12:56.62" />
                    <SPLIT distance="900" swimtime="00:13:41.13" />
                    <SPLIT distance="950" swimtime="00:14:25.60" />
                    <SPLIT distance="1000" swimtime="00:15:10.29" />
                    <SPLIT distance="1050" swimtime="00:15:54.79" />
                    <SPLIT distance="1100" swimtime="00:16:39.39" />
                    <SPLIT distance="1150" swimtime="00:17:24.38" />
                    <SPLIT distance="1200" swimtime="00:18:09.32" />
                    <SPLIT distance="1250" swimtime="00:18:53.80" />
                    <SPLIT distance="1300" swimtime="00:19:37.94" />
                    <SPLIT distance="1350" swimtime="00:20:21.74" />
                    <SPLIT distance="1400" swimtime="00:21:05.60" />
                    <SPLIT distance="1450" swimtime="00:21:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="275" swimtime="00:01:27.82" resultid="7669" heatid="9509" lane="6" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="308" reactiontime="+65" swimtime="00:02:30.92" resultid="7670" heatid="9553" lane="5" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="324" reactiontime="+71" swimtime="00:00:37.75" resultid="7671" heatid="9601" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="5636" points="308" reactiontime="+66" swimtime="00:05:25.78" resultid="7672" heatid="9616" lane="4" entrytime="00:05:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:01:58.41" />
                    <SPLIT distance="200" swimtime="00:02:40.49" />
                    <SPLIT distance="250" swimtime="00:03:21.83" />
                    <SPLIT distance="300" swimtime="00:04:03.88" />
                    <SPLIT distance="350" swimtime="00:04:45.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-02-11" firstname="Nadezda" gender="F" lastname="Davydova" nation="RUS" athleteid="7632">
              <RESULTS>
                <RESULT eventid="1212" points="249" reactiontime="+102" swimtime="00:03:20.40" resultid="7633" heatid="9338" lane="2" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:36.30" />
                    <SPLIT distance="150" swimtime="00:02:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="312" reactiontime="+106" swimtime="00:01:16.19" resultid="7634" heatid="9472" lane="4" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="208" reactiontime="+118" swimtime="00:00:41.21" resultid="7635" heatid="9515" lane="9" entrytime="00:00:41.50" />
                <RESULT eventid="5382" points="259" swimtime="00:02:57.17" resultid="7636" heatid="9545" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:23.08" />
                    <SPLIT distance="150" swimtime="00:02:10.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="255" swimtime="00:06:12.76" resultid="7637" heatid="9610" lane="1" entrytime="00:06:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="150" swimtime="00:02:11.44" />
                    <SPLIT distance="200" swimtime="00:03:00.17" />
                    <SPLIT distance="250" swimtime="00:03:48.29" />
                    <SPLIT distance="300" swimtime="00:04:37.48" />
                    <SPLIT distance="350" swimtime="00:05:26.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Tatiana" gender="F" lastname="Davydova" nation="RUS" athleteid="7648">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="7649" heatid="9311" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="7650" heatid="9594" lane="3" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-05" firstname="Elena" gender="F" lastname="Mekhteleva" nation="RUS" athleteid="7638">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="7639" heatid="9313" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="7640" heatid="9461" lane="0" entrytime="00:03:10.00" />
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="7641" heatid="9504" lane="2" entrytime="00:01:23.00" />
                <RESULT eventid="5314" status="DNS" swimtime="00:00:00.00" resultid="7642" heatid="9516" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="7643" heatid="9596" lane="7" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-06" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="7626">
              <RESULTS>
                <RESULT eventid="1133" points="291" reactiontime="+99" swimtime="00:00:35.69" resultid="7627" heatid="9311" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="1458" points="218" reactiontime="+84" swimtime="00:00:44.96" resultid="7628" heatid="9442" lane="3" entrytime="00:00:45.50" />
                <RESULT eventid="1527" points="301" swimtime="00:01:17.09" resultid="7629" heatid="9473" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="309" reactiontime="+90" swimtime="00:02:47.11" resultid="7630" heatid="9545" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="150" swimtime="00:02:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="296" reactiontime="+85" swimtime="00:05:54.46" resultid="7631" heatid="9610" lane="2" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:23.74" />
                    <SPLIT distance="150" swimtime="00:02:09.85" />
                    <SPLIT distance="200" swimtime="00:02:55.82" />
                    <SPLIT distance="250" swimtime="00:03:41.47" />
                    <SPLIT distance="300" swimtime="00:04:26.71" />
                    <SPLIT distance="350" swimtime="00:05:11.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="7677" heatid="9353" lane="5" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:00.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7662" number="1" reactiontime="+82" status="DSQ" />
                    <RELAYPOSITION athleteid="7638" number="2" reactiontime="+53" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RMKS " nation="POL" region="SLA" clubid="6575" name="Rmks Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" state="SLA" street="orzepowicka 22a/37" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="6576">
              <RESULTS>
                <RESULT eventid="1133" points="591" reactiontime="+76" swimtime="00:00:28.20" resultid="6577" heatid="9315" lane="2" entrytime="00:00:28.10" />
                <RESULT eventid="1212" points="486" reactiontime="+77" swimtime="00:02:40.37" resultid="6578" heatid="9340" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:02:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="526" swimtime="00:01:04.03" resultid="6579" heatid="9476" lane="9" entrytime="00:01:04.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="543" reactiontime="+74" swimtime="00:00:29.94" resultid="6580" heatid="9517" lane="5" entrytime="00:00:29.58" />
                <RESULT eventid="5499" points="494" reactiontime="+79" swimtime="00:01:10.17" resultid="6581" heatid="9571" lane="5" entrytime="00:01:08.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RSS" nation="POL" clubid="6686" name="Royal Swimmers Ślęza">
          <CONTACT name="Bloch" />
          <ATHLETES>
            <ATHLETE birthdate="1978-07-22" firstname="Magdalena" gender="F" lastname="Antonijczuk-Krzyśków" nation="POL" athleteid="6702">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="6703" heatid="9339" lane="7" entrytime="00:03:07.00" />
                <RESULT eventid="1458" status="DNS" swimtime="00:00:00.00" resultid="6704" heatid="9443" lane="3" entrytime="00:00:40.80" />
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="6705" heatid="9532" lane="0" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-11" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="6693">
              <RESULTS>
                <RESULT eventid="1458" points="262" reactiontime="+81" swimtime="00:00:42.26" resultid="6694" heatid="9443" lane="5" entrytime="00:00:40.80" />
                <RESULT eventid="1527" points="304" swimtime="00:01:16.87" resultid="6695" heatid="9473" lane="6" entrytime="00:01:15.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="226" reactiontime="+88" swimtime="00:00:40.09" resultid="6696" heatid="9515" lane="6" entrytime="00:00:38.24" />
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="6697" heatid="9544" lane="2" entrytime="00:03:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-05-16" firstname="Mariusz" gender="M" lastname="Maciaszek" nation="POL" athleteid="6698">
              <RESULTS>
                <RESULT eventid="1195" points="459" reactiontime="+92" swimtime="00:00:27.10" resultid="6699" heatid="9330" lane="9" entrytime="00:00:26.27" />
                <RESULT eventid="1544" points="456" reactiontime="+90" swimtime="00:01:00.93" resultid="6700" heatid="9486" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="447" reactiontime="+89" swimtime="00:00:29.32" resultid="6701" heatid="9524" lane="4" entrytime="00:00:30.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-07" firstname="Radosław" gender="M" lastname="Stefurak" nation="POL" athleteid="6687">
              <RESULTS>
                <RESULT eventid="1510" points="285" reactiontime="+95" swimtime="00:03:12.46" resultid="6688" heatid="9466" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:01:31.00" />
                    <SPLIT distance="150" swimtime="00:02:21.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="275" reactiontime="+98" swimtime="00:01:27.80" resultid="6689" heatid="9509" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="208" reactiontime="+96" swimtime="00:02:52.03" resultid="6690" heatid="9553" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:05.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="279" reactiontime="+90" swimtime="00:00:39.67" resultid="6691" heatid="9601" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="5636" points="214" swimtime="00:06:07.90" resultid="6692" heatid="9616" lane="1" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:20.94" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                    <SPLIT distance="200" swimtime="00:02:54.35" />
                    <SPLIT distance="250" swimtime="00:03:42.87" />
                    <SPLIT distance="300" swimtime="00:04:32.10" />
                    <SPLIT distance="350" swimtime="00:05:20.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RAAS" nation="POL" clubid="5776" name="Rydułtowska Akademia Aktywnego Seniora" name.en="Rydułtowska Akademia Aktywnego Seniora" shortname="Rydułtowska Akademia Aktywnego" shortname.en="Rydułtowska Akademia Aktywnego">
          <CONTACT name="Marian  Otlik" />
          <ATHLETES>
            <ATHLETE birthdate="1977-08-21" firstname="Michał" gender="M" lastname="Kądzioła" nation="POL" athleteid="5803">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="5804" heatid="9327" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="5805" heatid="9455" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="5806" heatid="9481" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="5807" heatid="9525" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="5808" heatid="9539" lane="7" entrytime="00:01:14.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="5809" heatid="9588" lane="7" entrytime="00:02:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-23" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="5794">
              <RESULTS>
                <RESULT eventid="1229" points="170" swimtime="00:03:25.55" resultid="5795" heatid="9344" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                    <SPLIT distance="100" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:02:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="173" reactiontime="+82" swimtime="00:26:01.36" resultid="5796" heatid="9367" lane="3" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="100" swimtime="00:01:36.48" />
                    <SPLIT distance="150" swimtime="00:02:28.35" />
                    <SPLIT distance="200" swimtime="00:03:20.41" />
                    <SPLIT distance="250" swimtime="00:04:13.86" />
                    <SPLIT distance="300" swimtime="00:05:06.48" />
                    <SPLIT distance="350" swimtime="00:05:59.47" />
                    <SPLIT distance="400" swimtime="00:06:51.36" />
                    <SPLIT distance="450" swimtime="00:07:44.20" />
                    <SPLIT distance="500" swimtime="00:08:35.78" />
                    <SPLIT distance="550" swimtime="00:09:28.56" />
                    <SPLIT distance="600" swimtime="00:10:20.31" />
                    <SPLIT distance="650" swimtime="00:11:12.74" />
                    <SPLIT distance="700" swimtime="00:12:05.27" />
                    <SPLIT distance="750" swimtime="00:12:58.36" />
                    <SPLIT distance="800" swimtime="00:13:51.44" />
                    <SPLIT distance="850" swimtime="00:14:45.00" />
                    <SPLIT distance="900" swimtime="00:15:37.48" />
                    <SPLIT distance="950" swimtime="00:16:30.68" />
                    <SPLIT distance="1000" swimtime="00:17:23.27" />
                    <SPLIT distance="1050" swimtime="00:18:16.01" />
                    <SPLIT distance="1100" swimtime="00:19:08.76" />
                    <SPLIT distance="1150" swimtime="00:20:01.65" />
                    <SPLIT distance="1200" swimtime="00:20:54.55" />
                    <SPLIT distance="1250" swimtime="00:21:46.98" />
                    <SPLIT distance="1300" swimtime="00:22:39.23" />
                    <SPLIT distance="1350" swimtime="00:23:31.05" />
                    <SPLIT distance="1400" swimtime="00:24:21.89" />
                    <SPLIT distance="1450" swimtime="00:25:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="205" reactiontime="+82" swimtime="00:00:40.74" resultid="5797" heatid="9451" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1578" points="91" reactiontime="+98" swimtime="00:04:07.86" resultid="5798" heatid="9494" lane="0" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:55.23" />
                    <SPLIT distance="150" swimtime="00:03:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="153" reactiontime="+80" swimtime="00:01:36.82" resultid="5799" heatid="9536" lane="5" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="142" reactiontime="+100" swimtime="00:07:46.67" resultid="5800" heatid="9565" lane="2" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                    <SPLIT distance="100" swimtime="00:01:54.13" />
                    <SPLIT distance="150" swimtime="00:02:53.93" />
                    <SPLIT distance="200" swimtime="00:03:52.10" />
                    <SPLIT distance="250" swimtime="00:04:59.63" />
                    <SPLIT distance="300" swimtime="00:06:05.91" />
                    <SPLIT distance="350" swimtime="00:06:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="134" reactiontime="+81" swimtime="00:01:37.15" resultid="5801" heatid="9573" lane="3" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="146" reactiontime="+89" swimtime="00:03:32.20" resultid="5802" heatid="9586" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:42.52" />
                    <SPLIT distance="150" swimtime="00:02:38.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="5777">
              <RESULTS>
                <RESULT eventid="1195" points="72" reactiontime="+118" swimtime="00:00:50.12" resultid="5778" heatid="9318" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1229" points="59" reactiontime="+98" swimtime="00:04:52.42" resultid="5779" heatid="9343" lane="8" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.06" />
                    <SPLIT distance="100" swimtime="00:02:26.75" />
                    <SPLIT distance="150" swimtime="00:03:47.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="52" reactiontime="+88" swimtime="00:01:04.18" resultid="5780" heatid="9449" lane="8" entrytime="00:00:55.00" />
                <RESULT eventid="1578" points="22" swimtime="00:06:32.39" resultid="5781" heatid="9493" lane="1" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.50" />
                    <SPLIT distance="100" swimtime="00:03:08.00" />
                    <SPLIT distance="150" swimtime="00:04:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="42" reactiontime="+106" swimtime="00:01:04.31" resultid="5782" heatid="9518" lane="4" entrytime="00:00:59.00" />
                <RESULT eventid="5467" points="50" swimtime="00:11:00.72" resultid="5783" heatid="9564" lane="6" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.94" />
                    <SPLIT distance="100" swimtime="00:02:51.03" />
                    <SPLIT distance="150" swimtime="00:04:16.10" />
                    <SPLIT distance="200" swimtime="00:05:39.35" />
                    <SPLIT distance="250" swimtime="00:07:09.49" />
                    <SPLIT distance="300" swimtime="00:08:35.63" />
                    <SPLIT distance="350" swimtime="00:09:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="30" reactiontime="+97" swimtime="00:02:39.64" resultid="5784" heatid="9572" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="56" reactiontime="+75" swimtime="00:04:50.90" resultid="5785" heatid="9584" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.04" />
                    <SPLIT distance="100" swimtime="00:02:26.89" />
                    <SPLIT distance="150" swimtime="00:03:42.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="5786">
              <RESULTS>
                <RESULT eventid="1195" points="23" reactiontime="+110" swimtime="00:01:12.85" resultid="5787" heatid="9317" lane="3" />
                <RESULT eventid="1476" points="12" reactiontime="+99" swimtime="00:01:44.01" resultid="5788" heatid="9447" lane="3" />
                <RESULT eventid="1544" points="27" reactiontime="+99" swimtime="00:02:35.47" resultid="5789" heatid="9477" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="11" reactiontime="+89" swimtime="00:03:50.98" resultid="5790" heatid="9534" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:50.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="25" swimtime="00:05:46.04" resultid="5791" heatid="9548" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.78" />
                    <SPLIT distance="100" swimtime="00:02:41.74" />
                    <SPLIT distance="150" swimtime="00:04:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="12" reactiontime="+82" swimtime="00:08:03.02" resultid="5792" heatid="9583" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.62" />
                    <SPLIT distance="100" swimtime="00:03:53.02" />
                    <SPLIT distance="150" swimtime="00:05:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="26" swimtime="00:12:21.88" resultid="5793" heatid="9619" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.21" />
                    <SPLIT distance="100" swimtime="00:02:41.11" />
                    <SPLIT distance="150" swimtime="00:04:14.60" />
                    <SPLIT distance="200" swimtime="00:05:49.31" />
                    <SPLIT distance="250" swimtime="00:07:27.36" />
                    <SPLIT distance="300" swimtime="00:09:07.76" />
                    <SPLIT distance="350" swimtime="00:10:48.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIKRET" nation="POL" clubid="5949" name="Sikret Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@tlen.pl" internet="www.sikret-plywanie.pl" name="Zagała Joanna" phone="601427257" state="ŚLĄSK" street="Kościuszki 35" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1940-04-20" firstname="Wojciech" gender="M" lastname="Kosiak" nation="POL" athleteid="5974">
              <RESULTS>
                <RESULT eventid="1195" points="132" reactiontime="+120" swimtime="00:00:41.06" resultid="5975" heatid="9319" lane="0" entrytime="00:00:43.00" />
                <RESULT eventid="1544" points="114" reactiontime="+125" swimtime="00:01:36.72" resultid="5976" heatid="9478" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="59" reactiontime="+118" swimtime="00:00:57.36" resultid="5977" heatid="9519" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="5399" points="91" reactiontime="+119" swimtime="00:03:46.58" resultid="5978" heatid="9549" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:51.22" />
                    <SPLIT distance="150" swimtime="00:02:52.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="5959">
              <RESULTS>
                <RESULT eventid="1133" points="146" reactiontime="+67" swimtime="00:00:44.91" resultid="5960" heatid="9310" lane="1" entrytime="00:00:43.00" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1263" status="DSQ" swimtime="00:00:00.00" resultid="5961" heatid="9356" lane="9" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.53" />
                    <SPLIT distance="100" swimtime="00:01:52.76" />
                    <SPLIT distance="150" swimtime="00:02:55.73" />
                    <SPLIT distance="200" swimtime="00:03:56.79" />
                    <SPLIT distance="250" swimtime="00:04:57.89" />
                    <SPLIT distance="300" swimtime="00:05:58.83" />
                    <SPLIT distance="350" swimtime="00:07:00.44" />
                    <SPLIT distance="400" swimtime="00:08:00.36" />
                    <SPLIT distance="450" swimtime="00:09:01.97" />
                    <SPLIT distance="500" swimtime="00:10:03.57" />
                    <SPLIT distance="550" swimtime="00:11:06.69" />
                    <SPLIT distance="600" swimtime="00:12:05.81" />
                    <SPLIT distance="650" swimtime="00:13:07.18" />
                    <SPLIT distance="700" swimtime="00:14:09.28" />
                    <SPLIT distance="750" swimtime="00:15:11.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="138" swimtime="00:04:28.81" resultid="5962" heatid="9459" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.22" />
                    <SPLIT distance="100" swimtime="00:02:10.28" />
                    <SPLIT distance="150" swimtime="00:03:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M5 - Pływak nie przeniósł ramion do przodu nad lustrem wody." eventid="1561" reactiontime="+93" status="DSQ" swimtime="00:05:57.72" resultid="5963" heatid="9491" lane="5" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.09" />
                    <SPLIT distance="100" swimtime="00:02:25.79" />
                    <SPLIT distance="150" swimtime="00:04:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="93" reactiontime="+95" swimtime="00:00:53.76" resultid="5964" heatid="9514" lane="7" entrytime="00:00:56.00" />
                <RESULT eventid="5382" points="118" swimtime="00:03:49.74" resultid="5965" heatid="9543" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.71" />
                    <SPLIT distance="100" swimtime="00:01:53.01" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="70" reactiontime="+107" swimtime="00:02:14.39" resultid="5966" heatid="9569" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="169" reactiontime="+98" swimtime="00:00:53.09" resultid="5967" heatid="9593" lane="9" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="5950">
              <RESULTS>
                <RESULT eventid="1133" points="227" reactiontime="+77" swimtime="00:00:38.78" resultid="5951" heatid="9310" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1297" points="179" swimtime="00:27:21.84" resultid="5952" heatid="9364" lane="6" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:42.74" />
                    <SPLIT distance="150" swimtime="00:02:38.48" />
                    <SPLIT distance="200" swimtime="00:03:34.67" />
                    <SPLIT distance="250" swimtime="00:04:30.50" />
                    <SPLIT distance="300" swimtime="00:05:26.55" />
                    <SPLIT distance="350" swimtime="00:06:22.26" />
                    <SPLIT distance="400" swimtime="00:07:18.44" />
                    <SPLIT distance="450" swimtime="00:08:13.01" />
                    <SPLIT distance="500" swimtime="00:09:09.09" />
                    <SPLIT distance="550" swimtime="00:10:04.83" />
                    <SPLIT distance="600" swimtime="00:11:01.10" />
                    <SPLIT distance="650" swimtime="00:11:56.28" />
                    <SPLIT distance="700" swimtime="00:12:51.87" />
                    <SPLIT distance="750" swimtime="00:13:47.37" />
                    <SPLIT distance="800" swimtime="00:14:42.92" />
                    <SPLIT distance="850" swimtime="00:15:38.55" />
                    <SPLIT distance="900" swimtime="00:16:34.20" />
                    <SPLIT distance="950" swimtime="00:17:29.86" />
                    <SPLIT distance="1000" swimtime="00:18:25.27" />
                    <SPLIT distance="1050" swimtime="00:19:19.46" />
                    <SPLIT distance="1100" swimtime="00:20:14.12" />
                    <SPLIT distance="1150" swimtime="00:21:08.69" />
                    <SPLIT distance="1200" swimtime="00:22:02.73" />
                    <SPLIT distance="1250" swimtime="00:22:57.04" />
                    <SPLIT distance="1300" swimtime="00:23:50.99" />
                    <SPLIT distance="1350" swimtime="00:24:45.21" />
                    <SPLIT distance="1400" swimtime="00:25:39.19" />
                    <SPLIT distance="1450" swimtime="00:26:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="135" reactiontime="+69" swimtime="00:00:52.69" resultid="5953" heatid="9441" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1527" points="210" reactiontime="+80" swimtime="00:01:26.99" resultid="5954" heatid="9471" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="160" reactiontime="+84" swimtime="00:01:58.01" resultid="5955" heatid="9501" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="192" swimtime="00:03:15.61" resultid="5956" heatid="9544" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:37.10" />
                    <SPLIT distance="150" swimtime="00:02:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="147" reactiontime="+96" swimtime="00:03:54.71" resultid="5957" heatid="9580" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.93" />
                    <SPLIT distance="100" swimtime="00:01:56.83" />
                    <SPLIT distance="150" swimtime="00:02:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="181" reactiontime="+89" swimtime="00:00:51.89" resultid="5958" heatid="9592" lane="7" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="5968">
              <RESULTS>
                <RESULT eventid="1229" points="239" reactiontime="+92" swimtime="00:03:03.53" resultid="5969" heatid="9344" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:23.38" />
                    <SPLIT distance="150" swimtime="00:02:20.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="324" reactiontime="+82" swimtime="00:00:34.97" resultid="5970" heatid="9453" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="5331" points="372" reactiontime="+89" swimtime="00:00:31.17" resultid="5971" heatid="9522" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="5972" heatid="9537" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="5636" points="249" reactiontime="+101" swimtime="00:05:49.75" resultid="5973" heatid="9617" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                    <SPLIT distance="200" swimtime="00:02:48.09" />
                    <SPLIT distance="250" swimtime="00:03:33.00" />
                    <SPLIT distance="300" swimtime="00:04:19.53" />
                    <SPLIT distance="350" swimtime="00:05:06.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1246" reactiontime="+75" status="DSQ" swimtime="00:02:38.12" resultid="5979" heatid="9353" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5959" number="1" reactiontime="+75" status="DSQ" />
                    <RELAYPOSITION athleteid="5974" number="2" reactiontime="+29" status="DSQ" />
                    <RELAYPOSITION athleteid="5950" number="3" reactiontime="+79" status="DSQ" />
                    <RELAYPOSITION athleteid="5968" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5602" status="DNS" swimtime="00:00:00.00" resultid="5980" heatid="9607" lane="0" entrytime="00:02:58.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5950" number="1" />
                    <RELAYPOSITION athleteid="5959" number="2" />
                    <RELAYPOSITION athleteid="5968" number="3" />
                    <RELAYPOSITION athleteid="5974" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STP" nation="POL" clubid="7040" name="St.P.P Legia Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1991-01-17" firstname="Aleksy" gender="M" lastname="Otłowski" nation="POL" athleteid="7039">
              <RESULTS>
                <RESULT eventid="5636" points="448" swimtime="00:04:47.60" resultid="7041" heatid="9613" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:01.51" />
                    <SPLIT distance="150" swimtime="00:01:36.81" />
                    <SPLIT distance="200" swimtime="00:02:14.56" />
                    <SPLIT distance="250" swimtime="00:02:52.76" />
                    <SPLIT distance="300" swimtime="00:03:31.27" />
                    <SPLIT distance="350" swimtime="00:04:10.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STP" nation="POL" clubid="7465" name="START Poznań">
          <CONTACT city="Poznań" email="kaczy4@autograf.pl" name="Kaczmarek" phone="603 434 586" street="Promenada 21" zip="60-375" />
          <ATHLETES>
            <ATHLETE birthdate="1982-10-03" firstname="Michał" gender="M" lastname="Kaczmarek" nation="POL" athleteid="7466">
              <RESULTS>
                <RESULT eventid="1195" points="288" reactiontime="+97" swimtime="00:00:31.66" resultid="7467" heatid="9323" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="7468" heatid="9343" lane="7" entrytime="00:04:00.00" />
                <RESULT eventid="1510" points="263" reactiontime="+106" swimtime="00:03:17.51" resultid="7469" heatid="9465" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:35.95" />
                    <SPLIT distance="150" swimtime="00:02:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="277" reactiontime="+102" swimtime="00:01:11.89" resultid="7470" heatid="9481" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="5297" points="262" reactiontime="+103" swimtime="00:01:29.24" resultid="7471" heatid="9508" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="191" reactiontime="+109" swimtime="00:00:38.89" resultid="7472" heatid="9520" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="5585" points="253" reactiontime="+101" swimtime="00:00:41.01" resultid="7473" heatid="9600" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-06" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="7502">
              <RESULTS>
                <RESULT eventid="1229" points="306" reactiontime="+86" swimtime="00:02:49.15" resultid="7503" heatid="9345" lane="4" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:02:09.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="305" reactiontime="+90" swimtime="00:03:08.12" resultid="7504" heatid="9465" lane="3" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:19.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="245" reactiontime="+90" swimtime="00:02:58.04" resultid="7505" heatid="9494" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="295" reactiontime="+84" swimtime="00:06:06.12" resultid="7506" heatid="9566" lane="3" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                    <SPLIT distance="200" swimtime="00:02:55.08" />
                    <SPLIT distance="250" swimtime="00:03:47.69" />
                    <SPLIT distance="300" swimtime="00:04:39.60" />
                    <SPLIT distance="350" swimtime="00:05:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="247" reactiontime="+86" swimtime="00:01:19.32" resultid="7507" heatid="9575" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-08-09" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="7490">
              <RESULTS>
                <RESULT eventid="1195" points="445" reactiontime="+80" swimtime="00:00:27.37" resultid="7491" heatid="9328" lane="3" entrytime="00:00:27.05" />
                <RESULT eventid="1229" points="401" reactiontime="+79" swimtime="00:02:34.50" resultid="7492" heatid="9348" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="473" reactiontime="+75" swimtime="00:01:00.17" resultid="7493" heatid="9488" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="468" reactiontime="+81" swimtime="00:02:11.34" resultid="7494" heatid="9557" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:04.41" />
                    <SPLIT distance="150" swimtime="00:01:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="379" reactiontime="+83" swimtime="00:05:36.72" resultid="7495" heatid="9567" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                    <SPLIT distance="200" swimtime="00:02:43.36" />
                    <SPLIT distance="250" swimtime="00:03:33.76" />
                    <SPLIT distance="300" swimtime="00:04:23.28" />
                    <SPLIT distance="350" swimtime="00:05:00.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="319" reactiontime="+80" swimtime="00:00:37.97" resultid="7496" heatid="9602" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="5636" points="428" swimtime="00:04:51.92" resultid="7497" heatid="9614" lane="6" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:47.93" />
                    <SPLIT distance="200" swimtime="00:02:26.90" />
                    <SPLIT distance="250" swimtime="00:03:03.47" />
                    <SPLIT distance="300" swimtime="00:03:40.03" />
                    <SPLIT distance="350" swimtime="00:04:16.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-08" firstname="Anna" gender="F" lastname="Rostkowska-Kaczmarek" nation="POL" athleteid="7484">
              <RESULTS>
                <RESULT eventid="1133" points="338" reactiontime="+101" swimtime="00:00:33.95" resultid="7485" heatid="9312" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1527" points="256" reactiontime="+98" swimtime="00:01:21.36" resultid="7486" heatid="9472" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="227" swimtime="00:03:05.09" resultid="7487" heatid="9544" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:30.64" />
                    <SPLIT distance="150" swimtime="00:02:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="238" reactiontime="+106" swimtime="00:00:47.44" resultid="7488" heatid="9594" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="5619" points="213" swimtime="00:06:35.88" resultid="7489" heatid="9611" lane="6" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:31.78" />
                    <SPLIT distance="150" swimtime="00:02:21.63" />
                    <SPLIT distance="200" swimtime="00:03:12.99" />
                    <SPLIT distance="250" swimtime="00:04:04.45" />
                    <SPLIT distance="300" swimtime="00:04:56.01" />
                    <SPLIT distance="350" swimtime="00:05:47.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-08" firstname="Łukasz" gender="M" lastname="Juskowiak" nation="POL" athleteid="7474">
              <RESULTS>
                <RESULT eventid="1195" points="344" reactiontime="+99" swimtime="00:00:29.83" resultid="7475" heatid="9325" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1476" points="211" reactiontime="+68" swimtime="00:00:40.33" resultid="7476" heatid="9454" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1544" points="332" reactiontime="+83" swimtime="00:01:07.70" resultid="7477" heatid="9486" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="295" reactiontime="+91" swimtime="00:00:33.68" resultid="7478" heatid="9524" lane="1" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-03-01" firstname="Adam" gender="M" lastname="Jędrychowski" nation="POL" athleteid="7479">
              <RESULTS>
                <RESULT eventid="1195" points="400" reactiontime="+75" swimtime="00:00:28.37" resultid="7480" heatid="9327" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="5297" points="426" reactiontime="+71" swimtime="00:01:15.91" resultid="7481" heatid="9512" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="346" reactiontime="+79" swimtime="00:00:31.94" resultid="7482" heatid="9524" lane="9" entrytime="00:00:31.50" />
                <RESULT eventid="5585" points="420" reactiontime="+70" swimtime="00:00:34.64" resultid="7483" heatid="9604" lane="0" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-08-03" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="7498">
              <RESULTS>
                <RESULT eventid="1510" points="300" swimtime="00:03:09.21" resultid="7499" heatid="9466" lane="9" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="312" reactiontime="+78" swimtime="00:01:24.17" resultid="7500" heatid="9509" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="325" reactiontime="+87" swimtime="00:00:37.71" resultid="7501" heatid="9601" lane="9" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="5433" status="DNS" swimtime="00:00:00.00" resultid="7508" heatid="9560" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7474" number="1" />
                    <RELAYPOSITION athleteid="7479" number="2" />
                    <RELAYPOSITION athleteid="7502" number="3" />
                    <RELAYPOSITION athleteid="7490" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1612" points="301" reactiontime="+88" swimtime="00:02:19.34" resultid="7509" heatid="9498" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7490" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="7466" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="7474" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="7479" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="5602" status="DNS" swimtime="00:00:00.00" resultid="7510" heatid="9606" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7502" number="1" />
                    <RELAYPOSITION athleteid="7479" number="2" />
                    <RELAYPOSITION athleteid="7490" number="3" />
                    <RELAYPOSITION athleteid="7484" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1246" status="DNS" swimtime="00:00:00.00" resultid="7511" heatid="9353" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7490" number="1" />
                    <RELAYPOSITION athleteid="7484" number="2" />
                    <RELAYPOSITION athleteid="7502" number="3" />
                    <RELAYPOSITION athleteid="7479" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="6333" name="Steef Wrocław">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="6334">
              <RESULTS>
                <RESULT eventid="1212" points="272" reactiontime="+84" swimtime="00:03:14.47" resultid="6335" heatid="9339" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="260" reactiontime="+94" swimtime="00:24:08.78" resultid="6336" heatid="9364" lane="5" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:02:17.90" />
                    <SPLIT distance="200" swimtime="00:03:06.33" />
                    <SPLIT distance="250" swimtime="00:03:56.38" />
                    <SPLIT distance="300" swimtime="00:04:45.20" />
                    <SPLIT distance="350" swimtime="00:05:33.62" />
                    <SPLIT distance="400" swimtime="00:06:22.75" />
                    <SPLIT distance="450" swimtime="00:07:11.21" />
                    <SPLIT distance="500" swimtime="00:07:59.99" />
                    <SPLIT distance="550" swimtime="00:08:48.10" />
                    <SPLIT distance="600" swimtime="00:09:37.10" />
                    <SPLIT distance="650" swimtime="00:10:25.50" />
                    <SPLIT distance="700" swimtime="00:11:14.55" />
                    <SPLIT distance="750" swimtime="00:12:03.69" />
                    <SPLIT distance="800" swimtime="00:12:52.58" />
                    <SPLIT distance="850" swimtime="00:13:41.58" />
                    <SPLIT distance="900" swimtime="00:14:30.38" />
                    <SPLIT distance="950" swimtime="00:15:19.08" />
                    <SPLIT distance="1000" swimtime="00:16:08.70" />
                    <SPLIT distance="1050" swimtime="00:16:56.93" />
                    <SPLIT distance="1100" swimtime="00:17:45.31" />
                    <SPLIT distance="1150" swimtime="00:18:33.98" />
                    <SPLIT distance="1200" swimtime="00:19:22.68" />
                    <SPLIT distance="1250" swimtime="00:20:10.60" />
                    <SPLIT distance="1300" swimtime="00:20:58.58" />
                    <SPLIT distance="1350" swimtime="00:21:46.76" />
                    <SPLIT distance="1400" swimtime="00:22:34.84" />
                    <SPLIT distance="1450" swimtime="00:23:22.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="278" reactiontime="+90" swimtime="00:00:41.44" resultid="6337" heatid="9443" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1561" status="DNS" swimtime="00:00:00.00" resultid="6338" heatid="9492" lane="8" entrytime="00:03:30.00" />
                <RESULT eventid="5348" points="273" reactiontime="+81" swimtime="00:01:29.50" resultid="6339" heatid="9532" lane="8" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="269" swimtime="00:06:52.30" resultid="6340" heatid="9563" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="100" swimtime="00:01:37.31" />
                    <SPLIT distance="150" swimtime="00:02:29.23" />
                    <SPLIT distance="200" swimtime="00:03:19.26" />
                    <SPLIT distance="250" swimtime="00:04:17.92" />
                    <SPLIT distance="300" swimtime="00:05:16.19" />
                    <SPLIT distance="350" swimtime="00:06:05.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="290" reactiontime="+80" swimtime="00:03:07.37" resultid="6341" heatid="9581" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                    <SPLIT distance="150" swimtime="00:02:18.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="251" swimtime="00:06:14.44" resultid="6342" heatid="9610" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:18.26" />
                    <SPLIT distance="200" swimtime="00:03:06.67" />
                    <SPLIT distance="250" swimtime="00:03:55.34" />
                    <SPLIT distance="300" swimtime="00:04:43.77" />
                    <SPLIT distance="350" swimtime="00:05:31.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STR" nation="POL" clubid="6861" name="Swim Tri Rzeszów">
          <CONTACT city="RZESZÓW" email="KLUB@SWIMTRI.PL" name="SWIM TRI RZESZÓW" street="KS. JERZEGO POPIEŁUSZKI 26 C" zip="35-328" />
          <ATHLETES>
            <ATHLETE birthdate="1963-11-15" firstname="Mariusz" gender="M" lastname="Faff" nation="POL" athleteid="6862">
              <RESULTS>
                <RESULT eventid="1195" points="373" reactiontime="+90" swimtime="00:00:29.03" resultid="6863" heatid="9325" lane="7" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1476" points="289" reactiontime="+78" swimtime="00:00:36.32" resultid="6864" heatid="9453" lane="1" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="373" reactiontime="+85" swimtime="00:01:05.16" resultid="6865" heatid="9485" lane="5" entrytime="00:01:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="327" reactiontime="+97" swimtime="00:00:32.55" resultid="6866" heatid="9523" lane="4" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="5399" points="310" swimtime="00:02:30.67" resultid="6867" heatid="9554" lane="1" entrytime="00:02:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMTS" nation="POL" clubid="8533" name="Swimming Masters Team Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="8560">
              <RESULTS>
                <RESULT eventid="1493" points="335" reactiontime="+93" swimtime="00:03:20.14" resultid="8561" heatid="9460" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:34.77" />
                    <SPLIT distance="150" swimtime="00:02:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="8562" heatid="9502" lane="2" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="8545">
              <RESULTS>
                <RESULT eventid="1195" points="500" reactiontime="+81" swimtime="00:00:26.34" resultid="8546" heatid="9329" lane="4" entrytime="00:00:26.30" />
                <RESULT eventid="1476" points="425" reactiontime="+77" swimtime="00:00:31.97" resultid="8547" heatid="9452" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1544" points="522" reactiontime="+81" swimtime="00:00:58.25" resultid="8548" heatid="9487" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="440" reactiontime="+84" swimtime="00:00:29.48" resultid="8549" heatid="9524" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="5365" points="382" reactiontime="+86" swimtime="00:01:11.43" resultid="8550" heatid="9539" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="409" reactiontime="+80" swimtime="00:01:07.11" resultid="8551" heatid="9576" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="366" reactiontime="+86" swimtime="00:00:36.26" resultid="8552" heatid="9601" lane="8" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-09-22" firstname="Szymon" gender="M" lastname="Zabawa" nation="POL" athleteid="8589">
              <RESULTS>
                <RESULT eventid="1476" points="410" reactiontime="+68" swimtime="00:00:32.35" resultid="8590" heatid="9452" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1544" points="456" reactiontime="+70" swimtime="00:01:00.92" resultid="8591" heatid="9487" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="8592" heatid="9540" lane="7" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="8571">
              <RESULTS>
                <RESULT eventid="5551" points="139" reactiontime="+82" swimtime="00:03:35.59" resultid="8572" heatid="9587" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:40.96" />
                    <SPLIT distance="150" swimtime="00:02:38.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-26" firstname="Grzegorz" gender="M" lastname="Król" nation="POL" athleteid="8556">
              <RESULTS>
                <RESULT eventid="1544" points="189" reactiontime="+100" swimtime="00:01:21.73" resultid="8557" heatid="9479" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="153" reactiontime="+99" swimtime="00:03:10.34" resultid="8558" heatid="9551" lane="0" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="150" swimtime="00:02:21.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="149" reactiontime="+104" swimtime="00:06:55.11" resultid="8559" heatid="9619" lane="5" entrytime="00:07:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:36.59" />
                    <SPLIT distance="150" swimtime="00:02:30.14" />
                    <SPLIT distance="200" swimtime="00:03:24.96" />
                    <SPLIT distance="250" swimtime="00:04:19.41" />
                    <SPLIT distance="300" swimtime="00:05:12.04" />
                    <SPLIT distance="350" swimtime="00:06:05.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="8534">
              <RESULTS>
                <RESULT eventid="1133" points="524" reactiontime="+86" swimtime="00:00:29.35" resultid="8535" heatid="9314" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1458" points="540" reactiontime="+80" swimtime="00:00:33.22" resultid="8536" heatid="9446" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="5348" points="521" reactiontime="+74" swimtime="00:01:12.20" resultid="8537" heatid="9533" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="283" reactiontime="+91" swimtime="00:00:44.77" resultid="8538" heatid="9595" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-12" firstname="Łukasz" gender="M" lastname="Rożek" nation="POL" athleteid="8581">
              <RESULTS>
                <RESULT eventid="1195" points="239" reactiontime="+89" swimtime="00:00:33.69" resultid="8582" heatid="9322" lane="0" entrytime="00:00:32.87" />
                <RESULT eventid="1314" reactiontime="+90" status="OTL" swimtime="00:00:00.00" resultid="8583" heatid="9367" lane="2" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                    <SPLIT distance="100" swimtime="00:01:37.43" />
                    <SPLIT distance="150" swimtime="00:02:31.82" />
                    <SPLIT distance="200" swimtime="00:03:27.34" />
                    <SPLIT distance="250" swimtime="00:04:22.84" />
                    <SPLIT distance="300" swimtime="00:05:18.95" />
                    <SPLIT distance="350" swimtime="00:06:16.24" />
                    <SPLIT distance="400" swimtime="00:07:13.00" />
                    <SPLIT distance="450" swimtime="00:08:09.79" />
                    <SPLIT distance="500" swimtime="00:09:08.31" />
                    <SPLIT distance="550" swimtime="00:10:05.97" />
                    <SPLIT distance="600" swimtime="00:11:04.44" />
                    <SPLIT distance="650" swimtime="00:12:02.17" />
                    <SPLIT distance="700" swimtime="00:12:59.86" />
                    <SPLIT distance="750" swimtime="00:13:56.00" />
                    <SPLIT distance="800" swimtime="00:14:53.41" />
                    <SPLIT distance="850" swimtime="00:15:51.34" />
                    <SPLIT distance="900" swimtime="00:16:47.75" />
                    <SPLIT distance="950" swimtime="00:17:44.53" />
                    <SPLIT distance="1000" swimtime="00:18:41.22" />
                    <SPLIT distance="1050" swimtime="00:19:39.70" />
                    <SPLIT distance="1100" swimtime="00:20:37.67" />
                    <SPLIT distance="1150" swimtime="00:21:36.68" />
                    <SPLIT distance="1200" swimtime="00:22:27.80" />
                    <SPLIT distance="1300" swimtime="00:22:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="218" swimtime="00:01:17.91" resultid="8584" heatid="9481" lane="9" entrytime="00:01:18.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="8585" heatid="9519" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="5399" points="171" reactiontime="+88" swimtime="00:03:03.46" resultid="8586" heatid="9551" lane="4" entrytime="00:02:58.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="152" reactiontime="+94" swimtime="00:00:48.52" resultid="8587" heatid="9598" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="5636" points="144" reactiontime="+89" swimtime="00:06:59.66" resultid="8588" heatid="9618" lane="7" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:33.74" />
                    <SPLIT distance="150" swimtime="00:02:26.94" />
                    <SPLIT distance="200" swimtime="00:03:21.44" />
                    <SPLIT distance="250" swimtime="00:04:17.57" />
                    <SPLIT distance="300" swimtime="00:05:13.57" />
                    <SPLIT distance="350" swimtime="00:06:09.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-29" firstname="Robert" gender="M" lastname="Szota" nation="POL" athleteid="8596">
              <RESULTS>
                <RESULT eventid="1195" points="337" reactiontime="+71" swimtime="00:00:30.02" resultid="8597" heatid="9324" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1280" points="318" swimtime="00:11:02.05" resultid="8598" heatid="9360" lane="6" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                    <SPLIT distance="200" swimtime="00:02:35.22" />
                    <SPLIT distance="250" swimtime="00:03:16.83" />
                    <SPLIT distance="300" swimtime="00:03:59.12" />
                    <SPLIT distance="350" swimtime="00:04:41.22" />
                    <SPLIT distance="400" swimtime="00:05:23.41" />
                    <SPLIT distance="450" swimtime="00:06:05.67" />
                    <SPLIT distance="500" swimtime="00:06:48.22" />
                    <SPLIT distance="550" swimtime="00:07:30.70" />
                    <SPLIT distance="600" swimtime="00:08:13.04" />
                    <SPLIT distance="650" swimtime="00:08:55.78" />
                    <SPLIT distance="700" swimtime="00:09:38.68" />
                    <SPLIT distance="750" swimtime="00:10:21.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="233" reactiontime="+72" swimtime="00:00:39.02" resultid="8599" heatid="9451" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1544" points="357" swimtime="00:01:06.07" resultid="8600" heatid="9484" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-13" firstname="Bogusław" gender="M" lastname="Michalak" nation="POL" athleteid="8593">
              <RESULTS>
                <RESULT eventid="1476" points="60" reactiontime="+106" swimtime="00:01:01.09" resultid="8594" heatid="9447" lane="8" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="8595" heatid="9534" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-27" firstname="Marek" gender="M" lastname="Piotrowski" nation="POL" athleteid="8553">
              <RESULTS>
                <RESULT eventid="5399" points="248" reactiontime="+76" swimtime="00:02:42.19" resultid="8554" heatid="9552" lane="7" entrytime="00:02:50.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="240" reactiontime="+76" swimtime="00:05:54.00" resultid="8555" heatid="9617" lane="3" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:02.05" />
                    <SPLIT distance="200" swimtime="00:02:47.37" />
                    <SPLIT distance="250" swimtime="00:03:33.55" />
                    <SPLIT distance="300" swimtime="00:04:20.55" />
                    <SPLIT distance="350" swimtime="00:05:08.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="8539">
              <RESULTS>
                <RESULT eventid="1195" points="414" reactiontime="+90" swimtime="00:00:28.04" resultid="8540" heatid="9324" lane="9" entrytime="00:00:30.02" />
                <RESULT eventid="1544" points="402" swimtime="00:01:03.56" resultid="8541" heatid="9484" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="341" swimtime="00:01:21.75" resultid="8542" heatid="9511" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="8543" heatid="9574" lane="5" entrytime="00:01:22.00" />
                <RESULT eventid="5585" points="389" reactiontime="+80" swimtime="00:00:35.53" resultid="8544" heatid="9603" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="8563">
              <RESULTS>
                <RESULT eventid="1212" points="415" reactiontime="+75" swimtime="00:02:49.00" resultid="8564" heatid="9340" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:02:09.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="369" swimtime="00:11:15.68" resultid="8565" heatid="9355" lane="1" entrytime="00:11:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                    <SPLIT distance="200" swimtime="00:02:43.33" />
                    <SPLIT distance="250" swimtime="00:03:26.63" />
                    <SPLIT distance="300" swimtime="00:04:10.49" />
                    <SPLIT distance="350" swimtime="00:04:54.28" />
                    <SPLIT distance="400" swimtime="00:05:38.07" />
                    <SPLIT distance="450" swimtime="00:06:21.70" />
                    <SPLIT distance="500" swimtime="00:07:05.53" />
                    <SPLIT distance="550" swimtime="00:07:48.68" />
                    <SPLIT distance="600" swimtime="00:08:31.89" />
                    <SPLIT distance="650" swimtime="00:09:14.14" />
                    <SPLIT distance="700" swimtime="00:09:56.29" />
                    <SPLIT distance="750" swimtime="00:10:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="387" reactiontime="+79" swimtime="00:00:37.11" resultid="8566" heatid="9445" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1527" points="428" reactiontime="+70" swimtime="00:01:08.57" resultid="8567" heatid="9475" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="393" reactiontime="+87" swimtime="00:01:19.29" resultid="8568" heatid="9533" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="394" swimtime="00:02:34.11" resultid="8569" heatid="9547" lane="9" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5534" points="400" reactiontime="+80" swimtime="00:02:48.27" resultid="8570" heatid="9582" lane="7" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:21.76" />
                    <SPLIT distance="150" swimtime="00:02:05.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="8573">
              <RESULTS>
                <RESULT eventid="1195" points="315" reactiontime="+77" swimtime="00:00:30.73" resultid="8574" heatid="9323" lane="5" entrytime="00:00:30.20" />
                <RESULT eventid="1229" points="215" reactiontime="+69" swimtime="00:03:10.12" resultid="8575" heatid="9344" lane="2" entrytime="00:03:11.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="150" swimtime="00:02:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="286" reactiontime="+73" swimtime="00:01:11.14" resultid="8576" heatid="9482" lane="2" entrytime="00:01:10.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="294" reactiontime="+72" swimtime="00:00:33.71" resultid="8577" heatid="9522" lane="0" entrytime="00:00:33.80" />
                <RESULT eventid="5399" points="227" reactiontime="+88" swimtime="00:02:46.98" resultid="8578" heatid="9552" lane="3" entrytime="00:02:47.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:03.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="250" swimtime="00:01:19.06" resultid="8579" heatid="9576" lane="1" entrytime="00:01:10.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="297" reactiontime="+81" swimtime="00:00:38.86" resultid="8580" heatid="9600" lane="5" entrytime="00:00:38.78" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="SMT Szczecin 1" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="371" reactiontime="+75" swimtime="00:02:10.02" resultid="8601" heatid="9498" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:40.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8545" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="8539" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="8573" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="8596" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5433" points="290" swimtime="00:02:08.09" resultid="8602" heatid="9561" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="100" swimtime="00:01:03.54" />
                    <SPLIT distance="150" swimtime="00:01:40.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8573" number="1" />
                    <RELAYPOSITION athleteid="8581" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="8556" number="3" />
                    <RELAYPOSITION athleteid="8539" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT Szczecin 1" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+87" swimtime="00:02:08.75" resultid="8603" heatid="9608" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:42.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8534" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="8539" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="8563" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="8545" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STP MASTER" nation="POL" region="ZAC" clubid="5932" name="Szczecineckie TP Masters">
          <CONTACT city="Szczecinek" email="szczecinekmasters@wp.pl" name="Wojnicz Andrzej" phone="887550761" state="ZACHO" street="Szczecińska" zip="78-400" />
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="5933">
              <RESULTS>
                <RESULT eventid="1195" points="54" swimtime="00:00:55.31" resultid="5934" heatid="9318" lane="9" entrytime="00:01:01.00" entrycourse="SCM" />
                <RESULT eventid="1280" points="51" swimtime="00:20:17.03" resultid="5935" heatid="9363" lane="3" entrytime="00:20:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.74" />
                    <SPLIT distance="100" swimtime="00:02:15.15" />
                    <SPLIT distance="150" swimtime="00:03:13.82" />
                    <SPLIT distance="200" swimtime="00:04:43.12" />
                    <SPLIT distance="250" swimtime="00:05:57.80" />
                    <SPLIT distance="300" swimtime="00:07:13.14" />
                    <SPLIT distance="350" swimtime="00:08:27.56" />
                    <SPLIT distance="400" swimtime="00:09:45.40" />
                    <SPLIT distance="450" swimtime="00:11:01.29" />
                    <SPLIT distance="500" swimtime="00:12:19.86" />
                    <SPLIT distance="550" swimtime="00:13:37.59" />
                    <SPLIT distance="600" swimtime="00:14:55.62" />
                    <SPLIT distance="650" swimtime="00:16:14.35" />
                    <SPLIT distance="700" swimtime="00:17:35.35" />
                    <SPLIT distance="750" swimtime="00:18:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="48" reactiontime="+133" swimtime="00:01:06.08" resultid="5936" heatid="9448" lane="9" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1544" points="55" swimtime="00:02:03.32" resultid="5937" heatid="9477" lane="3" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="38" reactiontime="+119" swimtime="00:02:33.33" resultid="5938" heatid="9534" lane="5" entrytime="00:02:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="50" swimtime="00:04:36.84" resultid="5939" heatid="9549" lane="9" entrytime="00:04:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.27" />
                    <SPLIT distance="100" swimtime="00:02:14.64" />
                    <SPLIT distance="150" swimtime="00:03:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="35" reactiontime="+123" swimtime="00:05:39.28" resultid="5940" heatid="9584" lane="9" entrytime="00:05:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.95" />
                    <SPLIT distance="100" swimtime="00:02:43.84" />
                    <SPLIT distance="150" swimtime="00:04:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="53" swimtime="00:09:45.36" resultid="5941" heatid="9619" lane="8" entrytime="00:09:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.84" />
                    <SPLIT distance="100" swimtime="00:02:23.09" />
                    <SPLIT distance="150" swimtime="00:03:34.91" />
                    <SPLIT distance="200" swimtime="00:04:50.40" />
                    <SPLIT distance="250" swimtime="00:06:04.46" />
                    <SPLIT distance="300" swimtime="00:07:19.71" />
                    <SPLIT distance="350" swimtime="00:08:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MO" nation="POL" clubid="6132" name="T.P.Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Samsel" nation="POL" athleteid="6145">
              <RESULTS>
                <RESULT eventid="1195" points="531" reactiontime="+72" swimtime="00:00:25.82" resultid="6146" heatid="9330" lane="4" entrytime="00:00:25.60" />
                <RESULT eventid="1476" points="399" reactiontime="+74" swimtime="00:00:32.64" resultid="6147" heatid="9455" lane="4" entrytime="00:00:31.76" />
                <RESULT eventid="1544" points="524" reactiontime="+72" swimtime="00:00:58.17" resultid="6148" heatid="9489" lane="5" entrytime="00:00:56.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="6149" heatid="9526" lane="8" entrytime="00:00:29.40" />
                <RESULT eventid="5365" points="348" reactiontime="+66" swimtime="00:01:13.65" resultid="6150" heatid="9540" lane="6" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="337" reactiontime="+72" swimtime="00:02:40.76" resultid="6151" heatid="9589" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:01:59.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="6133">
              <RESULTS>
                <RESULT eventid="5467" points="502" reactiontime="+69" swimtime="00:05:06.72" resultid="6134" heatid="9568" lane="8" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                    <SPLIT distance="200" swimtime="00:02:30.91" />
                    <SPLIT distance="250" swimtime="00:03:11.40" />
                    <SPLIT distance="300" swimtime="00:03:53.50" />
                    <SPLIT distance="350" swimtime="00:04:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="469" reactiontime="+67" swimtime="00:02:24.01" resultid="6135" heatid="9590" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="489" reactiontime="+79" swimtime="00:04:39.27" resultid="6136" heatid="9614" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:04.97" />
                    <SPLIT distance="150" swimtime="00:01:39.80" />
                    <SPLIT distance="200" swimtime="00:02:17.01" />
                    <SPLIT distance="250" swimtime="00:02:52.40" />
                    <SPLIT distance="300" swimtime="00:03:29.40" />
                    <SPLIT distance="350" swimtime="00:04:04.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="6152">
              <RESULTS>
                <RESULT eventid="1195" points="420" reactiontime="+72" swimtime="00:00:27.91" resultid="6153" heatid="9328" lane="0" entrytime="00:00:27.91" />
                <RESULT comment="Czas Lepszy od Rekordu Polski Kat. G" eventid="1476" points="459" reactiontime="+73" swimtime="00:00:31.16" resultid="6154" heatid="9456" lane="8" entrytime="00:00:31.27" />
                <RESULT eventid="5365" points="442" reactiontime="+63" swimtime="00:01:08.03" resultid="6155" heatid="9541" lane="9" entrytime="00:01:07.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski/ Czas lepszy od Rekordu Europy" eventid="5551" points="442" reactiontime="+66" swimtime="00:02:26.90" resultid="6156" heatid="9590" lane="7" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:49.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="6137">
              <RESULTS>
                <RESULT eventid="1195" points="104" reactiontime="+128" swimtime="00:00:44.35" resultid="6138" heatid="9318" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1476" points="55" reactiontime="+98" swimtime="00:01:02.88" resultid="6139" heatid="9448" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="1544" points="51" reactiontime="+116" swimtime="00:02:06.08" resultid="6140" heatid="9478" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="40" reactiontime="+91" swimtime="00:02:30.56" resultid="6141" heatid="9535" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="6142" heatid="9550" lane="0" entrytime="00:03:45.00" />
                <RESULT eventid="5551" points="31" reactiontime="+92" swimtime="00:05:56.11" resultid="6143" heatid="9583" lane="4" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.31" />
                    <SPLIT distance="100" swimtime="00:02:54.21" />
                    <SPLIT distance="150" swimtime="00:04:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="33" reactiontime="+122" swimtime="00:01:20.23" resultid="6144" heatid="9597" lane="5" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="6157">
              <RESULTS>
                <RESULT eventid="1133" points="514" reactiontime="+82" swimtime="00:00:29.53" resultid="6158" heatid="9314" lane="7" entrytime="00:00:30.22" />
                <RESULT eventid="1458" points="569" reactiontime="+71" swimtime="00:00:32.65" resultid="6159" heatid="9446" lane="7" entrytime="00:00:33.14" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5348" points="567" reactiontime="+65" swimtime="00:01:10.16" resultid="6160" heatid="9533" lane="4" entrytime="00:01:10.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5534" points="526" reactiontime="+68" swimtime="00:02:33.59" resultid="6161" heatid="9582" lane="4" entrytime="00:02:31.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4215" nation="POL" region="PO" clubid="7055" name="Tarnowskie Termy">
          <CONTACT email="damiandelfin@o2.pl" name="Jerszyński" phone="500276047" />
          <ATHLETES>
            <ATHLETE birthdate="1992-06-14" firstname="Alicja" gender="F" lastname="Szwarc" nation="POL" athleteid="7056">
              <RESULTS>
                <RESULT eventid="1263" points="346" reactiontime="+72" swimtime="00:11:30.34" resultid="7057" heatid="9355" lane="3" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:54.38" />
                    <SPLIT distance="200" swimtime="00:02:36.21" />
                    <SPLIT distance="250" swimtime="00:03:18.39" />
                    <SPLIT distance="300" swimtime="00:04:01.76" />
                    <SPLIT distance="350" swimtime="00:04:46.12" />
                    <SPLIT distance="400" swimtime="00:05:30.84" />
                    <SPLIT distance="450" swimtime="00:06:15.52" />
                    <SPLIT distance="500" swimtime="00:06:59.97" />
                    <SPLIT distance="550" swimtime="00:07:45.23" />
                    <SPLIT distance="600" swimtime="00:08:30.82" />
                    <SPLIT distance="650" swimtime="00:09:16.30" />
                    <SPLIT distance="700" swimtime="00:10:01.27" />
                    <SPLIT distance="750" swimtime="00:10:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="381" reactiontime="+70" swimtime="00:02:47.93" resultid="7058" heatid="9492" lane="5" entrytime="00:02:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:02.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="418" reactiontime="+68" swimtime="00:02:31.00" resultid="7059" heatid="9546" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-12-27" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="7060">
              <RESULTS>
                <RESULT eventid="1133" points="544" reactiontime="+74" swimtime="00:00:28.99" resultid="7061" heatid="9314" lane="4" entrytime="00:00:29.33" />
                <RESULT eventid="1458" points="527" reactiontime="+76" swimtime="00:00:33.50" resultid="7062" heatid="9446" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="5314" points="497" reactiontime="+76" swimtime="00:00:30.84" resultid="7063" heatid="9517" lane="2" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-07-08" firstname="Tomasz" gender="M" lastname="Rybak" nation="POL" athleteid="7068">
              <RESULTS>
                <RESULT eventid="1195" points="389" reactiontime="+84" swimtime="00:00:28.63" resultid="7069" heatid="9327" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="5331" points="403" reactiontime="+76" swimtime="00:00:30.36" resultid="7070" heatid="9524" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-05-24" firstname="Bartosz" gender="M" lastname="Jaraszkiewicz" nation="POL" athleteid="7064">
              <RESULTS>
                <RESULT eventid="1476" points="558" reactiontime="+61" swimtime="00:00:29.19" resultid="7065" heatid="9457" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="5365" points="546" reactiontime="+61" swimtime="00:01:03.42" resultid="7066" heatid="9541" lane="3" entrytime="00:01:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="500" reactiontime="+56" swimtime="00:02:20.98" resultid="7067" heatid="9590" lane="4" entrytime="00:02:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:44.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+55" swimtime="00:02:08.79" resultid="7072" heatid="9606" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:40.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7064" number="1" reactiontime="+55" />
                    <RELAYPOSITION athleteid="7060" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7056" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7068" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TKKF" nation="POL" region="ZAC" clubid="7798" name="TKKF Koszalin Masters">
          <CONTACT email="rpieslak@wp.pl" name="Pieślak Roman" phone="600227112" />
          <ATHLETES>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="7836">
              <RESULTS>
                <RESULT eventid="1195" points="362" reactiontime="+99" swimtime="00:00:29.32" resultid="7837" heatid="9327" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="1544" points="361" reactiontime="+78" swimtime="00:01:05.83" resultid="7838" heatid="9485" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="299" reactiontime="+83" swimtime="00:00:33.51" resultid="7839" heatid="9523" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="7846">
              <RESULTS>
                <RESULT eventid="1297" points="212" reactiontime="+101" swimtime="00:25:50.69" resultid="7847" heatid="9364" lane="3" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="150" swimtime="00:02:25.91" />
                    <SPLIT distance="200" swimtime="00:03:18.40" />
                    <SPLIT distance="250" swimtime="00:04:10.77" />
                    <SPLIT distance="300" swimtime="00:05:03.46" />
                    <SPLIT distance="350" swimtime="00:05:55.86" />
                    <SPLIT distance="400" swimtime="00:06:48.00" />
                    <SPLIT distance="450" swimtime="00:07:40.27" />
                    <SPLIT distance="500" swimtime="00:08:32.56" />
                    <SPLIT distance="550" swimtime="00:09:24.66" />
                    <SPLIT distance="600" swimtime="00:10:16.62" />
                    <SPLIT distance="650" swimtime="00:10:58.63" />
                    <SPLIT distance="700" swimtime="00:12:00.90" />
                    <SPLIT distance="750" swimtime="00:12:52.78" />
                    <SPLIT distance="800" swimtime="00:13:44.22" />
                    <SPLIT distance="850" swimtime="00:14:35.94" />
                    <SPLIT distance="900" swimtime="00:15:27.63" />
                    <SPLIT distance="950" swimtime="00:16:19.90" />
                    <SPLIT distance="1000" swimtime="00:17:11.82" />
                    <SPLIT distance="1050" swimtime="00:18:04.00" />
                    <SPLIT distance="1100" swimtime="00:18:56.40" />
                    <SPLIT distance="1150" swimtime="00:19:49.16" />
                    <SPLIT distance="1200" swimtime="00:20:40.97" />
                    <SPLIT distance="1250" swimtime="00:21:33.57" />
                    <SPLIT distance="1300" swimtime="00:22:25.25" />
                    <SPLIT distance="1350" swimtime="00:23:16.87" />
                    <SPLIT distance="1400" swimtime="00:24:08.22" />
                    <SPLIT distance="1450" swimtime="00:25:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="175" reactiontime="+79" swimtime="00:00:48.33" resultid="7848" heatid="9442" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1527" points="196" swimtime="00:01:28.87" resultid="7849" heatid="9472" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="159" reactiontime="+98" swimtime="00:01:58.31" resultid="7850" heatid="9502" lane="0" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="202" reactiontime="+100" swimtime="00:07:33.93" resultid="7851" heatid="9562" lane="3" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:48.32" />
                    <SPLIT distance="150" swimtime="00:02:45.81" />
                    <SPLIT distance="200" swimtime="00:03:42.00" />
                    <SPLIT distance="250" swimtime="00:04:46.32" />
                    <SPLIT distance="300" swimtime="00:05:52.22" />
                    <SPLIT distance="350" swimtime="00:06:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="177" reactiontime="+70" swimtime="00:03:40.64" resultid="7852" heatid="9580" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.58" />
                    <SPLIT distance="100" swimtime="00:01:48.12" />
                    <SPLIT distance="150" swimtime="00:02:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="197" reactiontime="+99" swimtime="00:06:45.71" resultid="7853" heatid="9611" lane="4" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:34.35" />
                    <SPLIT distance="150" swimtime="00:02:25.87" />
                    <SPLIT distance="200" swimtime="00:03:17.74" />
                    <SPLIT distance="250" swimtime="00:04:10.43" />
                    <SPLIT distance="300" swimtime="00:05:03.16" />
                    <SPLIT distance="350" swimtime="00:05:55.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-28" firstname="Roman" gender="M" lastname="Pieślak" nation="POL" athleteid="7828">
              <RESULTS>
                <RESULT eventid="1195" points="360" reactiontime="+80" swimtime="00:00:29.37" resultid="7829" heatid="9325" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="1510" points="314" reactiontime="+81" swimtime="00:03:06.31" resultid="7830" heatid="9466" lane="3" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="364" swimtime="00:01:05.67" resultid="7831" heatid="9485" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="315" reactiontime="+70" swimtime="00:01:23.92" resultid="7832" heatid="9510" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="310" reactiontime="+73" swimtime="00:02:30.57" resultid="7833" heatid="9555" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:51.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="354" reactiontime="+60" swimtime="00:00:36.66" resultid="7834" heatid="9601" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="5636" points="278" reactiontime="+79" swimtime="00:05:36.87" resultid="7835" heatid="9615" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                    <SPLIT distance="200" swimtime="00:02:46.55" />
                    <SPLIT distance="250" swimtime="00:03:30.03" />
                    <SPLIT distance="300" swimtime="00:04:14.17" />
                    <SPLIT distance="350" swimtime="00:04:57.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="7840">
              <RESULTS>
                <RESULT eventid="1133" points="315" reactiontime="+86" swimtime="00:00:34.77" resultid="7841" heatid="9311" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1458" points="308" reactiontime="+71" swimtime="00:00:40.06" resultid="7842" heatid="9444" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1527" points="286" reactiontime="+78" swimtime="00:01:18.44" resultid="7843" heatid="9472" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="278" reactiontime="+74" swimtime="00:01:28.96" resultid="7844" heatid="9532" lane="9" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="239" reactiontime="+77" swimtime="00:03:19.70" resultid="7845" heatid="9581" lane="0" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                    <SPLIT distance="150" swimtime="00:02:30.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="7813">
              <RESULTS>
                <RESULT eventid="1229" points="309" reactiontime="+80" swimtime="00:02:48.60" resultid="7814" heatid="9346" lane="0" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="272" reactiontime="+93" swimtime="00:22:23.73" resultid="7815" heatid="9366" lane="5" entrytime="00:21:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:01.43" />
                    <SPLIT distance="200" swimtime="00:02:44.55" />
                    <SPLIT distance="250" swimtime="00:03:27.28" />
                    <SPLIT distance="300" swimtime="00:04:10.28" />
                    <SPLIT distance="350" swimtime="00:04:53.48" />
                    <SPLIT distance="400" swimtime="00:05:37.34" />
                    <SPLIT distance="450" swimtime="00:06:21.11" />
                    <SPLIT distance="500" swimtime="00:07:05.22" />
                    <SPLIT distance="550" swimtime="00:07:49.90" />
                    <SPLIT distance="600" swimtime="00:08:34.90" />
                    <SPLIT distance="650" swimtime="00:10:51.58" />
                    <SPLIT distance="700" swimtime="00:10:05.82" />
                    <SPLIT distance="750" swimtime="00:12:23.54" />
                    <SPLIT distance="800" swimtime="00:11:37.74" />
                    <SPLIT distance="850" swimtime="00:13:56.52" />
                    <SPLIT distance="900" swimtime="00:13:10.22" />
                    <SPLIT distance="950" swimtime="00:15:29.23" />
                    <SPLIT distance="1000" swimtime="00:14:43.15" />
                    <SPLIT distance="1050" swimtime="00:17:03.82" />
                    <SPLIT distance="1100" swimtime="00:16:15.67" />
                    <SPLIT distance="1150" swimtime="00:18:37.56" />
                    <SPLIT distance="1200" swimtime="00:17:50.85" />
                    <SPLIT distance="1250" swimtime="00:20:11.35" />
                    <SPLIT distance="1300" swimtime="00:19:24.94" />
                    <SPLIT distance="1350" swimtime="00:21:42.05" />
                    <SPLIT distance="1400" swimtime="00:20:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="368" reactiontime="+77" swimtime="00:00:33.54" resultid="7816" heatid="9454" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="5365" points="330" reactiontime="+73" swimtime="00:01:15.02" resultid="7817" heatid="9538" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="7818" heatid="9566" lane="5" entrytime="00:06:09.00" />
                <RESULT eventid="5551" points="280" reactiontime="+78" swimtime="00:02:50.95" resultid="7819" heatid="9588" lane="1" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:23.96" />
                    <SPLIT distance="150" swimtime="00:02:09.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="301" swimtime="00:05:28.19" resultid="7820" heatid="9615" lane="6" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:01:59.58" />
                    <SPLIT distance="200" swimtime="00:02:42.10" />
                    <SPLIT distance="250" swimtime="00:03:24.84" />
                    <SPLIT distance="300" swimtime="00:04:07.01" />
                    <SPLIT distance="350" swimtime="00:04:48.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-25" firstname="Tomasz" gender="M" lastname="Szymanowski" nation="POL" athleteid="7854">
              <RESULTS>
                <RESULT eventid="1195" points="385" reactiontime="+90" swimtime="00:00:28.73" resultid="7855" heatid="9325" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1280" points="272" reactiontime="+99" swimtime="00:11:37.39" resultid="7856" heatid="9361" lane="5" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:17.37" />
                    <SPLIT distance="150" swimtime="00:01:59.99" />
                    <SPLIT distance="200" swimtime="00:02:43.17" />
                    <SPLIT distance="250" swimtime="00:03:27.04" />
                    <SPLIT distance="300" swimtime="00:04:11.41" />
                    <SPLIT distance="350" swimtime="00:04:55.71" />
                    <SPLIT distance="400" swimtime="00:05:40.24" />
                    <SPLIT distance="450" swimtime="00:06:25.28" />
                    <SPLIT distance="500" swimtime="00:07:10.59" />
                    <SPLIT distance="550" swimtime="00:07:56.47" />
                    <SPLIT distance="600" swimtime="00:08:41.90" />
                    <SPLIT distance="650" swimtime="00:09:27.29" />
                    <SPLIT distance="700" swimtime="00:10:12.30" />
                    <SPLIT distance="750" swimtime="00:10:57.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="346" reactiontime="+89" swimtime="00:00:34.23" resultid="7857" heatid="9454" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="5365" points="311" reactiontime="+89" swimtime="00:01:16.50" resultid="7858" heatid="9538" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="280" reactiontime="+94" swimtime="00:02:50.97" resultid="7859" heatid="9588" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:08.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-14" firstname="Leszek" gender="M" lastname="Szwed" nation="POL" athleteid="7860">
              <RESULTS>
                <RESULT eventid="1195" points="83" reactiontime="+100" swimtime="00:00:47.79" resultid="7861" heatid="9318" lane="2" entrytime="00:00:47.68" />
                <RESULT eventid="1476" points="99" reactiontime="+101" swimtime="00:00:51.96" resultid="7862" heatid="9449" lane="7" entrytime="00:00:52.01" />
                <RESULT eventid="1544" points="83" swimtime="00:01:47.44" resultid="7863" heatid="9478" lane="9" entrytime="00:01:50.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="83" reactiontime="+91" swimtime="00:01:58.51" resultid="7864" heatid="9535" lane="2" entrytime="00:01:58.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="87" reactiontime="+92" swimtime="00:04:12.09" resultid="7865" heatid="9585" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.00" />
                    <SPLIT distance="100" swimtime="00:02:07.00" />
                    <SPLIT distance="150" swimtime="00:03:10.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-29" firstname="Lidia" gender="F" lastname="Mikołajczyk" nation="POL" athleteid="7799">
              <RESULTS>
                <RESULT eventid="1212" points="380" reactiontime="+90" swimtime="00:02:54.07" resultid="7800" heatid="9340" lane="0" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="150" swimtime="00:02:12.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="359" reactiontime="+98" swimtime="00:03:15.61" resultid="7801" heatid="9461" lane="8" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:32.88" />
                    <SPLIT distance="150" swimtime="00:02:24.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="413" reactiontime="+92" swimtime="00:01:09.39" resultid="7802" heatid="9474" lane="4" entrytime="00:01:10.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="358" reactiontime="+102" swimtime="00:01:30.31" resultid="7803" heatid="9504" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="337" swimtime="00:06:22.64" resultid="7804" heatid="9563" lane="6" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:28.84" />
                    <SPLIT distance="150" swimtime="00:02:20.25" />
                    <SPLIT distance="200" swimtime="00:03:09.76" />
                    <SPLIT distance="250" swimtime="00:04:03.65" />
                    <SPLIT distance="300" swimtime="00:04:54.54" />
                    <SPLIT distance="350" swimtime="00:05:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="364" reactiontime="+100" swimtime="00:00:41.15" resultid="7805" heatid="9595" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-28" firstname="Michał" gender="M" lastname="Pieślak" nation="POL" athleteid="7821">
              <RESULTS>
                <RESULT eventid="1195" points="382" reactiontime="+98" swimtime="00:00:28.80" resultid="7822" heatid="9326" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1544" points="379" swimtime="00:01:04.77" resultid="7823" heatid="9486" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" status="DNS" swimtime="00:00:00.00" resultid="7824" heatid="9509" lane="7" entrytime="00:01:28.00" />
                <RESULT eventid="5399" points="312" reactiontime="+91" swimtime="00:02:30.37" resultid="7825" heatid="9554" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:52.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="297" reactiontime="+86" swimtime="00:00:38.86" resultid="7826" heatid="9600" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="5636" points="316" reactiontime="+88" swimtime="00:05:23.00" resultid="7827" heatid="9615" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                    <SPLIT distance="200" swimtime="00:02:37.45" />
                    <SPLIT distance="250" swimtime="00:03:19.02" />
                    <SPLIT distance="300" swimtime="00:04:00.79" />
                    <SPLIT distance="350" swimtime="00:04:42.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="7806">
              <RESULTS>
                <RESULT eventid="1133" points="325" reactiontime="+88" swimtime="00:00:34.40" resultid="7807" heatid="9313" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1527" points="315" swimtime="00:01:15.97" resultid="7808" heatid="9474" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="206" reactiontime="+91" swimtime="00:01:48.45" resultid="7809" heatid="9502" lane="8" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="287" swimtime="00:02:51.24" resultid="7810" heatid="9546" lane="1" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="241" reactiontime="+96" swimtime="00:00:47.23" resultid="7811" heatid="9594" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="5619" points="246" reactiontime="+92" swimtime="00:06:17.03" resultid="7812" heatid="9610" lane="4" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:27.21" />
                    <SPLIT distance="150" swimtime="00:02:15.00" />
                    <SPLIT distance="200" swimtime="00:03:03.40" />
                    <SPLIT distance="250" swimtime="00:03:53.44" />
                    <SPLIT distance="300" swimtime="00:04:42.96" />
                    <SPLIT distance="350" swimtime="00:05:31.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1612" points="351" reactiontime="+80" swimtime="00:02:12.39" resultid="7869" heatid="9499" lane="9" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:10.50" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7813" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="7828" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="7836" number="3" />
                    <RELAYPOSITION athleteid="7821" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="5433" points="403" reactiontime="+79" swimtime="00:01:54.81" resultid="7871" heatid="9561" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:00:57.50" />
                    <SPLIT distance="150" swimtime="00:01:25.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7854" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="7828" number="2" reactiontime="+7" />
                    <RELAYPOSITION athleteid="7836" number="3" reactiontime="-12" />
                    <RELAYPOSITION athleteid="7821" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1595" points="293" reactiontime="+72" swimtime="00:02:39.75" resultid="7868" heatid="9497" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:31.68" />
                    <SPLIT distance="150" swimtime="00:02:06.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7840" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7846" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7799" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="7806" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="5416" points="327" reactiontime="+83" swimtime="00:02:20.17" resultid="7870" heatid="9559" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="150" swimtime="00:01:46.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7840" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="7846" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="7799" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="7806" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" swimtime="00:02:01.45" resultid="7866" heatid="9354" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:00:59.98" />
                    <SPLIT distance="150" swimtime="00:01:32.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7828" number="1" />
                    <RELAYPOSITION athleteid="7799" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="7806" number="3" />
                    <RELAYPOSITION athleteid="7854" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1246" reactiontime="+73" status="DSQ" swimtime="00:02:10.18" resultid="7867" heatid="9353" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="150" swimtime="00:01:41.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7840" number="1" reactiontime="+73" status="DSQ" />
                    <RELAYPOSITION athleteid="7836" number="2" reactiontime="-13" status="DSQ" />
                    <RELAYPOSITION athleteid="7846" number="3" reactiontime="+44" status="DSQ" />
                    <RELAYPOSITION athleteid="7821" number="4" reactiontime="+17" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+69" swimtime="00:02:19.73" resultid="7872" heatid="9607" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7840" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="7828" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="7799" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="7854" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+77" swimtime="00:02:59.71" resultid="7873" heatid="9607" lane="8" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                    <SPLIT distance="100" swimtime="00:01:50.81" />
                    <SPLIT distance="150" swimtime="00:02:24.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7860" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="7846" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="7813" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="7806" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="505815" nation="POL" region="WIE" clubid="6716" name="Tma Barracuda Kalisz">
          <CONTACT city="KALISZ" email="GALCZYNSKIWOJ@OP.PL" name="GAŁCZYŃSKI WOJCIECH" phone="790690666" state="WLKP" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1958-11-02" firstname="Anna" gender="F" lastname="Gałczyńska" nation="POL" athleteid="6724">
              <RESULTS>
                <RESULT eventid="1458" status="DNS" swimtime="00:00:00.00" resultid="6725" heatid="9440" lane="3" />
                <RESULT eventid="5279" status="DNS" swimtime="00:00:00.00" resultid="6726" heatid="9500" lane="3" entrytime="00:02:30.00" />
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="6727" heatid="9530" lane="8" entrytime="00:02:30.00" />
                <RESULT eventid="5568" status="DNS" swimtime="00:00:00.00" resultid="6728" heatid="9591" lane="4" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-12-13" firstname="Paweł" gender="M" lastname="Przybylski" nation="POL" athleteid="6754">
              <RESULTS>
                <RESULT eventid="1195" points="168" reactiontime="+118" swimtime="00:00:37.89" resultid="6755" heatid="9320" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1544" points="140" swimtime="00:01:30.17" resultid="6756" heatid="9478" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="95" reactiontime="+111" swimtime="00:03:43.29" resultid="6757" heatid="9549" lane="5" entrytime="00:03:49.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:42.16" />
                    <SPLIT distance="150" swimtime="00:02:41.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-13" firstname="Agata" gender="F" lastname="Gałczyńska" nation="POL" athleteid="6768">
              <RESULTS>
                <RESULT eventid="1458" points="87" reactiontime="+75" swimtime="00:01:00.84" resultid="6769" heatid="9441" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="5279" points="87" swimtime="00:02:24.59" resultid="6770" heatid="9501" lane="9" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="6771" heatid="9530" lane="7" entrytime="00:02:25.00" />
                <RESULT eventid="5568" points="89" swimtime="00:01:05.75" resultid="6772" heatid="9592" lane="1" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-11" firstname="Patrycja" gender="F" lastname="Rupa" nation="POL" athleteid="6717">
              <RESULTS>
                <RESULT eventid="1133" points="457" reactiontime="+76" swimtime="00:00:30.71" resultid="6718" heatid="9308" lane="5" />
                <RESULT eventid="1212" points="361" reactiontime="+84" swimtime="00:02:57.10" resultid="6719" heatid="9339" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:19.12" />
                    <SPLIT distance="150" swimtime="00:02:13.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="478" reactiontime="+59" swimtime="00:00:34.60" resultid="6720" heatid="9446" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="5314" status="DNS" swimtime="00:00:00.00" resultid="6721" heatid="9514" lane="9" />
                <RESULT eventid="5348" points="484" reactiontime="+61" swimtime="00:01:13.98" resultid="6722" heatid="9533" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="443" reactiontime="+57" swimtime="00:02:42.68" resultid="6723" heatid="9582" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:01.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-04" firstname="Elzbieta" gender="F" lastname="Tomczyk" nation="POL" athleteid="6748">
              <RESULTS>
                <RESULT eventid="1133" points="125" reactiontime="+107" swimtime="00:00:47.30" resultid="6749" heatid="9309" lane="6" entrytime="00:00:51.00" />
                <RESULT eventid="1527" points="119" swimtime="00:01:45.01" resultid="6751" heatid="9470" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="127" reactiontime="+89" swimtime="00:03:44.53" resultid="6752" heatid="9543" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:45.57" />
                    <SPLIT distance="150" swimtime="00:02:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="118" swimtime="00:08:01.62" resultid="6753" heatid="9612" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.54" />
                    <SPLIT distance="100" swimtime="00:01:52.58" />
                    <SPLIT distance="150" swimtime="00:02:53.12" />
                    <SPLIT distance="200" swimtime="00:03:55.11" />
                    <SPLIT distance="250" swimtime="00:04:58.55" />
                    <SPLIT distance="300" swimtime="00:06:00.91" />
                    <SPLIT distance="350" swimtime="00:07:02.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-30" firstname="Magdalena" gender="F" lastname="Kolera" nation="POL" athleteid="6759">
              <RESULTS>
                <RESULT eventid="1133" points="212" reactiontime="+115" swimtime="00:00:39.66" resultid="6760" heatid="9310" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1458" points="232" reactiontime="+70" swimtime="00:00:44.00" resultid="6762" heatid="9442" lane="2" entrytime="00:00:46.00" />
                <RESULT eventid="1527" points="183" reactiontime="+108" swimtime="00:01:30.98" resultid="6763" heatid="9471" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="193" reactiontime="+79" swimtime="00:01:40.39" resultid="6764" heatid="9531" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="6765" heatid="9543" lane="3" entrytime="00:03:30.00" />
                <RESULT eventid="5534" points="188" reactiontime="+85" swimtime="00:03:36.47" resultid="6766" heatid="9581" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.94" />
                    <SPLIT distance="100" swimtime="00:01:45.66" />
                    <SPLIT distance="150" swimtime="00:02:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="125" reactiontime="+116" swimtime="00:07:52.54" resultid="6767" heatid="9612" lane="0" entrytime="00:07:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:48.04" />
                    <SPLIT distance="150" swimtime="00:02:51.50" />
                    <SPLIT distance="200" swimtime="00:03:53.92" />
                    <SPLIT distance="250" swimtime="00:04:57.36" />
                    <SPLIT distance="300" swimtime="00:05:58.41" />
                    <SPLIT distance="350" swimtime="00:06:58.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-12" firstname="Wojciech" gender="M" lastname="Gałczyński" nation="POL" athleteid="6773">
              <RESULTS>
                <RESULT eventid="1195" points="461" reactiontime="+67" swimtime="00:00:27.05" resultid="6774" heatid="9330" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1476" points="360" reactiontime="+67" swimtime="00:00:33.78" resultid="6775" heatid="9447" lane="1" />
                <RESULT eventid="1510" points="321" reactiontime="+71" swimtime="00:03:04.91" resultid="6776" heatid="9466" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="309" reactiontime="+67" swimtime="00:01:24.45" resultid="6777" heatid="9511" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="331" reactiontime="+66" swimtime="00:01:14.90" resultid="6778" heatid="9539" lane="6" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="418" reactiontime="+76" swimtime="00:00:34.70" resultid="6779" heatid="9603" lane="8" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="6734">
              <RESULTS>
                <RESULT eventid="1195" points="257" reactiontime="+75" swimtime="00:00:32.86" resultid="6735" heatid="9322" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1229" points="217" swimtime="00:03:09.48" resultid="6736" heatid="9345" lane="9" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:02:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="230" reactiontime="+81" swimtime="00:03:26.51" resultid="6737" heatid="9464" lane="4" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:39.37" />
                    <SPLIT distance="150" swimtime="00:02:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="112" swimtime="00:03:50.76" resultid="6738" heatid="9494" lane="1" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                    <SPLIT distance="100" swimtime="00:01:42.83" />
                    <SPLIT distance="150" swimtime="00:02:45.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="213" swimtime="00:01:35.55" resultid="6739" heatid="9508" lane="6" entrytime="00:01:30.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="209" reactiontime="+76" swimtime="00:01:27.27" resultid="6740" heatid="9537" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="153" reactiontime="+76" swimtime="00:01:32.98" resultid="6741" heatid="9573" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="251" reactiontime="+61" swimtime="00:00:41.11" resultid="6742" heatid="9600" lane="1" entrytime="00:00:39.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-27" firstname="Małgorzata" gender="F" lastname="Rembowska-Świeboda" nation="POL" athleteid="6729">
              <RESULTS>
                <RESULT eventid="1133" points="383" reactiontime="+86" swimtime="00:00:32.57" resultid="6730" heatid="9312" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1458" points="383" reactiontime="+71" swimtime="00:00:37.23" resultid="6731" heatid="9444" lane="3" entrytime="00:00:39.40" />
                <RESULT eventid="1527" points="342" reactiontime="+86" swimtime="00:01:13.93" resultid="6732" heatid="9473" lane="7" entrytime="00:01:16.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="342" reactiontime="+76" swimtime="00:01:23.07" resultid="6733" heatid="9532" lane="1" entrytime="00:01:26.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-18" firstname="Marek" gender="M" lastname="Gola" nation="POL" athleteid="6743">
              <RESULTS>
                <RESULT eventid="1476" points="93" reactiontime="+124" swimtime="00:00:52.89" resultid="6744" heatid="9447" lane="7" />
                <RESULT eventid="1544" points="138" reactiontime="+106" swimtime="00:01:30.74" resultid="6745" heatid="9479" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="130" reactiontime="+93" swimtime="00:01:52.50" resultid="6746" heatid="9507" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="80" reactiontime="+99" swimtime="00:00:51.95" resultid="6747" heatid="9520" lane="9" entrytime="00:00:44.05" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="BARRACUDA MEN" number="1">
              <RESULTS>
                <RESULT eventid="5433" points="229" reactiontime="+100" swimtime="00:02:18.61" resultid="6782" heatid="9560" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="150" swimtime="00:01:50.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6754" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="6743" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="6734" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="6773" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="BARRACUDA MEN" number="2">
              <RESULTS>
                <RESULT eventid="1612" points="220" reactiontime="+60" swimtime="00:02:34.62" resultid="6781" heatid="9498" lane="6" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:01:57.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6773" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6743" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6734" number="3" />
                    <RELAYPOSITION athleteid="6754" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="BARRACUDA WOMEN" number="3">
              <RESULTS>
                <RESULT eventid="5416" points="167" swimtime="00:02:55.25" resultid="6780" heatid="9559" lane="1" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.60" />
                    <SPLIT distance="100" swimtime="00:01:38.95" />
                    <SPLIT distance="150" swimtime="00:02:23.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6768" number="1" />
                    <RELAYPOSITION athleteid="6759" number="2" />
                    <RELAYPOSITION athleteid="6748" number="3" />
                    <RELAYPOSITION athleteid="6729" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="BARRACUDA WOMEN" number="4">
              <RESULTS>
                <RESULT eventid="1595" points="173" reactiontime="+81" swimtime="00:03:10.24" resultid="6783" heatid="9497" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                    <SPLIT distance="100" swimtime="00:01:49.83" />
                    <SPLIT distance="150" swimtime="00:02:25.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6759" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="6768" number="2" />
                    <RELAYPOSITION athleteid="6729" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="6748" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="BARRACUDA MIX" number="5">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+85" swimtime="00:02:10.84" resultid="6784" heatid="9354" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                    <SPLIT distance="150" swimtime="00:01:44.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6759" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="6734" number="2" reactiontime="+4" />
                    <RELAYPOSITION athleteid="6729" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6773" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="BARRACUDA MIX" number="6">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+80" swimtime="00:02:27.88" resultid="6785" heatid="9607" lane="3" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:19.98" />
                    <SPLIT distance="150" swimtime="00:01:55.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6759" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6773" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="6734" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="6729" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03302" nation="POL" region="KUJ" clubid="8818" name="TMKS Champions Toruń">
          <CONTACT city="Toruń" email="slawekpredki@gmail.com" name="Prędki" phone="692449265" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1977-07-25" firstname="Sławomir" gender="M" lastname="Prędki" nation="POL" athleteid="8819">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1510" points="499" reactiontime="+79" swimtime="00:02:39.60" resultid="8820" heatid="9468" lane="0" entrytime="00:02:44.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="520" reactiontime="+77" swimtime="00:00:58.30" resultid="8821" heatid="9488" lane="0" entrytime="00:00:59.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="481" reactiontime="+76" swimtime="00:01:12.88" resultid="8822" heatid="9512" lane="3" entrytime="00:01:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="486" reactiontime="+77" swimtime="00:00:28.52" resultid="8823" heatid="9527" lane="1" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="8604" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="8631">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="8632" heatid="9318" lane="6" entrytime="00:00:46.21" />
                <RESULT eventid="1476" points="82" reactiontime="+82" swimtime="00:00:55.32" resultid="8633" heatid="9449" lane="1" entrytime="00:00:52.21" />
                <RESULT eventid="1510" points="94" reactiontime="+85" swimtime="00:04:37.88" resultid="8634" heatid="9463" lane="0" entrytime="00:04:27.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.57" />
                    <SPLIT distance="100" swimtime="00:02:10.22" />
                    <SPLIT distance="150" swimtime="00:03:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="97" reactiontime="+84" swimtime="00:02:04.09" resultid="8635" heatid="9506" lane="0" entrytime="00:02:02.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="8636" heatid="9535" lane="7" entrytime="00:02:05.31" />
                <RESULT eventid="5585" points="119" reactiontime="+119" swimtime="00:00:52.71" resultid="8637" heatid="9597" lane="4" entrytime="00:00:52.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-24" firstname="Anita" gender="F" lastname="Śliwa" nation="POL" athleteid="8665">
              <RESULTS>
                <RESULT eventid="1263" points="196" swimtime="00:13:53.58" resultid="8666" heatid="9356" lane="1" entrytime="00:13:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:32.90" />
                    <SPLIT distance="150" swimtime="00:02:24.74" />
                    <SPLIT distance="200" swimtime="00:03:17.51" />
                    <SPLIT distance="250" swimtime="00:04:10.48" />
                    <SPLIT distance="300" swimtime="00:05:04.16" />
                    <SPLIT distance="350" swimtime="00:05:58.02" />
                    <SPLIT distance="400" swimtime="00:06:51.54" />
                    <SPLIT distance="450" swimtime="00:07:44.86" />
                    <SPLIT distance="500" swimtime="00:08:37.97" />
                    <SPLIT distance="550" swimtime="00:09:31.16" />
                    <SPLIT distance="600" swimtime="00:10:25.38" />
                    <SPLIT distance="650" swimtime="00:11:17.50" />
                    <SPLIT distance="700" swimtime="00:12:10.72" />
                    <SPLIT distance="750" swimtime="00:13:03.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="221" reactiontime="+100" swimtime="00:00:44.72" resultid="8667" heatid="9443" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="5348" points="191" reactiontime="+86" swimtime="00:01:40.77" resultid="8668" heatid="9531" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="206" reactiontime="+91" swimtime="00:03:29.93" resultid="8669" heatid="9580" lane="5" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="150" swimtime="00:02:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="204" reactiontime="+96" swimtime="00:06:41.10" resultid="8670" heatid="9611" lane="2" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:23.96" />
                    <SPLIT distance="200" swimtime="00:03:15.51" />
                    <SPLIT distance="250" swimtime="00:04:07.13" />
                    <SPLIT distance="300" swimtime="00:04:59.78" />
                    <SPLIT distance="350" swimtime="00:05:52.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="8638">
              <RESULTS>
                <RESULT comment="Czas Lepszy od Rekordu Polski Kat A" eventid="1280" points="600" reactiontime="+76" swimtime="00:08:55.97" resultid="8639" heatid="9359" lane="4" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:36.68" />
                    <SPLIT distance="200" swimtime="00:02:10.76" />
                    <SPLIT distance="250" swimtime="00:02:44.90" />
                    <SPLIT distance="300" swimtime="00:03:18.82" />
                    <SPLIT distance="350" swimtime="00:03:52.76" />
                    <SPLIT distance="400" swimtime="00:04:26.77" />
                    <SPLIT distance="450" swimtime="00:05:00.65" />
                    <SPLIT distance="500" swimtime="00:05:34.66" />
                    <SPLIT distance="550" swimtime="00:06:08.77" />
                    <SPLIT distance="600" swimtime="00:06:43.00" />
                    <SPLIT distance="650" swimtime="00:07:16.95" />
                    <SPLIT distance="700" swimtime="00:07:51.38" />
                    <SPLIT distance="750" swimtime="00:08:24.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="624" reactiontime="+63" swimtime="00:02:28.23" resultid="8640" heatid="9468" lane="4" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="527" reactiontime="+71" swimtime="00:01:10.70" resultid="8641" heatid="9513" lane="0" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5467" points="587" swimtime="00:04:51.11" resultid="8642" heatid="9568" lane="6" entrytime="00:04:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                    <SPLIT distance="200" swimtime="00:02:28.67" />
                    <SPLIT distance="250" swimtime="00:03:08.22" />
                    <SPLIT distance="300" swimtime="00:03:47.41" />
                    <SPLIT distance="350" swimtime="00:04:20.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="563" reactiontime="+73" swimtime="00:00:31.42" resultid="8643" heatid="9604" lane="4" entrytime="00:00:31.90" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5636" points="629" reactiontime="+80" swimtime="00:04:16.78" resultid="8644" heatid="9613" lane="4" entrytime="00:04:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:33.30" />
                    <SPLIT distance="200" swimtime="00:02:06.19" />
                    <SPLIT distance="250" swimtime="00:02:39.24" />
                    <SPLIT distance="300" swimtime="00:03:12.33" />
                    <SPLIT distance="350" swimtime="00:03:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="8645">
              <RESULTS>
                <RESULT eventid="1195" points="259" reactiontime="+85" swimtime="00:00:32.80" resultid="8646" heatid="9323" lane="9" entrytime="00:00:31.30" />
                <RESULT eventid="1280" status="DNS" swimtime="00:00:00.00" resultid="8647" heatid="9360" lane="9" entrytime="00:11:45.00" />
                <RESULT eventid="1544" points="253" reactiontime="+87" swimtime="00:01:14.13" resultid="8648" heatid="9482" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="306" reactiontime="+87" swimtime="00:00:33.27" resultid="8649" heatid="9522" lane="1" entrytime="00:00:33.30" />
                <RESULT eventid="5399" points="236" reactiontime="+83" swimtime="00:02:44.90" resultid="8650" heatid="9552" lane="5" entrytime="00:02:47.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="208" reactiontime="+84" swimtime="00:01:24.03" resultid="8651" heatid="9575" lane="2" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="8671">
              <RESULTS>
                <RESULT eventid="1133" points="82" reactiontime="+130" swimtime="00:00:54.28" resultid="8672" heatid="9309" lane="7" entrytime="00:00:54.25" />
                <RESULT eventid="1458" points="76" reactiontime="+99" swimtime="00:01:03.79" resultid="8673" heatid="9441" lane="0" entrytime="00:01:03.39" />
                <RESULT eventid="1527" points="77" reactiontime="+126" swimtime="00:02:01.20" resultid="8674" heatid="9470" lane="0" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="79" reactiontime="+103" swimtime="00:02:15.09" resultid="8675" heatid="9530" lane="2" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="71" reactiontime="+90" swimtime="00:04:58.51" resultid="8676" heatid="9579" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.99" />
                    <SPLIT distance="100" swimtime="00:02:25.72" />
                    <SPLIT distance="150" swimtime="00:03:45.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="8658">
              <RESULTS>
                <RESULT eventid="1280" points="404" reactiontime="+62" swimtime="00:10:11.33" resultid="8659" heatid="9359" lane="7" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:44.31" />
                    <SPLIT distance="200" swimtime="00:02:21.66" />
                    <SPLIT distance="250" swimtime="00:02:59.49" />
                    <SPLIT distance="300" swimtime="00:03:37.61" />
                    <SPLIT distance="350" swimtime="00:04:16.25" />
                    <SPLIT distance="400" swimtime="00:04:55.46" />
                    <SPLIT distance="450" swimtime="00:05:34.90" />
                    <SPLIT distance="500" swimtime="00:06:15.00" />
                    <SPLIT distance="550" swimtime="00:06:54.83" />
                    <SPLIT distance="600" swimtime="00:07:34.77" />
                    <SPLIT distance="650" swimtime="00:08:14.75" />
                    <SPLIT distance="700" swimtime="00:08:54.15" />
                    <SPLIT distance="750" swimtime="00:09:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="459" reactiontime="+73" swimtime="00:02:44.10" resultid="8660" heatid="9468" lane="8" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="522" swimtime="00:01:10.93" resultid="8661" heatid="9513" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="471" reactiontime="+78" swimtime="00:02:11.03" resultid="8662" heatid="9557" lane="5" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="532" reactiontime="+80" swimtime="00:00:32.02" resultid="8663" heatid="9604" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="5636" points="455" swimtime="00:04:46.09" resultid="8664" heatid="9613" lane="9" entrytime="00:04:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:43.32" />
                    <SPLIT distance="200" swimtime="00:02:20.27" />
                    <SPLIT distance="250" swimtime="00:02:57.13" />
                    <SPLIT distance="300" swimtime="00:03:34.56" />
                    <SPLIT distance="350" swimtime="00:04:11.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="8627">
              <RESULTS>
                <RESULT eventid="1195" points="21" reactiontime="+131" swimtime="00:01:14.76" resultid="8628" heatid="9317" lane="4" entrytime="00:01:05.40" />
                <RESULT eventid="1476" points="18" reactiontime="+114" swimtime="00:01:30.44" resultid="8629" heatid="9447" lane="5" entrytime="00:01:58.45" />
                <RESULT eventid="5585" points="13" reactiontime="+130" swimtime="00:01:48.18" resultid="8630" heatid="9597" lane="8" entrytime="00:01:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="8677">
              <RESULTS>
                <RESULT eventid="1133" points="481" reactiontime="+84" swimtime="00:00:30.19" resultid="8678" heatid="9314" lane="6" entrytime="00:00:29.99" />
                <RESULT eventid="1212" points="455" swimtime="00:02:43.93" resultid="8679" heatid="9340" lane="6" entrytime="00:02:39.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:05.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="412" reactiontime="+74" swimtime="00:03:06.90" resultid="8680" heatid="9460" lane="4" entrytime="00:03:13.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:02:17.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="441" swimtime="00:01:07.91" resultid="8681" heatid="9475" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="386" swimtime="00:01:28.02" resultid="8682" heatid="9504" lane="1" entrytime="00:01:25.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="426" reactiontime="+73" swimtime="00:02:30.05" resultid="8683" heatid="9546" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:01:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="406" reactiontime="+78" swimtime="00:00:39.70" resultid="8684" heatid="9595" lane="3" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-11" firstname="Kamil" gender="M" lastname="Kordowski" nation="POL" athleteid="8653">
              <RESULTS>
                <RESULT eventid="1195" points="416" reactiontime="+82" swimtime="00:00:28.01" resultid="8654" heatid="9327" lane="7" entrytime="00:00:28.14" />
                <RESULT eventid="1544" points="419" reactiontime="+75" swimtime="00:01:02.67" resultid="8655" heatid="9485" lane="4" entrytime="00:01:03.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="356" reactiontime="+93" swimtime="00:00:31.63" resultid="8656" heatid="9523" lane="9" entrytime="00:00:32.29" />
                <RESULT eventid="5517" points="270" swimtime="00:01:17.02" resultid="8657" heatid="9575" lane="6" entrytime="00:01:17.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-04" firstname="Andrzej" gender="M" lastname="Marchewka" nation="POL" athleteid="8694">
              <RESULTS>
                <RESULT eventid="1476" points="394" reactiontime="+71" swimtime="00:00:32.77" resultid="8695" heatid="9456" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="5365" points="335" reactiontime="+79" swimtime="00:01:14.59" resultid="8696" heatid="9540" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="273" reactiontime="+74" swimtime="00:02:52.36" resultid="8697" heatid="9588" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:10.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="8611">
              <RESULTS>
                <RESULT eventid="1195" points="88" reactiontime="+116" swimtime="00:00:46.92" resultid="8612" heatid="9319" lane="2" entrytime="00:00:40.72" />
                <RESULT eventid="1229" points="47" reactiontime="+120" swimtime="00:05:15.10" resultid="8613" heatid="9342" lane="5" entrytime="00:05:07.26">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:49.21" />
                    <SPLIT distance="150" swimtime="00:04:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="32" reactiontime="+103" swimtime="00:01:15.03" resultid="8614" heatid="9447" lane="4" entrytime="00:01:10.41" />
                <RESULT eventid="1578" points="29" reactiontime="+117" swimtime="00:06:02.47" resultid="8615" heatid="9493" lane="0" entrytime="00:05:30.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.99" />
                    <SPLIT distance="100" swimtime="00:03:00.23" />
                    <SPLIT distance="150" swimtime="00:04:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="55" reactiontime="+130" swimtime="00:04:27.81" resultid="8616" heatid="9549" lane="7" entrytime="00:04:03.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:02:13.15" />
                    <SPLIT distance="150" swimtime="00:03:27.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="46" reactiontime="+115" swimtime="00:11:20.21" resultid="8617" heatid="9564" lane="2" entrytime="00:10:59.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.70" />
                    <SPLIT distance="100" swimtime="00:02:48.13" />
                    <SPLIT distance="150" swimtime="00:04:24.08" />
                    <SPLIT distance="200" swimtime="00:05:57.88" />
                    <SPLIT distance="250" swimtime="00:07:33.93" />
                    <SPLIT distance="300" swimtime="00:09:05.72" />
                    <SPLIT distance="350" swimtime="00:10:15.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="29" reactiontime="+114" swimtime="00:02:41.52" resultid="8618" heatid="9572" lane="7" entrytime="00:02:35.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="8686">
              <RESULTS>
                <RESULT eventid="1195" points="260" reactiontime="+89" swimtime="00:00:32.72" resultid="8687" heatid="9322" lane="8" entrytime="00:00:32.80" />
                <RESULT eventid="1280" points="179" swimtime="00:13:21.31" resultid="8688" heatid="9361" lane="7" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:33.95" />
                    <SPLIT distance="150" swimtime="00:02:24.41" />
                    <SPLIT distance="200" swimtime="00:03:15.57" />
                    <SPLIT distance="250" swimtime="00:04:06.94" />
                    <SPLIT distance="300" swimtime="00:04:58.31" />
                    <SPLIT distance="350" swimtime="00:05:49.48" />
                    <SPLIT distance="400" swimtime="00:06:40.53" />
                    <SPLIT distance="450" swimtime="00:07:32.49" />
                    <SPLIT distance="500" swimtime="00:08:24.08" />
                    <SPLIT distance="550" swimtime="00:09:15.44" />
                    <SPLIT distance="600" swimtime="00:10:07.17" />
                    <SPLIT distance="650" swimtime="00:10:57.36" />
                    <SPLIT distance="700" swimtime="00:11:47.85" />
                    <SPLIT distance="750" swimtime="00:12:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="239" reactiontime="+84" swimtime="00:01:15.54" resultid="8689" heatid="9481" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="221" reactiontime="+79" swimtime="00:00:37.05" resultid="8690" heatid="9521" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="5399" points="191" reactiontime="+88" swimtime="00:02:56.91" resultid="8691" heatid="9552" lane="0" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:28.38" />
                    <SPLIT distance="150" swimtime="00:02:14.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="162" swimtime="00:01:31.22" resultid="8692" heatid="9573" lane="6" entrytime="00:01:35.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="188" reactiontime="+78" swimtime="00:06:23.69" resultid="8693" heatid="9617" lane="7" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                    <SPLIT distance="200" swimtime="00:03:10.44" />
                    <SPLIT distance="250" swimtime="00:03:59.96" />
                    <SPLIT distance="300" swimtime="00:04:49.06" />
                    <SPLIT distance="350" swimtime="00:05:38.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="8620">
              <RESULTS>
                <RESULT eventid="1195" points="118" reactiontime="+119" swimtime="00:00:42.62" resultid="8621" heatid="9319" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1476" points="50" reactiontime="+86" swimtime="00:01:04.95" resultid="8622" heatid="9448" lane="0" entrytime="00:01:05.25" />
                <RESULT eventid="1544" points="89" reactiontime="+97" swimtime="00:01:44.85" resultid="8623" heatid="9478" lane="7" entrytime="00:01:43.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="41" reactiontime="+72" swimtime="00:02:29.54" resultid="8624" heatid="9535" lane="8" entrytime="00:02:12.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="66" reactiontime="+112" swimtime="00:04:12.24" resultid="8625" heatid="9549" lane="4" entrytime="00:03:48.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.27" />
                    <SPLIT distance="100" swimtime="00:02:01.52" />
                    <SPLIT distance="150" swimtime="00:03:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="45" reactiontime="+87" swimtime="00:05:13.73" resultid="8626" heatid="9584" lane="1" entrytime="00:04:48.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.98" />
                    <SPLIT distance="100" swimtime="00:02:35.08" />
                    <SPLIT distance="150" swimtime="00:03:56.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1612" points="458" reactiontime="+73" swimtime="00:02:01.14" resultid="8700" heatid="9499" lane="2" entrytime="00:02:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:02.88" />
                    <SPLIT distance="150" swimtime="00:01:35.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8694" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="8638" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="8645" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="8658" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5433" points="459" reactiontime="+86" swimtime="00:01:49.99" resultid="8701" heatid="9561" lane="7" entrytime="00:01:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="100" swimtime="00:00:57.10" />
                    <SPLIT distance="150" swimtime="00:01:23.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8658" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="8645" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="8694" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="8638" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1612" points="83" reactiontime="+88" swimtime="00:03:34.04" resultid="8702" heatid="9498" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.10" />
                    <SPLIT distance="100" swimtime="00:02:08.39" />
                    <SPLIT distance="150" swimtime="00:02:50.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8611" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="8631" number="2" reactiontime="+96" />
                    <RELAYPOSITION athleteid="8686" number="3" />
                    <RELAYPOSITION athleteid="8620" number="4" reactiontime="+92" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5433" points="115" reactiontime="+74" swimtime="00:02:54.13" resultid="8703" heatid="9560" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:02:06.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8686" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="8620" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="8631" number="3" />
                    <RELAYPOSITION athleteid="8611" number="4" reactiontime="+101" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+93" swimtime="00:02:38.19" resultid="8698" heatid="9353" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:07.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8686" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="8671" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="8665" number="3" />
                    <RELAYPOSITION athleteid="8645" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5602" reactiontime="+85" swimtime="00:02:57.31" resultid="8699" heatid="9606" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8665" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="8671" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="8645" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="8686" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="8244" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="8253">
              <RESULTS>
                <RESULT eventid="1280" points="119" reactiontime="+104" swimtime="00:15:16.80" resultid="8254" heatid="9362" lane="8" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.00" />
                    <SPLIT distance="100" swimtime="00:01:48.91" />
                    <SPLIT distance="150" swimtime="00:02:46.38" />
                    <SPLIT distance="200" swimtime="00:03:44.74" />
                    <SPLIT distance="250" swimtime="00:04:42.93" />
                    <SPLIT distance="300" swimtime="00:05:41.99" />
                    <SPLIT distance="350" swimtime="00:06:39.35" />
                    <SPLIT distance="400" swimtime="00:07:40.09" />
                    <SPLIT distance="450" swimtime="00:08:37.00" />
                    <SPLIT distance="500" swimtime="00:09:35.18" />
                    <SPLIT distance="550" swimtime="00:10:33.13" />
                    <SPLIT distance="600" swimtime="00:11:30.66" />
                    <SPLIT distance="650" swimtime="00:12:27.55" />
                    <SPLIT distance="700" swimtime="00:13:26.25" />
                    <SPLIT distance="750" swimtime="00:14:23.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="157" reactiontime="+87" swimtime="00:00:44.47" resultid="8255" heatid="9450" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="5365" points="116" reactiontime="+85" swimtime="00:01:46.31" resultid="8256" heatid="9536" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="8257" heatid="9585" lane="7" entrytime="00:03:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-01" firstname="Lech" gender="M" lastname="Sarnowski" nation="POL" athleteid="8245">
              <RESULTS>
                <RESULT eventid="1195" points="68" swimtime="00:00:51.04" resultid="8246" heatid="9318" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1476" points="39" reactiontime="+74" swimtime="00:01:10.45" resultid="8247" heatid="9448" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="5585" points="89" reactiontime="+104" swimtime="00:00:58.10" resultid="8248" heatid="9597" lane="6" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Agnieszka" gender="F" lastname="Rybak-Starczak" nation="POL" athleteid="8290">
              <RESULTS>
                <RESULT eventid="1212" points="274" reactiontime="+117" swimtime="00:03:14.14" resultid="8291" heatid="9338" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:33.04" />
                    <SPLIT distance="150" swimtime="00:02:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="280" swimtime="00:03:32.55" resultid="8292" heatid="9460" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:42.75" />
                    <SPLIT distance="150" swimtime="00:02:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="295" reactiontime="+104" swimtime="00:01:36.27" resultid="8293" heatid="9503" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="8249">
              <RESULTS>
                <RESULT eventid="1476" points="137" reactiontime="+79" swimtime="00:00:46.61" resultid="8250" heatid="9450" lane="9" entrytime="00:00:46.00" />
                <RESULT eventid="5365" points="119" reactiontime="+78" swimtime="00:01:45.35" resultid="8251" heatid="9536" lane="9" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="108" reactiontime="+76" swimtime="00:03:54.41" resultid="8252" heatid="9585" lane="2" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.63" />
                    <SPLIT distance="100" swimtime="00:01:53.82" />
                    <SPLIT distance="150" swimtime="00:02:55.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Wojciech" gender="M" lastname="Niewitecki" nation="POL" athleteid="8266">
              <RESULTS>
                <RESULT eventid="1476" points="205" reactiontime="+93" swimtime="00:00:40.77" resultid="8267" heatid="9452" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="5365" points="173" reactiontime="+81" swimtime="00:01:32.99" resultid="8268" heatid="9536" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="8269">
              <RESULTS>
                <RESULT eventid="1510" points="302" reactiontime="+81" swimtime="00:03:08.68" resultid="8270" heatid="9465" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:29.23" />
                    <SPLIT distance="150" swimtime="00:02:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="325" reactiontime="+81" swimtime="00:01:23.05" resultid="8271" heatid="9509" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="322" reactiontime="+81" swimtime="00:00:37.83" resultid="8272" heatid="9601" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="8282">
              <RESULTS>
                <RESULT eventid="1133" points="191" reactiontime="+90" swimtime="00:00:41.05" resultid="8283" heatid="9310" lane="2" entrytime="00:00:41.00" />
                <RESULT comment="Czas Lepszy od Rekordu Polski Kat. I" eventid="1297" points="149" swimtime="00:29:04.19" resultid="8284" heatid="9364" lane="7" entrytime="00:34:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:47.16" />
                    <SPLIT distance="150" swimtime="00:02:45.05" />
                    <SPLIT distance="200" swimtime="00:03:43.39" />
                    <SPLIT distance="250" swimtime="00:04:41.41" />
                    <SPLIT distance="300" swimtime="00:05:38.81" />
                    <SPLIT distance="350" swimtime="00:06:37.17" />
                    <SPLIT distance="400" swimtime="00:07:36.06" />
                    <SPLIT distance="450" swimtime="00:08:35.54" />
                    <SPLIT distance="500" swimtime="00:09:34.18" />
                    <SPLIT distance="550" swimtime="00:10:33.28" />
                    <SPLIT distance="600" swimtime="00:11:31.94" />
                    <SPLIT distance="650" swimtime="00:12:32.10" />
                    <SPLIT distance="700" swimtime="00:13:31.90" />
                    <SPLIT distance="750" swimtime="00:14:31.35" />
                    <SPLIT distance="800" swimtime="00:15:30.35" />
                    <SPLIT distance="850" swimtime="00:16:29.74" />
                    <SPLIT distance="900" swimtime="00:17:29.18" />
                    <SPLIT distance="950" swimtime="00:18:28.42" />
                    <SPLIT distance="1000" swimtime="00:19:27.36" />
                    <SPLIT distance="1050" swimtime="00:20:26.96" />
                    <SPLIT distance="1100" swimtime="00:21:25.40" />
                    <SPLIT distance="1150" swimtime="00:22:24.60" />
                    <SPLIT distance="1200" swimtime="00:23:23.02" />
                    <SPLIT distance="1250" swimtime="00:24:22.71" />
                    <SPLIT distance="1300" swimtime="00:25:20.65" />
                    <SPLIT distance="1350" swimtime="00:26:19.31" />
                    <SPLIT distance="1400" swimtime="00:27:16.87" />
                    <SPLIT distance="1450" swimtime="00:28:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="139" reactiontime="+85" swimtime="00:00:52.12" resultid="8285" heatid="9442" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="5314" points="111" reactiontime="+93" swimtime="00:00:50.76" resultid="8286" heatid="9514" lane="2" entrytime="00:00:53.00" />
                <RESULT eventid="5382" points="166" swimtime="00:03:25.30" resultid="8287" heatid="9543" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:41.31" />
                    <SPLIT distance="150" swimtime="00:02:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="135" reactiontime="+74" swimtime="00:04:01.69" resultid="8288" heatid="9580" lane="0" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.45" />
                    <SPLIT distance="100" swimtime="00:01:58.73" />
                    <SPLIT distance="150" swimtime="00:03:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="148" swimtime="00:07:26.83" resultid="8289" heatid="9611" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:47.61" />
                    <SPLIT distance="150" swimtime="00:02:46.32" />
                    <SPLIT distance="200" swimtime="00:03:44.43" />
                    <SPLIT distance="250" swimtime="00:04:41.51" />
                    <SPLIT distance="300" swimtime="00:05:37.02" />
                    <SPLIT distance="350" swimtime="00:06:33.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="8259">
              <RESULTS>
                <RESULT eventid="1229" points="198" reactiontime="+89" swimtime="00:03:15.58" resultid="8260" heatid="9344" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="150" swimtime="00:02:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="186" swimtime="00:13:11.33" resultid="8261" heatid="9361" lane="6" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                    <SPLIT distance="200" swimtime="00:03:14.32" />
                    <SPLIT distance="250" swimtime="00:04:04.89" />
                    <SPLIT distance="300" swimtime="00:04:56.14" />
                    <SPLIT distance="350" swimtime="00:05:47.01" />
                    <SPLIT distance="400" swimtime="00:06:37.35" />
                    <SPLIT distance="450" swimtime="00:07:27.23" />
                    <SPLIT distance="500" swimtime="00:08:16.90" />
                    <SPLIT distance="550" swimtime="00:09:06.48" />
                    <SPLIT distance="600" swimtime="00:09:55.82" />
                    <SPLIT distance="650" swimtime="00:10:45.24" />
                    <SPLIT distance="700" swimtime="00:11:34.75" />
                    <SPLIT distance="750" swimtime="00:12:23.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="182" reactiontime="+82" swimtime="00:00:42.38" resultid="8262" heatid="9451" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="5365" points="175" reactiontime="+91" swimtime="00:01:32.69" resultid="8263" heatid="9537" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="201" swimtime="00:06:55.83" resultid="8264" heatid="9566" lane="9" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.20" />
                    <SPLIT distance="100" swimtime="00:01:50.05" />
                    <SPLIT distance="150" swimtime="00:02:41.77" />
                    <SPLIT distance="200" swimtime="00:03:32.25" />
                    <SPLIT distance="250" swimtime="00:04:28.38" />
                    <SPLIT distance="300" swimtime="00:05:24.86" />
                    <SPLIT distance="350" swimtime="00:06:10.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="185" reactiontime="+80" swimtime="00:03:16.13" resultid="8265" heatid="9586" lane="6" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:36.98" />
                    <SPLIT distance="150" swimtime="00:02:27.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Jacek" gender="M" lastname="Matyszczak" nation="POL" athleteid="8273">
              <RESULTS>
                <RESULT eventid="1195" points="389" reactiontime="+86" swimtime="00:00:28.64" resultid="8274" heatid="9327" lane="0" entrytime="00:00:28.50" />
                <RESULT eventid="1229" points="270" reactiontime="+91" swimtime="00:02:56.31" resultid="8275" heatid="9345" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="233" reactiontime="+87" swimtime="00:00:39.03" resultid="8276" heatid="9452" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1544" points="355" reactiontime="+88" swimtime="00:01:06.19" resultid="8277" heatid="9484" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="314" reactiontime="+103" swimtime="00:00:32.99" resultid="8278" heatid="9523" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="5399" points="291" swimtime="00:02:33.83" resultid="8279" heatid="9553" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="190" reactiontime="+80" swimtime="00:03:14.44" resultid="8280" heatid="9587" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:34.55" />
                    <SPLIT distance="150" swimtime="00:02:25.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="268" reactiontime="+100" swimtime="00:05:41.12" resultid="8281" heatid="9616" lane="7" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                    <SPLIT distance="200" swimtime="00:02:43.26" />
                    <SPLIT distance="250" swimtime="00:03:27.40" />
                    <SPLIT distance="300" swimtime="00:04:12.07" />
                    <SPLIT distance="350" swimtime="00:04:58.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="210" reactiontime="+79" swimtime="00:02:37.16" resultid="8294" heatid="9498" lane="2" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:23.32" />
                    <SPLIT distance="150" swimtime="00:01:59.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8266" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="8259" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="8269" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="8253" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="100413" nation="POL" region="WAR" clubid="6630" name="UKP Jedynka Elbląg">
          <CONTACT name="Wysocki" phone="696427414" />
          <ATHLETES>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="6631">
              <RESULTS>
                <RESULT eventid="1212" points="104" reactiontime="+122" swimtime="00:04:27.47" resultid="6632" heatid="9337" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                    <SPLIT distance="100" swimtime="00:02:09.61" />
                    <SPLIT distance="150" swimtime="00:03:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="152" reactiontime="+111" swimtime="00:28:53.21" resultid="6633" heatid="9364" lane="2" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:48.79" />
                    <SPLIT distance="150" swimtime="00:02:45.99" />
                    <SPLIT distance="200" swimtime="00:03:44.62" />
                    <SPLIT distance="250" swimtime="00:04:43.63" />
                    <SPLIT distance="300" swimtime="00:05:42.56" />
                    <SPLIT distance="350" swimtime="00:06:41.01" />
                    <SPLIT distance="400" swimtime="00:07:39.28" />
                    <SPLIT distance="450" swimtime="00:08:37.85" />
                    <SPLIT distance="500" swimtime="00:09:35.59" />
                    <SPLIT distance="550" swimtime="00:10:33.47" />
                    <SPLIT distance="600" swimtime="00:11:33.14" />
                    <SPLIT distance="650" swimtime="00:12:30.98" />
                    <SPLIT distance="700" swimtime="00:13:30.09" />
                    <SPLIT distance="750" swimtime="00:14:27.90" />
                    <SPLIT distance="800" swimtime="00:15:25.47" />
                    <SPLIT distance="850" swimtime="00:16:23.13" />
                    <SPLIT distance="900" swimtime="00:17:20.96" />
                    <SPLIT distance="950" swimtime="00:18:18.78" />
                    <SPLIT distance="1000" swimtime="00:19:17.03" />
                    <SPLIT distance="1050" swimtime="00:20:14.64" />
                    <SPLIT distance="1100" swimtime="00:21:12.72" />
                    <SPLIT distance="1150" swimtime="00:22:10.32" />
                    <SPLIT distance="1200" swimtime="00:23:08.22" />
                    <SPLIT distance="1250" swimtime="00:24:05.90" />
                    <SPLIT distance="1300" swimtime="00:25:04.17" />
                    <SPLIT distance="1350" swimtime="00:26:02.01" />
                    <SPLIT distance="1400" swimtime="00:27:00.25" />
                    <SPLIT distance="1450" swimtime="00:27:57.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="114" reactiontime="+106" swimtime="00:01:46.63" resultid="6634" heatid="9471" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="99" swimtime="00:04:22.55" resultid="6635" heatid="9491" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.06" />
                    <SPLIT distance="100" swimtime="00:02:04.88" />
                    <SPLIT distance="150" swimtime="00:03:15.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" status="DNS" swimtime="00:00:00.00" resultid="6636" heatid="9543" lane="2" entrytime="00:03:35.00" />
                <RESULT eventid="5450" points="105" reactiontime="+117" swimtime="00:09:24.11" resultid="6637" heatid="9562" lane="8" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                    <SPLIT distance="100" swimtime="00:02:08.19" />
                    <SPLIT distance="150" swimtime="00:03:21.31" />
                    <SPLIT distance="200" swimtime="00:04:36.11" />
                    <SPLIT distance="250" swimtime="00:06:00.48" />
                    <SPLIT distance="300" swimtime="00:07:25.19" />
                    <SPLIT distance="350" swimtime="00:08:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" status="DNS" swimtime="00:00:00.00" resultid="6638" heatid="9611" lane="9" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:39.40" />
                    <SPLIT distance="150" swimtime="00:02:33.39" />
                    <SPLIT distance="200" swimtime="00:03:28.15" />
                    <SPLIT distance="250" swimtime="00:04:23.44" />
                    <SPLIT distance="300" swimtime="00:05:19.19" />
                    <SPLIT distance="350" swimtime="00:06:14.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="6639">
              <RESULTS>
                <RESULT eventid="1133" points="146" reactiontime="+101" swimtime="00:00:44.91" resultid="6640" heatid="9310" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1263" reactiontime="+94" status="OTL" swimtime="00:00:00.00" resultid="6641" heatid="9356" lane="2" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                    <SPLIT distance="100" swimtime="00:01:49.02" />
                    <SPLIT distance="150" swimtime="00:02:48.39" />
                    <SPLIT distance="200" swimtime="00:03:48.26" />
                    <SPLIT distance="250" swimtime="00:04:48.58" />
                    <SPLIT distance="300" swimtime="00:05:47.99" />
                    <SPLIT distance="350" swimtime="00:06:47.21" />
                    <SPLIT distance="400" swimtime="00:07:46.78" />
                    <SPLIT distance="450" swimtime="00:08:46.44" />
                    <SPLIT distance="500" swimtime="00:09:45.71" />
                    <SPLIT distance="550" swimtime="00:10:45.10" />
                    <SPLIT distance="600" swimtime="00:11:43.30" />
                    <SPLIT distance="650" swimtime="00:12:41.75" />
                    <SPLIT distance="700" swimtime="00:13:39.96" />
                    <SPLIT distance="750" swimtime="00:14:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="144" reactiontime="+98" swimtime="00:01:38.50" resultid="6642" heatid="9470" lane="4" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="156" swimtime="00:03:29.57" resultid="6643" heatid="9543" lane="6" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="153" reactiontime="+100" swimtime="00:07:21.86" resultid="6644" heatid="9611" lane="8" entrytime="00:07:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                    <SPLIT distance="100" swimtime="00:01:46.22" />
                    <SPLIT distance="150" swimtime="00:02:43.65" />
                    <SPLIT distance="200" swimtime="00:03:41.26" />
                    <SPLIT distance="250" swimtime="00:04:36.96" />
                    <SPLIT distance="300" swimtime="00:05:34.29" />
                    <SPLIT distance="350" swimtime="00:06:29.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="6645">
              <RESULTS>
                <RESULT comment="Z3 - Pływak ukończył poszczególne odcinki niezgodnie z przepisami o zakończeniu wyścigu w danym stylu., /K14" eventid="1229" reactiontime="+72" status="DSQ" swimtime="00:02:35.33" resultid="6646" heatid="9347" lane="2" entrytime="00:02:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="444" reactiontime="+75" swimtime="00:02:13.64" resultid="6647" heatid="9556" lane="4" entrytime="00:02:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                    <SPLIT distance="150" swimtime="00:01:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6648" heatid="9576" lane="4" entrytime="00:01:08.00" />
                <RESULT eventid="5636" points="434" reactiontime="+80" swimtime="00:04:50.51" resultid="6649" heatid="9614" lane="3" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                    <SPLIT distance="200" swimtime="00:02:21.59" />
                    <SPLIT distance="250" swimtime="00:02:58.64" />
                    <SPLIT distance="300" swimtime="00:03:36.46" />
                    <SPLIT distance="350" swimtime="00:04:14.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="7073">
              <RESULTS>
                <RESULT eventid="1263" status="OTL" swimtime="00:20:59.40" resultid="7074" heatid="9357" lane="6" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.72" />
                    <SPLIT distance="100" swimtime="00:02:29.69" />
                    <SPLIT distance="150" swimtime="00:03:49.51" />
                    <SPLIT distance="200" swimtime="00:05:07.60" />
                    <SPLIT distance="250" swimtime="00:09:05.50" />
                    <SPLIT distance="300" swimtime="00:07:46.46" />
                    <SPLIT distance="350" swimtime="00:11:43.68" />
                    <SPLIT distance="400" swimtime="00:10:24.37" />
                    <SPLIT distance="450" swimtime="00:14:22.61" />
                    <SPLIT distance="500" swimtime="00:13:02.93" />
                    <SPLIT distance="550" swimtime="00:17:03.56" />
                    <SPLIT distance="600" swimtime="00:15:42.97" />
                    <SPLIT distance="650" swimtime="00:19:43.05" />
                    <SPLIT distance="700" swimtime="00:18:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="59" reactiontime="+88" swimtime="00:01:09.35" resultid="7075" heatid="9440" lane="4" entrytime="00:01:07.00" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1493" status="DSQ" swimtime="00:06:18.87" resultid="7076" heatid="9458" lane="7" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.51" />
                    <SPLIT distance="100" swimtime="00:03:11.68" />
                    <SPLIT distance="150" swimtime="00:04:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="5279" status="DSQ" swimtime="00:03:12.77" resultid="7077" heatid="9500" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="46" reactiontime="+167" swimtime="00:02:41.48" resultid="7078" heatid="9529" lane="4" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="48" reactiontime="+87" swimtime="00:05:39.35" resultid="7079" heatid="9579" lane="6" entrytime="00:05:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.90" />
                    <SPLIT distance="100" swimtime="00:02:48.97" />
                    <SPLIT distance="150" swimtime="00:04:16.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08314" nation="POL" region="MAZ" clubid="6852" name="UKS Delfin Garwolin">
          <CONTACT name="Mianowski" />
          <ATHLETES>
            <ATHLETE birthdate="1996-12-29" firstname="Mateusz" gender="M" lastname="Szczypek" nation="POL" athleteid="6853">
              <RESULTS>
                <RESULT eventid="1195" points="428" reactiontime="+81" swimtime="00:00:27.73" resultid="6854" heatid="9328" lane="7" entrytime="00:00:27.47" />
                <RESULT eventid="1280" points="372" reactiontime="+55" swimtime="00:10:28.24" resultid="6855" heatid="9360" lane="7" entrytime="00:11:04.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                    <SPLIT distance="200" swimtime="00:02:29.99" />
                    <SPLIT distance="250" swimtime="00:03:10.71" />
                    <SPLIT distance="300" swimtime="00:03:51.09" />
                    <SPLIT distance="350" swimtime="00:04:30.93" />
                    <SPLIT distance="400" swimtime="00:05:11.12" />
                    <SPLIT distance="450" swimtime="00:05:51.04" />
                    <SPLIT distance="500" swimtime="00:06:31.19" />
                    <SPLIT distance="550" swimtime="00:07:11.52" />
                    <SPLIT distance="600" swimtime="00:07:51.92" />
                    <SPLIT distance="650" swimtime="00:08:32.01" />
                    <SPLIT distance="700" swimtime="00:09:11.83" />
                    <SPLIT distance="750" swimtime="00:09:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="464" swimtime="00:01:00.59" resultid="6856" heatid="9487" lane="1" entrytime="00:01:00.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="448" reactiontime="+83" swimtime="00:00:29.30" resultid="6857" heatid="9525" lane="5" entrytime="00:00:29.60" />
                <RESULT eventid="5399" points="410" reactiontime="+79" swimtime="00:02:17.25" resultid="6858" heatid="9556" lane="2" entrytime="00:02:18.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                    <SPLIT distance="150" swimtime="00:01:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="448" reactiontime="+82" swimtime="00:00:33.91" resultid="6859" heatid="9603" lane="6" entrytime="00:00:33.68" />
                <RESULT eventid="5636" points="391" reactiontime="+78" swimtime="00:05:00.78" resultid="6860" heatid="9615" lane="3" entrytime="00:05:11.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.32" />
                    <SPLIT distance="200" swimtime="00:02:25.88" />
                    <SPLIT distance="250" swimtime="00:03:04.85" />
                    <SPLIT distance="300" swimtime="00:03:43.79" />
                    <SPLIT distance="350" swimtime="00:04:23.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="WA" clubid="5831" name="Uks Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="0-601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1990-05-19" firstname="Dawid" gender="M" lastname="Szulich" nation="POL" license="101414700035" athleteid="5832">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5585" points="693" reactiontime="+70" swimtime="00:00:29.32" resultid="5833" heatid="9605" lane="4" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" athleteid="5834">
              <RESULTS>
                <RESULT eventid="1195" points="615" reactiontime="+79" swimtime="00:00:24.58" resultid="5835" heatid="9332" lane="9" entrytime="00:00:24.77" />
                <RESULT eventid="1544" points="590" swimtime="00:00:55.90" resultid="5836" heatid="9490" lane="6" entrytime="00:00:54.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="578" reactiontime="+70" swimtime="00:01:08.57" resultid="5837" heatid="9513" lane="5" entrytime="00:01:06.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="581" reactiontime="+71" swimtime="00:00:26.87" resultid="5838" heatid="9527" lane="3" entrytime="00:00:27.25" />
                <RESULT eventid="5585" points="682" reactiontime="+68" swimtime="00:00:29.47" resultid="5839" heatid="9605" lane="2" entrytime="00:00:29.97" />
                <RESULT eventid="5636" points="342" reactiontime="+74" swimtime="00:05:14.53" resultid="5840" heatid="9614" lane="7" entrytime="00:04:56.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                    <SPLIT distance="200" swimtime="00:02:28.10" />
                    <SPLIT distance="250" swimtime="00:03:10.55" />
                    <SPLIT distance="300" swimtime="00:03:52.20" />
                    <SPLIT distance="350" swimtime="00:04:35.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-23" firstname="Krzysztof" gender="M" lastname="Żbikowski" nation="POL" athleteid="5841">
              <RESULTS>
                <RESULT eventid="1195" points="504" reactiontime="+72" swimtime="00:00:26.27" resultid="5842" heatid="9330" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1476" points="423" reactiontime="+74" swimtime="00:00:32.00" resultid="5843" heatid="9457" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1510" points="520" reactiontime="+106" swimtime="00:02:37.52" resultid="5844" heatid="9468" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="586" reactiontime="+65" swimtime="00:01:08.24" resultid="5845" heatid="9513" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="475" reactiontime="+73" swimtime="00:00:28.73" resultid="5846" heatid="9527" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="5585" points="637" reactiontime="+70" swimtime="00:00:30.15" resultid="5847" heatid="9605" lane="1" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-05" firstname="Karolina" gender="F" lastname="Modzelan" nation="POL" athleteid="5848">
              <RESULTS>
                <RESULT eventid="1133" points="426" reactiontime="+75" swimtime="00:00:31.45" resultid="5849" heatid="9315" lane="0" entrytime="00:00:29.14" />
                <RESULT eventid="1527" points="407" swimtime="00:01:09.75" resultid="5850" heatid="9475" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="378" reactiontime="+74" swimtime="00:01:28.69" resultid="5851" heatid="9503" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="397" reactiontime="+77" swimtime="00:00:40.00" resultid="5852" heatid="9595" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="7217" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="7254">
              <RESULTS>
                <RESULT eventid="1195" points="321" reactiontime="+79" swimtime="00:00:30.52" resultid="7255" heatid="9323" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1314" points="260" swimtime="00:22:44.40" resultid="7256" heatid="9366" lane="7" entrytime="00:22:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                    <SPLIT distance="200" swimtime="00:02:50.31" />
                    <SPLIT distance="250" swimtime="00:03:35.01" />
                    <SPLIT distance="300" swimtime="00:04:19.90" />
                    <SPLIT distance="350" swimtime="00:05:04.91" />
                    <SPLIT distance="400" swimtime="00:05:50.77" />
                    <SPLIT distance="450" swimtime="00:06:36.13" />
                    <SPLIT distance="500" swimtime="00:07:22.33" />
                    <SPLIT distance="550" swimtime="00:08:08.31" />
                    <SPLIT distance="600" swimtime="00:08:54.47" />
                    <SPLIT distance="650" swimtime="00:09:40.04" />
                    <SPLIT distance="700" swimtime="00:10:25.71" />
                    <SPLIT distance="750" swimtime="00:11:11.61" />
                    <SPLIT distance="800" swimtime="00:11:57.20" />
                    <SPLIT distance="850" swimtime="00:12:42.70" />
                    <SPLIT distance="900" swimtime="00:13:28.94" />
                    <SPLIT distance="950" swimtime="00:14:15.36" />
                    <SPLIT distance="1000" swimtime="00:15:02.24" />
                    <SPLIT distance="1050" swimtime="00:15:48.81" />
                    <SPLIT distance="1100" swimtime="00:16:35.26" />
                    <SPLIT distance="1150" swimtime="00:17:22.04" />
                    <SPLIT distance="1200" swimtime="00:18:08.63" />
                    <SPLIT distance="1250" swimtime="00:18:55.79" />
                    <SPLIT distance="1300" swimtime="00:19:42.35" />
                    <SPLIT distance="1350" swimtime="00:20:29.09" />
                    <SPLIT distance="1400" swimtime="00:21:15.58" />
                    <SPLIT distance="1450" swimtime="00:22:01.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="338" reactiontime="+73" swimtime="00:01:07.29" resultid="7257" heatid="9483" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="181" swimtime="00:03:16.83" resultid="7258" heatid="9494" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                    <SPLIT distance="100" swimtime="00:01:33.34" />
                    <SPLIT distance="150" swimtime="00:02:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="268" reactiontime="+74" swimtime="00:02:38.16" resultid="7259" heatid="9553" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:01:59.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="237" reactiontime="+83" swimtime="00:06:33.64" resultid="7260" heatid="9566" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:23.14" />
                    <SPLIT distance="200" swimtime="00:03:14.83" />
                    <SPLIT distance="250" swimtime="00:04:12.30" />
                    <SPLIT distance="300" swimtime="00:05:09.40" />
                    <SPLIT distance="350" swimtime="00:05:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="223" reactiontime="+95" swimtime="00:03:04.54" resultid="7261" heatid="9587" lane="9" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:18.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="283" reactiontime="+78" swimtime="00:05:34.91" resultid="7262" heatid="9616" lane="2" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:00.82" />
                    <SPLIT distance="200" swimtime="00:02:44.02" />
                    <SPLIT distance="250" swimtime="00:03:27.59" />
                    <SPLIT distance="300" swimtime="00:04:11.39" />
                    <SPLIT distance="350" swimtime="00:04:55.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="7226">
              <RESULTS>
                <RESULT eventid="1133" points="379" reactiontime="+80" swimtime="00:00:32.69" resultid="7227" heatid="9313" lane="8" entrytime="00:00:32.57" />
                <RESULT eventid="1458" points="290" reactiontime="+76" swimtime="00:00:40.87" resultid="7228" heatid="9443" lane="4" entrytime="00:00:40.27" />
                <RESULT eventid="1527" points="365" reactiontime="+69" swimtime="00:01:12.34" resultid="7229" heatid="9474" lane="5" entrytime="00:01:11.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="243" swimtime="00:00:39.13" resultid="7230" heatid="9515" lane="3" entrytime="00:00:37.39" />
                <RESULT eventid="5382" points="293" swimtime="00:02:50.09" resultid="7231" heatid="9545" lane="6" entrytime="00:02:50.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:02:07.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="234" reactiontime="+93" swimtime="00:01:29.92" resultid="7232" heatid="9570" lane="5" entrytime="00:01:28.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="269" swimtime="00:00:45.49" resultid="7233" heatid="9594" lane="7" entrytime="00:00:44.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="7270">
              <RESULTS>
                <RESULT eventid="1133" points="331" reactiontime="+92" swimtime="00:00:34.21" resultid="7271" heatid="9312" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1212" points="301" reactiontime="+77" swimtime="00:03:08.18" resultid="7272" heatid="9339" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:30.56" />
                    <SPLIT distance="150" swimtime="00:02:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="270" reactiontime="+91" swimtime="00:00:41.82" resultid="7273" heatid="9444" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1493" points="262" swimtime="00:03:37.24" resultid="7274" heatid="9460" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:01:44.90" />
                    <SPLIT distance="150" swimtime="00:02:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="282" swimtime="00:01:37.69" resultid="7275" heatid="9502" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5450" points="246" swimtime="00:07:04.92" resultid="7276" heatid="9563" lane="9" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:38.05" />
                    <SPLIT distance="150" swimtime="00:02:32.77" />
                    <SPLIT distance="200" swimtime="00:03:25.37" />
                    <SPLIT distance="250" swimtime="00:04:26.22" />
                    <SPLIT distance="300" swimtime="00:05:26.70" />
                    <SPLIT distance="350" swimtime="00:06:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="184" reactiontime="+94" swimtime="00:01:37.45" resultid="7277" heatid="9570" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="302" reactiontime="+83" swimtime="00:00:43.79" resultid="7278" heatid="9594" lane="2" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="7238">
              <RESULTS>
                <RESULT eventid="1229" points="296" swimtime="00:02:50.96" resultid="7239" heatid="9346" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:02:09.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="213" reactiontime="+79" swimtime="00:12:36.80" resultid="7240" heatid="9360" lane="8" entrytime="00:11:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:19.80" />
                    <SPLIT distance="150" swimtime="00:02:05.28" />
                    <SPLIT distance="200" swimtime="00:02:53.12" />
                    <SPLIT distance="250" swimtime="00:03:41.71" />
                    <SPLIT distance="300" swimtime="00:04:30.45" />
                    <SPLIT distance="350" swimtime="00:05:19.28" />
                    <SPLIT distance="400" swimtime="00:06:08.73" />
                    <SPLIT distance="450" swimtime="00:06:57.82" />
                    <SPLIT distance="500" swimtime="00:07:47.45" />
                    <SPLIT distance="550" swimtime="00:08:36.67" />
                    <SPLIT distance="600" swimtime="00:09:25.93" />
                    <SPLIT distance="650" swimtime="00:10:14.84" />
                    <SPLIT distance="700" swimtime="00:11:03.12" />
                    <SPLIT distance="750" swimtime="00:11:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="332" reactiontime="+79" swimtime="00:03:02.84" resultid="7241" heatid="9467" lane="3" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:13.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="346" reactiontime="+74" swimtime="00:01:21.35" resultid="7242" heatid="9511" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="7243" heatid="9523" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="5585" points="377" reactiontime="+72" swimtime="00:00:35.92" resultid="7244" heatid="9602" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="7218">
              <RESULTS>
                <RESULT eventid="1263" points="315" swimtime="00:11:52.38" resultid="7219" heatid="9355" lane="7" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                    <SPLIT distance="200" swimtime="00:02:50.87" />
                    <SPLIT distance="250" swimtime="00:03:36.00" />
                    <SPLIT distance="300" swimtime="00:04:21.53" />
                    <SPLIT distance="350" swimtime="00:05:06.68" />
                    <SPLIT distance="400" swimtime="00:05:52.10" />
                    <SPLIT distance="450" swimtime="00:06:37.71" />
                    <SPLIT distance="500" swimtime="00:07:23.86" />
                    <SPLIT distance="550" swimtime="00:08:09.13" />
                    <SPLIT distance="600" swimtime="00:08:54.67" />
                    <SPLIT distance="650" swimtime="00:09:40.03" />
                    <SPLIT distance="700" swimtime="00:10:25.59" />
                    <SPLIT distance="750" swimtime="00:11:10.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="316" reactiontime="+75" swimtime="00:00:39.70" resultid="7220" heatid="9444" lane="7" entrytime="00:00:39.50" />
                <RESULT eventid="1527" points="350" swimtime="00:01:13.34" resultid="7221" heatid="9474" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="344" reactiontime="+72" swimtime="00:01:22.90" resultid="7222" heatid="9532" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="327" reactiontime="+88" swimtime="00:02:43.91" resultid="7223" heatid="9546" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" points="359" reactiontime="+74" swimtime="00:02:54.46" resultid="7224" heatid="9582" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="317" reactiontime="+87" swimtime="00:05:46.49" resultid="7225" heatid="9609" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:21.62" />
                    <SPLIT distance="150" swimtime="00:02:05.74" />
                    <SPLIT distance="200" swimtime="00:02:50.10" />
                    <SPLIT distance="250" swimtime="00:03:35.26" />
                    <SPLIT distance="300" swimtime="00:04:20.06" />
                    <SPLIT distance="350" swimtime="00:05:04.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="7246">
              <RESULTS>
                <RESULT eventid="1195" points="335" reactiontime="+81" swimtime="00:00:30.10" resultid="7247" heatid="9326" lane="6" entrytime="00:00:28.99" />
                <RESULT eventid="1510" points="287" reactiontime="+76" swimtime="00:03:11.86" resultid="7248" heatid="9467" lane="8" entrytime="00:02:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:22.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="7249" heatid="9486" lane="9" entrytime="00:01:03.79" />
                <RESULT eventid="5297" points="284" reactiontime="+77" swimtime="00:01:26.89" resultid="7250" heatid="9510" lane="3" entrytime="00:01:21.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="7251" heatid="9523" lane="0" entrytime="00:00:32.07" />
                <RESULT eventid="5585" points="324" reactiontime="+79" swimtime="00:00:37.78" resultid="7252" heatid="9602" lane="1" entrytime="00:00:36.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="7234">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1195" status="DSQ" swimtime="00:00:26.84" resultid="7235" heatid="9323" lane="3" entrytime="00:00:30.34" />
                <RESULT eventid="1544" points="468" reactiontime="+86" swimtime="00:01:00.42" resultid="7236" heatid="9485" lane="0" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="429" reactiontime="+86" swimtime="00:02:15.21" resultid="7237" heatid="9555" lane="3" entrytime="00:02:22.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:41.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="7263">
              <RESULTS>
                <RESULT eventid="1314" status="OTL" swimtime="00:21:04.03" resultid="7264" heatid="9365" lane="7" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:55.15" />
                    <SPLIT distance="200" swimtime="00:02:36.35" />
                    <SPLIT distance="250" swimtime="00:03:18.24" />
                    <SPLIT distance="300" swimtime="00:04:01.20" />
                    <SPLIT distance="350" swimtime="00:04:43.99" />
                    <SPLIT distance="400" swimtime="00:05:26.75" />
                    <SPLIT distance="450" swimtime="00:06:08.52" />
                    <SPLIT distance="500" swimtime="00:06:51.25" />
                    <SPLIT distance="550" swimtime="00:07:33.91" />
                    <SPLIT distance="600" swimtime="00:08:16.31" />
                    <SPLIT distance="650" swimtime="00:08:58.14" />
                    <SPLIT distance="700" swimtime="00:09:40.68" />
                    <SPLIT distance="750" swimtime="00:10:22.51" />
                    <SPLIT distance="800" swimtime="00:11:04.86" />
                    <SPLIT distance="850" swimtime="00:11:47.28" />
                    <SPLIT distance="900" swimtime="00:12:30.43" />
                    <SPLIT distance="950" swimtime="00:13:13.32" />
                    <SPLIT distance="1000" swimtime="00:13:56.50" />
                    <SPLIT distance="1050" swimtime="00:14:39.86" />
                    <SPLIT distance="1100" swimtime="00:15:23.13" />
                    <SPLIT distance="1150" swimtime="00:16:06.47" />
                    <SPLIT distance="1200" swimtime="00:16:49.59" />
                    <SPLIT distance="1250" swimtime="00:17:32.45" />
                    <SPLIT distance="1300" swimtime="00:18:15.18" />
                    <SPLIT distance="1350" swimtime="00:18:57.84" />
                    <SPLIT distance="1400" swimtime="00:19:40.00" />
                    <SPLIT distance="1450" swimtime="00:20:22.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="454" reactiontime="+72" swimtime="00:02:44.75" resultid="7265" heatid="9468" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                    <SPLIT distance="150" swimtime="00:02:02.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="411" reactiontime="+67" swimtime="00:01:16.80" resultid="7266" heatid="9513" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="7267" heatid="9567" lane="0" entrytime="00:06:00.00" />
                <RESULT eventid="5585" points="437" reactiontime="+85" swimtime="00:00:34.19" resultid="7268" heatid="9605" lane="8" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="338" reactiontime="+92" swimtime="00:02:14.12" resultid="7281" heatid="9499" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7254" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="7263" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="7246" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="7238" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5433" points="373" swimtime="00:01:57.86" resultid="7282" heatid="9561" lane="1" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="100" swimtime="00:01:00.50" />
                    <SPLIT distance="150" swimtime="00:01:30.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7238" number="1" />
                    <RELAYPOSITION athleteid="7254" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="7246" number="3" />
                    <RELAYPOSITION athleteid="7263" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+78" swimtime="00:02:04.76" resultid="7279" heatid="9354" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:02.10" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7238" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="7226" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="7246" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="7218" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="5602" reactiontime="+76" swimtime="00:02:20.23" resultid="7280" heatid="9608" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:01:47.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7218" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="7238" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="7246" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="7226" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="6407" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska 2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="6408">
              <RESULTS>
                <RESULT eventid="1229" points="78" swimtime="00:04:25.70" resultid="6409" heatid="9343" lane="6" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.09" />
                    <SPLIT distance="100" swimtime="00:02:06.29" />
                    <SPLIT distance="150" swimtime="00:03:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="90" reactiontime="+104" swimtime="00:16:46.29" resultid="6410" heatid="9363" lane="4" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.59" />
                    <SPLIT distance="100" swimtime="00:01:59.29" />
                    <SPLIT distance="150" swimtime="00:03:04.71" />
                    <SPLIT distance="200" swimtime="00:04:09.38" />
                    <SPLIT distance="250" swimtime="00:05:14.49" />
                    <SPLIT distance="300" swimtime="00:06:18.94" />
                    <SPLIT distance="350" swimtime="00:07:24.00" />
                    <SPLIT distance="400" swimtime="00:08:27.62" />
                    <SPLIT distance="450" swimtime="00:09:32.18" />
                    <SPLIT distance="500" swimtime="00:10:36.65" />
                    <SPLIT distance="550" swimtime="00:11:40.25" />
                    <SPLIT distance="600" swimtime="00:12:42.05" />
                    <SPLIT distance="650" swimtime="00:13:43.68" />
                    <SPLIT distance="700" swimtime="00:14:45.83" />
                    <SPLIT distance="750" swimtime="00:15:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="78" swimtime="00:04:55.38" resultid="6411" heatid="9463" lane="9" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.73" />
                    <SPLIT distance="100" swimtime="00:02:23.98" />
                    <SPLIT distance="150" swimtime="00:03:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="52" swimtime="00:04:58.75" resultid="6412" heatid="9493" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.27" />
                    <SPLIT distance="100" swimtime="00:02:25.03" />
                    <SPLIT distance="150" swimtime="00:03:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="75" reactiontime="+83" swimtime="00:02:02.42" resultid="6413" heatid="9535" lane="3" entrytime="00:01:55.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="80" reactiontime="+92" swimtime="00:09:25.23" resultid="6414" heatid="9564" lane="4" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.86" />
                    <SPLIT distance="100" swimtime="00:02:24.32" />
                    <SPLIT distance="150" swimtime="00:03:35.99" />
                    <SPLIT distance="200" swimtime="00:04:44.47" />
                    <SPLIT distance="250" swimtime="00:06:02.78" />
                    <SPLIT distance="300" swimtime="00:07:24.40" />
                    <SPLIT distance="350" swimtime="00:08:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="49" swimtime="00:02:15.36" resultid="6415" heatid="9572" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="89" reactiontime="+79" swimtime="00:04:09.99" resultid="6416" heatid="9585" lane="0" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.41" />
                    <SPLIT distance="100" swimtime="00:02:05.67" />
                    <SPLIT distance="150" swimtime="00:03:10.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="107414" nation="POL" region="OL" clubid="6092" name="UKS Manta Warszawa Włochy">
          <CONTACT name="Barański" phone="510835478" />
          <ATHLETES>
            <ATHLETE birthdate="1993-09-09" firstname="Michał" gender="M" lastname="Bielawski" nation="POL" license="107414700127" athleteid="6093">
              <RESULTS>
                <RESULT eventid="1195" points="642" reactiontime="+66" swimtime="00:00:24.23" resultid="6094" heatid="9332" lane="4" entrytime="00:00:23.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1544" points="740" reactiontime="+61" swimtime="00:00:51.85" resultid="6095" heatid="9490" lane="4" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02201" nation="POL" region="DOL" clubid="6559" name="Uks Shark Rudna">
          <CONTACT name="SZAJNICKI" />
          <ATHLETES>
            <ATHLETE birthdate="1995-07-19" firstname="Katarzyna" gender="F" lastname="Kita" nation="POL" license="102201600078" athleteid="6569">
              <RESULTS>
                <RESULT eventid="1133" points="650" reactiontime="+67" swimtime="00:00:27.32" resultid="6570" heatid="9315" lane="4" entrytime="00:00:26.82" />
                <RESULT eventid="1458" points="412" reactiontime="+85" swimtime="00:00:36.35" resultid="6571" heatid="9445" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1527" points="630" reactiontime="+66" swimtime="00:01:00.29" resultid="6572" heatid="9476" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="420" reactiontime="+75" swimtime="00:00:32.62" resultid="6573" heatid="9517" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="5382" points="552" reactiontime="+69" swimtime="00:02:17.65" resultid="6574" heatid="9547" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                    <SPLIT distance="150" swimtime="00:01:43.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-11" firstname="Agnieszka" gender="F" lastname="Gajdowska" nation="POL" license="102201600071" athleteid="6560">
              <RESULTS>
                <RESULT eventid="1133" points="555" swimtime="00:00:28.80" resultid="6561" heatid="9315" lane="3" entrytime="00:00:27.89" />
                <RESULT eventid="1212" points="440" swimtime="00:02:45.80" resultid="6562" heatid="9340" lane="1" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="150" swimtime="00:02:07.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="464" reactiontime="+75" swimtime="00:00:34.93" resultid="6563" heatid="9446" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1527" points="587" swimtime="00:01:01.75" resultid="6564" heatid="9476" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="478" reactiontime="+74" swimtime="00:00:31.23" resultid="6565" heatid="9517" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="5382" points="489" reactiontime="+68" swimtime="00:02:23.39" resultid="6566" heatid="9547" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="410" reactiontime="+70" swimtime="00:00:39.57" resultid="6567" heatid="9596" lane="2" entrytime="00:00:36.78" />
                <RESULT eventid="5619" points="462" reactiontime="+69" swimtime="00:05:05.73" resultid="6568" heatid="9609" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:53.56" />
                    <SPLIT distance="200" swimtime="00:02:33.63" />
                    <SPLIT distance="250" swimtime="00:03:12.78" />
                    <SPLIT distance="300" swimtime="00:03:51.63" />
                    <SPLIT distance="350" swimtime="00:04:30.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SP8" nation="POL" region="MAL" clubid="5715" name="UKS SP 8 Chrzanow">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański" phone="692076808" state="MAŁ" street="Niepodległości 7 / 46" zip="32 500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="5716">
              <RESULTS>
                <RESULT eventid="1195" points="275" reactiontime="+92" swimtime="00:00:32.15" resultid="5717" heatid="9322" lane="1" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1280" points="167" reactiontime="+107" swimtime="00:13:40.92" resultid="5718" heatid="9361" lane="8" entrytime="00:13:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                    <SPLIT distance="200" swimtime="00:03:14.24" />
                    <SPLIT distance="250" swimtime="00:04:07.32" />
                    <SPLIT distance="300" swimtime="00:04:59.48" />
                    <SPLIT distance="350" swimtime="00:05:52.00" />
                    <SPLIT distance="400" swimtime="00:06:43.96" />
                    <SPLIT distance="450" swimtime="00:07:36.37" />
                    <SPLIT distance="500" swimtime="00:08:29.10" />
                    <SPLIT distance="550" swimtime="00:09:22.24" />
                    <SPLIT distance="600" swimtime="00:10:15.11" />
                    <SPLIT distance="650" swimtime="00:11:08.15" />
                    <SPLIT distance="700" swimtime="00:12:01.64" />
                    <SPLIT distance="750" swimtime="00:12:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="172" reactiontime="+79" swimtime="00:00:43.20" resultid="5719" heatid="9451" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1544" points="265" reactiontime="+94" swimtime="00:01:12.99" resultid="5720" heatid="9481" lane="4" entrytime="00:01:13.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="204" swimtime="00:02:53.24" resultid="5721" heatid="9552" lane="1" entrytime="00:02:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:09.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="176" reactiontime="+96" swimtime="00:06:32.46" resultid="5722" heatid="9617" lane="8" entrytime="00:06:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:31.18" />
                    <SPLIT distance="150" swimtime="00:02:20.77" />
                    <SPLIT distance="200" swimtime="00:03:10.98" />
                    <SPLIT distance="250" swimtime="00:04:01.48" />
                    <SPLIT distance="300" swimtime="00:04:51.58" />
                    <SPLIT distance="350" swimtime="00:05:43.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPOOB" nation="POL" region="WIE" clubid="5817" name="UKS Sportowiec Oborniki">
          <CONTACT city="Oborniki" email="ukssportowiec.oborniki@gmail.com" name="Kolendowicz" phone="606267334" state="WIE" street="Czarnkowska  57" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1988-05-16" firstname="Łukasz" gender="M" lastname="Kolendowicz" nation="POL" license="505715700037" athleteid="5818">
              <RESULTS>
                <RESULT eventid="1314" points="411" reactiontime="+97" swimtime="00:19:31.14" resultid="5819" heatid="9365" lane="5" entrytime="00:18:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                    <SPLIT distance="200" swimtime="00:02:24.14" />
                    <SPLIT distance="250" swimtime="00:03:02.01" />
                    <SPLIT distance="300" swimtime="00:03:40.50" />
                    <SPLIT distance="350" swimtime="00:04:19.44" />
                    <SPLIT distance="400" swimtime="00:04:58.33" />
                    <SPLIT distance="450" swimtime="00:05:37.81" />
                    <SPLIT distance="500" swimtime="00:06:17.27" />
                    <SPLIT distance="550" swimtime="00:06:56.82" />
                    <SPLIT distance="600" swimtime="00:07:36.69" />
                    <SPLIT distance="650" swimtime="00:08:16.43" />
                    <SPLIT distance="700" swimtime="00:08:56.38" />
                    <SPLIT distance="750" swimtime="00:09:36.18" />
                    <SPLIT distance="800" swimtime="00:10:16.19" />
                    <SPLIT distance="850" swimtime="00:10:56.21" />
                    <SPLIT distance="900" swimtime="00:11:35.94" />
                    <SPLIT distance="950" swimtime="00:12:15.98" />
                    <SPLIT distance="1000" swimtime="00:12:56.06" />
                    <SPLIT distance="1050" swimtime="00:13:36.37" />
                    <SPLIT distance="1100" swimtime="00:14:16.74" />
                    <SPLIT distance="1150" swimtime="00:14:56.54" />
                    <SPLIT distance="1200" swimtime="00:15:36.51" />
                    <SPLIT distance="1250" swimtime="00:16:15.81" />
                    <SPLIT distance="1300" swimtime="00:16:55.62" />
                    <SPLIT distance="1350" swimtime="00:17:35.18" />
                    <SPLIT distance="1400" swimtime="00:18:14.21" />
                    <SPLIT distance="1450" swimtime="00:18:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" reactiontime="+95" status="DNS" swimtime="00:00:00.00" resultid="5821" heatid="9613" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRCZ" nation="POL" clubid="5673" name="UKS Trójka Częstochowa">
          <ATHLETES>
            <ATHLETE birthdate="1995-06-07" firstname="Mateusz" gender="M" lastname="Chowaniec" nation="POL" license="100111700079" athleteid="5672">
              <RESULTS>
                <RESULT eventid="1195" points="493" reactiontime="+74" swimtime="00:00:26.46" resultid="5674" heatid="9329" lane="2" entrytime="00:00:26.69" />
                <RESULT eventid="1229" points="370" reactiontime="+75" swimtime="00:02:38.71" resultid="5675" heatid="9342" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:58.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="419" swimtime="00:02:49.15" resultid="5676" heatid="9462" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:20.53" />
                    <SPLIT distance="150" swimtime="00:02:05.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="467" reactiontime="+69" swimtime="00:01:13.60" resultid="5677" heatid="9512" lane="2" entrytime="00:01:13.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="346" reactiontime="+75" swimtime="00:00:31.94" resultid="5678" heatid="9518" lane="3" />
                <RESULT eventid="5585" points="518" reactiontime="+73" swimtime="00:00:32.31" resultid="5679" heatid="9604" lane="8" entrytime="00:00:32.92" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="KA" clubid="7985" name="UKS Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="8025">
              <RESULTS>
                <RESULT eventid="1195" points="290" reactiontime="+89" swimtime="00:00:31.59" resultid="8026" heatid="9322" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1510" points="300" reactiontime="+93" swimtime="00:03:09.04" resultid="8027" heatid="9466" lane="8" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:30.35" />
                    <SPLIT distance="150" swimtime="00:02:19.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="316" reactiontime="+84" swimtime="00:01:23.84" resultid="8028" heatid="9510" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="364" reactiontime="+90" swimtime="00:00:36.32" resultid="8029" heatid="9602" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="8020">
              <RESULTS>
                <RESULT eventid="1195" points="328" reactiontime="+108" swimtime="00:00:30.30" resultid="8021" heatid="9325" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1544" points="286" reactiontime="+101" swimtime="00:01:11.14" resultid="8022" heatid="9483" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5331" points="341" reactiontime="+102" swimtime="00:00:32.10" resultid="8023" heatid="9523" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="5517" points="240" swimtime="00:01:20.10" resultid="8024" heatid="9575" lane="1" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="8006">
              <RESULTS>
                <RESULT eventid="1458" status="DNS" swimtime="00:00:00.00" resultid="8008" heatid="9441" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="8009" heatid="9530" lane="3" entrytime="00:02:05.00" />
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="8010" heatid="9580" lane="9" entrytime="00:04:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="8011">
              <RESULTS>
                <RESULT eventid="1195" points="359" reactiontime="+86" swimtime="00:00:29.40" resultid="8012" heatid="9325" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1280" points="289" reactiontime="+103" swimtime="00:11:23.40" resultid="8013" heatid="9360" lane="5" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:55.61" />
                    <SPLIT distance="200" swimtime="00:02:38.62" />
                    <SPLIT distance="250" swimtime="00:03:22.01" />
                    <SPLIT distance="300" swimtime="00:04:05.81" />
                    <SPLIT distance="350" swimtime="00:04:49.75" />
                    <SPLIT distance="400" swimtime="00:05:34.03" />
                    <SPLIT distance="450" swimtime="00:06:18.20" />
                    <SPLIT distance="500" swimtime="00:07:01.03" />
                    <SPLIT distance="550" swimtime="00:07:45.05" />
                    <SPLIT distance="600" swimtime="00:08:28.91" />
                    <SPLIT distance="650" swimtime="00:09:13.18" />
                    <SPLIT distance="700" swimtime="00:09:56.78" />
                    <SPLIT distance="750" swimtime="00:10:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G2 - Pływak zanurzył się całkowicie w trakcie wyścigu (z wyjątkiem 15 m po starcie lub nawrocie)." eventid="1476" reactiontime="+96" status="DSQ" swimtime="00:00:37.75" resultid="8014" heatid="9453" lane="9" entrytime="00:00:36.50" />
                <RESULT eventid="1544" points="352" reactiontime="+89" swimtime="00:01:06.39" resultid="8015" heatid="9484" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="260" reactiontime="+98" swimtime="00:01:21.22" resultid="8016" heatid="9538" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="292" reactiontime="+95" swimtime="00:02:33.71" resultid="8017" heatid="9555" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="234" reactiontime="+96" swimtime="00:03:01.38" resultid="8018" heatid="9587" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:26.95" />
                    <SPLIT distance="150" swimtime="00:02:14.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="279" reactiontime="+81" swimtime="00:05:36.45" resultid="8019" heatid="9615" lane="8" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                    <SPLIT distance="200" swimtime="00:02:42.55" />
                    <SPLIT distance="250" swimtime="00:03:26.47" />
                    <SPLIT distance="300" swimtime="00:04:10.56" />
                    <SPLIT distance="350" swimtime="00:04:54.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01711" nation="POL" region="11" clubid="6118" name="UKS WODNIK Siemianowice Ślaskie" shortname="UKS WODNIK Siemianowice Ślaski">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek Leszek" phone="534033934" state="ŚLĄSK" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="6119">
              <RESULTS>
                <RESULT eventid="1229" points="228" swimtime="00:03:06.56" resultid="6120" heatid="9344" lane="1" entrytime="00:03:15.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:29.49" />
                    <SPLIT distance="150" swimtime="00:02:24.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="229" reactiontime="+72" swimtime="00:23:42.82" resultid="6121" heatid="9366" lane="0" entrytime="00:23:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:02:16.05" />
                    <SPLIT distance="200" swimtime="00:03:04.50" />
                    <SPLIT distance="250" swimtime="00:03:54.32" />
                    <SPLIT distance="300" swimtime="00:04:43.03" />
                    <SPLIT distance="350" swimtime="00:05:31.66" />
                    <SPLIT distance="400" swimtime="00:06:19.55" />
                    <SPLIT distance="450" swimtime="00:07:06.74" />
                    <SPLIT distance="500" swimtime="00:07:55.36" />
                    <SPLIT distance="550" swimtime="00:08:43.53" />
                    <SPLIT distance="600" swimtime="00:09:31.05" />
                    <SPLIT distance="650" swimtime="00:10:18.62" />
                    <SPLIT distance="700" swimtime="00:11:05.81" />
                    <SPLIT distance="750" swimtime="00:11:53.45" />
                    <SPLIT distance="800" swimtime="00:12:41.60" />
                    <SPLIT distance="850" swimtime="00:13:30.54" />
                    <SPLIT distance="900" swimtime="00:14:17.81" />
                    <SPLIT distance="950" swimtime="00:15:05.93" />
                    <SPLIT distance="1000" swimtime="00:15:53.36" />
                    <SPLIT distance="1050" swimtime="00:16:40.54" />
                    <SPLIT distance="1100" swimtime="00:17:27.62" />
                    <SPLIT distance="1150" swimtime="00:18:14.33" />
                    <SPLIT distance="1200" swimtime="00:19:01.44" />
                    <SPLIT distance="1250" swimtime="00:19:48.66" />
                    <SPLIT distance="1300" swimtime="00:20:35.48" />
                    <SPLIT distance="1350" swimtime="00:21:22.63" />
                    <SPLIT distance="1400" swimtime="00:22:09.91" />
                    <SPLIT distance="1450" swimtime="00:22:57.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="151" reactiontime="+48" swimtime="00:03:29.01" resultid="6122" heatid="9494" lane="7" entrytime="00:03:24.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:39.76" />
                    <SPLIT distance="150" swimtime="00:02:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="6123" heatid="9521" lane="1" entrytime="00:00:36.60" />
                <RESULT eventid="5467" points="207" swimtime="00:06:51.71" resultid="6124" heatid="9566" lane="1" entrytime="00:06:31.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                    <SPLIT distance="150" swimtime="00:02:31.62" />
                    <SPLIT distance="200" swimtime="00:03:24.86" />
                    <SPLIT distance="250" swimtime="00:04:23.53" />
                    <SPLIT distance="300" swimtime="00:05:22.99" />
                    <SPLIT distance="350" swimtime="00:06:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6125" heatid="9574" lane="9" entrytime="00:01:27.40" />
                <RESULT eventid="5636" points="214" swimtime="00:06:07.63" resultid="6126" heatid="9616" lane="9" entrytime="00:05:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:13.48" />
                    <SPLIT distance="200" swimtime="00:03:00.77" />
                    <SPLIT distance="250" swimtime="00:03:48.26" />
                    <SPLIT distance="300" swimtime="00:04:36.25" />
                    <SPLIT distance="350" swimtime="00:05:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="6183" name="Unia Oświęcim Masters">
          <ATHLETES>
            <ATHLETE birthdate="1952-07-01" firstname="Barbara" gender="F" lastname="Lipniarska-Skubis" nation="POL" license="501006600377" athleteid="6184">
              <RESULTS>
                <RESULT eventid="1263" points="94" swimtime="00:17:45.94" resultid="6185" heatid="9357" lane="7" entrytime="00:18:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                    <SPLIT distance="100" swimtime="00:01:59.63" />
                    <SPLIT distance="150" swimtime="00:03:06.56" />
                    <SPLIT distance="200" swimtime="00:04:13.15" />
                    <SPLIT distance="250" swimtime="00:05:20.94" />
                    <SPLIT distance="300" swimtime="00:06:27.81" />
                    <SPLIT distance="350" swimtime="00:07:35.84" />
                    <SPLIT distance="400" swimtime="00:08:43.07" />
                    <SPLIT distance="450" swimtime="00:09:51.16" />
                    <SPLIT distance="500" swimtime="00:10:58.37" />
                    <SPLIT distance="550" swimtime="00:12:08.06" />
                    <SPLIT distance="600" swimtime="00:13:15.47" />
                    <SPLIT distance="650" swimtime="00:14:24.38" />
                    <SPLIT distance="700" swimtime="00:15:31.47" />
                    <SPLIT distance="750" swimtime="00:16:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="87" swimtime="00:01:56.32" resultid="6186" heatid="9470" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="84" reactiontime="+99" swimtime="00:04:17.32" resultid="6187" heatid="9542" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.05" />
                    <SPLIT distance="100" swimtime="00:02:01.60" />
                    <SPLIT distance="150" swimtime="00:03:10.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="97" swimtime="00:08:32.98" resultid="6188" heatid="9612" lane="2" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.08" />
                    <SPLIT distance="100" swimtime="00:02:00.93" />
                    <SPLIT distance="150" swimtime="00:03:06.51" />
                    <SPLIT distance="200" swimtime="00:04:12.88" />
                    <SPLIT distance="250" swimtime="00:05:18.17" />
                    <SPLIT distance="300" swimtime="00:06:24.48" />
                    <SPLIT distance="350" swimtime="00:07:29.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="6540" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="6541">
              <RESULTS>
                <RESULT eventid="1195" points="361" reactiontime="+77" swimtime="00:00:29.34" resultid="6542" heatid="9325" lane="1" entrytime="00:00:29.30" />
                <RESULT eventid="1544" points="369" reactiontime="+88" swimtime="00:01:05.37" resultid="6543" heatid="9484" lane="5" entrytime="00:01:04.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="325" reactiontime="+93" swimtime="00:00:32.60" resultid="6544" heatid="9521" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="5399" points="309" reactiontime="+79" swimtime="00:02:30.72" resultid="6545" heatid="9554" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6546" heatid="9574" lane="1" entrytime="00:01:26.00" />
                <RESULT eventid="5636" points="300" reactiontime="+83" swimtime="00:05:28.65" resultid="6547" heatid="9616" lane="5" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:15.94" />
                    <SPLIT distance="150" swimtime="00:01:58.21" />
                    <SPLIT distance="200" swimtime="00:02:41.77" />
                    <SPLIT distance="250" swimtime="00:03:24.80" />
                    <SPLIT distance="300" swimtime="00:04:07.20" />
                    <SPLIT distance="350" swimtime="00:04:49.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031/05" nation="POL" region="LOD" clubid="6189" name="UTW &quot;Masters&quot; Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1949-02-07" firstname="Krzysztof" gender="M" lastname="Wojciechowski" nation="POL" license="503105700024" athleteid="6224">
              <RESULTS>
                <RESULT eventid="1510" points="171" swimtime="00:03:47.80" resultid="6225" heatid="9464" lane="9" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                    <SPLIT distance="100" swimtime="00:01:49.30" />
                    <SPLIT distance="150" swimtime="00:02:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="194" reactiontime="+96" swimtime="00:01:38.57" resultid="6226" heatid="9508" lane="0" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="236" reactiontime="+98" swimtime="00:00:41.95" resultid="6227" heatid="9599" lane="1" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-03" firstname="Yuriy" gender="M" lastname="Danylchenko" nation="POL" license="503105700" athleteid="6255">
              <RESULTS>
                <RESULT eventid="1195" points="256" reactiontime="+109" swimtime="00:00:32.91" resultid="6256" heatid="9321" lane="7" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1314" reactiontime="+103" status="OTL" swimtime="00:00:00.00" resultid="6257" heatid="9368" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:01:31.50" />
                    <SPLIT distance="150" swimtime="00:02:27.78" />
                    <SPLIT distance="200" swimtime="00:03:25.22" />
                    <SPLIT distance="250" swimtime="00:04:24.29" />
                    <SPLIT distance="300" swimtime="00:05:22.23" />
                    <SPLIT distance="350" swimtime="00:06:20.63" />
                    <SPLIT distance="400" swimtime="00:07:19.96" />
                    <SPLIT distance="450" swimtime="00:08:18.20" />
                    <SPLIT distance="500" swimtime="00:09:16.36" />
                    <SPLIT distance="550" swimtime="00:10:14.97" />
                    <SPLIT distance="600" swimtime="00:11:15.63" />
                    <SPLIT distance="650" swimtime="00:12:14.34" />
                    <SPLIT distance="700" swimtime="00:13:13.27" />
                    <SPLIT distance="750" swimtime="00:14:14.65" />
                    <SPLIT distance="800" swimtime="00:15:13.64" />
                    <SPLIT distance="850" swimtime="00:16:13.93" />
                    <SPLIT distance="900" swimtime="00:17:12.38" />
                    <SPLIT distance="950" swimtime="00:18:12.65" />
                    <SPLIT distance="1000" swimtime="00:19:11.91" />
                    <SPLIT distance="1050" swimtime="00:20:12.23" />
                    <SPLIT distance="1100" swimtime="00:21:11.16" />
                    <SPLIT distance="1150" swimtime="00:22:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6258" heatid="9481" lane="2" entrytime="00:01:15.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="6190">
              <RESULTS>
                <RESULT eventid="1476" points="158" reactiontime="+82" swimtime="00:00:44.40" resultid="6191" heatid="9450" lane="1" entrytime="00:00:46.00" entrycourse="LCM" />
                <RESULT eventid="1510" points="209" reactiontime="+102" swimtime="00:03:33.32" resultid="6192" heatid="9464" lane="2" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.62" />
                    <SPLIT distance="100" swimtime="00:01:43.85" />
                    <SPLIT distance="150" swimtime="00:02:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="208" swimtime="00:01:36.36" resultid="6193" heatid="9508" lane="1" entrytime="00:01:34.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="152" reactiontime="+86" swimtime="00:01:36.97" resultid="6194" heatid="9536" lane="7" entrytime="00:01:37.00" entrycourse="LCM" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5551" points="154" reactiontime="+86" swimtime="00:03:28.71" resultid="6195" heatid="9585" lane="3" entrytime="00:03:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="231" reactiontime="+100" swimtime="00:00:42.29" resultid="6196" heatid="9599" lane="5" entrytime="00:00:41.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-06" firstname="Robert" gender="M" lastname="Szalbierz" nation="POL" license="503105700056" athleteid="6197">
              <RESULTS>
                <RESULT eventid="1195" points="311" reactiontime="+46" swimtime="00:00:30.83" resultid="6198" heatid="9324" lane="3" entrytime="00:00:29.60" entrycourse="LCM" />
                <RESULT eventid="1544" points="300" swimtime="00:01:10.06" resultid="6199" heatid="9483" lane="9" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="296" reactiontime="+94" swimtime="00:00:33.63" resultid="6200" heatid="9522" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6201" heatid="9575" lane="9" entrytime="00:01:20.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Woźniak" nation="POL" license="503157000390" athleteid="6263">
              <RESULTS>
                <RESULT eventid="1476" points="470" reactiontime="+59" swimtime="00:00:30.91" resultid="6264" heatid="9456" lane="1" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="5331" points="479" reactiontime="+76" swimtime="00:00:28.66" resultid="6265" heatid="9518" lane="6" />
                <RESULT eventid="5365" points="452" reactiontime="+59" swimtime="00:01:07.56" resultid="6266" heatid="9540" lane="5" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="413" reactiontime="+79" swimtime="00:01:06.85" resultid="6267" heatid="9572" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="420" reactiontime="+61" swimtime="00:02:29.36" resultid="6268" heatid="9590" lane="2" entrytime="00:02:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:50.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="6228">
              <RESULTS>
                <RESULT eventid="1212" points="450" reactiontime="+83" swimtime="00:02:44.54" resultid="6229" heatid="9339" lane="4" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1458" points="385" reactiontime="+79" swimtime="00:00:37.17" resultid="6230" heatid="9445" lane="4" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1561" points="334" reactiontime="+87" swimtime="00:02:55.39" resultid="6231" heatid="9492" lane="3" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.67" />
                    <SPLIT distance="150" swimtime="00:02:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas równy Rekordowi Polski" eventid="5314" points="432" swimtime="00:00:32.30" resultid="6232" heatid="9516" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="5348" points="355" reactiontime="+83" swimtime="00:01:22.01" resultid="6233" heatid="9533" lane="2" entrytime="00:01:13.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="446" reactiontime="+80" swimtime="00:01:12.61" resultid="6234" heatid="9571" lane="2" entrytime="00:01:13.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="6269">
              <RESULTS>
                <RESULT eventid="1133" points="365" reactiontime="+86" swimtime="00:00:33.12" resultid="6270" heatid="9313" lane="1" entrytime="00:00:32.40" entrycourse="LCM" />
                <RESULT eventid="1458" points="323" reactiontime="+77" swimtime="00:00:39.41" resultid="6271" heatid="9444" lane="4" entrytime="00:00:38.30" entrycourse="LCM" />
                <RESULT eventid="1561" points="207" reactiontime="+95" swimtime="00:03:25.81" resultid="6272" heatid="9492" lane="7" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:40.82" />
                    <SPLIT distance="150" swimtime="00:02:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="324" reactiontime="+87" swimtime="00:00:35.56" resultid="6273" heatid="9516" lane="1" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="5348" points="257" reactiontime="+77" swimtime="00:01:31.35" resultid="6274" heatid="9532" lane="3" entrytime="00:01:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="251" swimtime="00:01:27.90" resultid="6275" heatid="9571" lane="9" entrytime="00:01:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" athleteid="7532">
              <RESULTS>
                <RESULT eventid="1195" points="489" reactiontime="+78" swimtime="00:00:26.53" resultid="7533" heatid="9331" lane="9" entrytime="00:00:25.50" />
                <RESULT eventid="5331" points="521" reactiontime="+72" swimtime="00:00:27.87" resultid="7534" heatid="9528" lane="0" entrytime="00:00:26.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="6211">
              <RESULTS>
                <RESULT eventid="1229" points="257" reactiontime="+82" swimtime="00:02:59.30" resultid="6212" heatid="9345" lane="7" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:02:18.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="271" reactiontime="+78" swimtime="00:00:37.13" resultid="6213" heatid="9452" lane="5" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="324" swimtime="00:01:08.28" resultid="6214" heatid="9483" lane="6" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="282" reactiontime="+89" swimtime="00:00:34.20" resultid="6215" heatid="9522" lane="8" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="5399" points="270" reactiontime="+89" swimtime="00:02:37.72" resultid="6216" heatid="9554" lane="0" entrytime="00:02:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:57.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="211" reactiontime="+77" swimtime="00:03:07.70" resultid="6217" heatid="9587" lane="3" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                    <SPLIT distance="100" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:02:20.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-10" firstname="Sonia" gender="F" lastname="Bochyńska" nation="POL" license="503105600046" athleteid="6251">
              <RESULTS>
                <RESULT eventid="1133" points="562" reactiontime="+77" swimtime="00:00:28.67" resultid="6252" heatid="9315" lane="6" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1458" points="592" reactiontime="+70" swimtime="00:00:32.22" resultid="6253" heatid="9446" lane="4" entrytime="00:00:32.10" entrycourse="LCM" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="6254" heatid="9476" lane="8" entrytime="00:01:03.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="6242">
              <RESULTS>
                <RESULT eventid="1195" points="542" reactiontime="+72" swimtime="00:00:25.64" resultid="6243" heatid="9329" lane="1" entrytime="00:00:26.95" entrycourse="LCM" />
                <RESULT eventid="1229" points="447" reactiontime="+76" swimtime="00:02:29.07" resultid="6244" heatid="9347" lane="7" entrytime="00:02:38.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:53.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="460" reactiontime="+83" swimtime="00:00:31.12" resultid="6245" heatid="9453" lane="6" entrytime="00:00:35.80" entrycourse="LCM" />
                <RESULT eventid="1544" points="515" reactiontime="+70" swimtime="00:00:58.52" resultid="6246" heatid="9488" lane="8" entrytime="00:00:59.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="481" reactiontime="+72" swimtime="00:01:12.90" resultid="6247" heatid="9510" lane="4" entrytime="00:01:18.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="462" reactiontime="+78" swimtime="00:00:29.01" resultid="6248" heatid="9525" lane="6" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6249" heatid="9576" lane="8" entrytime="00:01:11.55" entrycourse="LCM" />
                <RESULT eventid="5585" points="495" reactiontime="+72" swimtime="00:00:32.79" resultid="6250" heatid="9603" lane="4" entrytime="00:00:33.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="6218">
              <RESULTS>
                <RESULT eventid="1133" points="359" reactiontime="+73" swimtime="00:00:33.30" resultid="6219" heatid="9313" lane="9" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1493" points="277" swimtime="00:03:33.30" resultid="6220" heatid="9460" lane="1" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                    <SPLIT distance="100" swimtime="00:01:42.97" />
                    <SPLIT distance="150" swimtime="00:02:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="353" reactiontime="+70" swimtime="00:01:30.69" resultid="6221" heatid="9503" lane="3" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="285" reactiontime="+72" swimtime="00:02:51.63" resultid="6222" heatid="9546" lane="8" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="364" reactiontime="+68" swimtime="00:00:41.16" resultid="6223" heatid="9595" lane="0" entrytime="00:00:40.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="6202">
              <RESULTS>
                <RESULT eventid="1195" points="112" reactiontime="+82" swimtime="00:00:43.26" resultid="6203" heatid="9319" lane="1" entrytime="00:00:42.08" entrycourse="LCM" />
                <RESULT eventid="1229" points="72" reactiontime="+86" swimtime="00:04:33.11" resultid="6204" heatid="9343" lane="0" entrytime="00:04:26.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.90" />
                    <SPLIT distance="100" swimtime="00:02:12.61" />
                    <SPLIT distance="150" swimtime="00:03:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="72" reactiontime="+90" swimtime="00:00:57.59" resultid="6205" heatid="9448" lane="5" entrytime="00:00:58.05" entrycourse="LCM" />
                <RESULT eventid="1544" points="117" reactiontime="+90" swimtime="00:01:35.80" resultid="6206" heatid="9478" lane="5" entrytime="00:01:36.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="69" reactiontime="+102" swimtime="00:02:06.35" resultid="6207" heatid="9535" lane="1" entrytime="00:02:12.27" entrycourse="LCM" />
                <RESULT eventid="5399" points="95" reactiontime="+98" swimtime="00:03:42.80" resultid="6208" heatid="9550" lane="8" entrytime="00:03:40.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                    <SPLIT distance="100" swimtime="00:01:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="64" reactiontime="+113" swimtime="00:04:38.96" resultid="6209" heatid="9584" lane="7" entrytime="00:04:47.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:03:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="91" reactiontime="+102" swimtime="00:08:08.40" resultid="6210" heatid="9619" lane="2" entrytime="00:07:57.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.58" />
                    <SPLIT distance="100" swimtime="00:01:54.81" />
                    <SPLIT distance="150" swimtime="00:03:00.29" />
                    <SPLIT distance="200" swimtime="00:04:03.97" />
                    <SPLIT distance="300" swimtime="00:06:11.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="6235">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="6236" heatid="9320" lane="3" entrytime="00:00:35.50" entrycourse="LCM" />
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="6237" heatid="9449" lane="5" entrytime="00:00:47.00" entrycourse="LCM" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6238" heatid="9480" lane="3" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="5331" status="DNS" swimtime="00:00:00.00" resultid="6239" heatid="9520" lane="6" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="5365" status="DNS" swimtime="00:00:00.00" resultid="6240" heatid="9536" lane="8" entrytime="00:01:40.00" entrycourse="LCM" />
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="6241" heatid="9573" lane="8" entrytime="00:01:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="6259">
              <RESULTS>
                <RESULT eventid="1510" points="157" reactiontime="+96" swimtime="00:03:54.31" resultid="6260" heatid="9463" lane="7" entrytime="00:03:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.79" />
                    <SPLIT distance="100" swimtime="00:01:53.99" />
                    <SPLIT distance="150" swimtime="00:02:55.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="181" reactiontime="+91" swimtime="00:01:40.82" resultid="6261" heatid="9507" lane="4" entrytime="00:01:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" status="DNS" swimtime="00:00:00.00" resultid="6262" heatid="9599" lane="4" entrytime="00:00:40.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105700035" athleteid="6401">
              <RESULTS>
                <RESULT eventid="1195" points="252" reactiontime="+105" swimtime="00:00:33.07" resultid="6402" heatid="9322" lane="7" entrytime="00:00:32.40" entrycourse="LCM" />
                <RESULT eventid="1476" points="105" reactiontime="+83" swimtime="00:00:50.88" resultid="6403" heatid="9450" lane="0" entrytime="00:00:46.00" entrycourse="LCM" />
                <RESULT eventid="1544" points="227" swimtime="00:01:16.81" resultid="6404" heatid="9482" lane="1" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="152" swimtime="00:01:46.94" resultid="6405" heatid="9507" lane="6" entrytime="00:01:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="197" reactiontime="+104" swimtime="00:00:44.53" resultid="6406" heatid="9598" lane="6" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1612" points="291" reactiontime="+60" swimtime="00:02:20.87" resultid="6281" heatid="9498" lane="3" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:46.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6263" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6259" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="6197" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="6401" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="5433" points="212" reactiontime="+84" swimtime="00:02:22.11" resultid="6282" heatid="9560" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.93" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6211" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="6224" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="6190" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="6259" number="4" reactiontime="+88" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1612" points="163" reactiontime="+79" swimtime="00:02:50.83" resultid="6283" heatid="9498" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:19.25" />
                    <SPLIT distance="150" swimtime="00:02:14.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6211" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="6190" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="6202" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="6224" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="5433" points="266" reactiontime="+92" swimtime="00:02:11.84" resultid="6284" heatid="9560" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:43.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6401" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="6202" number="2" reactiontime="+7" />
                    <RELAYPOSITION athleteid="6197" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="6263" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+75" swimtime="00:01:59.39" resultid="6276" heatid="9354" lane="5" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:02.15" />
                    <SPLIT distance="150" swimtime="00:01:32.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6251" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6228" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="6197" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="6242" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+80" swimtime="00:02:30.18" resultid="6280" heatid="9607" lane="6" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6211" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6190" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="6269" number="3" />
                    <RELAYPOSITION athleteid="6218" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1246" swimtime="00:02:12.92" resultid="6277" heatid="9354" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:40.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6269" number="1" />
                    <RELAYPOSITION athleteid="6224" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="6218" number="3" />
                    <RELAYPOSITION athleteid="6211" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WTM" nation="POL" clubid="7043" name="Wandzioch Team Maters">
          <ATHLETES>
            <ATHLETE birthdate="1992-12-08" firstname="Monika" gender="F" lastname="Matyszczyk" nation="POL" athleteid="7042">
              <RESULTS>
                <RESULT eventid="1458" points="136" reactiontime="+85" swimtime="00:00:52.57" resultid="7044" heatid="9441" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="5348" points="118" reactiontime="+76" swimtime="00:01:58.36" resultid="7045" heatid="9531" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-16" firstname="Krzysztof" gender="M" lastname="Wandzioch" nation="POL" athleteid="7046">
              <RESULTS>
                <RESULT eventid="1314" reactiontime="+75" status="OTL" swimtime="00:20:40.57" resultid="7047" heatid="9365" lane="2" entrytime="00:19:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:55.28" />
                    <SPLIT distance="200" swimtime="00:02:35.78" />
                    <SPLIT distance="250" swimtime="00:03:17.10" />
                    <SPLIT distance="300" swimtime="00:03:58.30" />
                    <SPLIT distance="350" swimtime="00:04:39.76" />
                    <SPLIT distance="400" swimtime="00:05:20.96" />
                    <SPLIT distance="450" swimtime="00:06:02.77" />
                    <SPLIT distance="500" swimtime="00:06:43.74" />
                    <SPLIT distance="550" swimtime="00:07:24.67" />
                    <SPLIT distance="600" swimtime="00:08:05.63" />
                    <SPLIT distance="650" swimtime="00:08:47.38" />
                    <SPLIT distance="700" swimtime="00:09:28.99" />
                    <SPLIT distance="750" swimtime="00:10:10.74" />
                    <SPLIT distance="800" swimtime="00:10:52.38" />
                    <SPLIT distance="850" swimtime="00:11:33.94" />
                    <SPLIT distance="900" swimtime="00:12:15.73" />
                    <SPLIT distance="950" swimtime="00:12:57.61" />
                    <SPLIT distance="1000" swimtime="00:13:39.89" />
                    <SPLIT distance="1050" swimtime="00:14:22.27" />
                    <SPLIT distance="1100" swimtime="00:15:04.50" />
                    <SPLIT distance="1150" swimtime="00:15:46.95" />
                    <SPLIT distance="1200" swimtime="00:16:29.00" />
                    <SPLIT distance="1250" swimtime="00:17:11.59" />
                    <SPLIT distance="1300" swimtime="00:17:53.36" />
                    <SPLIT distance="1350" swimtime="00:18:35.93" />
                    <SPLIT distance="1400" swimtime="00:19:17.89" />
                    <SPLIT distance="1450" swimtime="00:20:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="248" reactiontime="+81" swimtime="00:02:57.30" resultid="7048" heatid="9494" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="150" swimtime="00:02:12.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="312" reactiontime="+74" swimtime="00:05:59.35" resultid="7049" heatid="9566" lane="2" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:22.80" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                    <SPLIT distance="200" swimtime="00:02:54.98" />
                    <SPLIT distance="250" swimtime="00:03:49.16" />
                    <SPLIT distance="300" swimtime="00:04:42.21" />
                    <SPLIT distance="350" swimtime="00:05:21.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="7050" heatid="9574" lane="4" entrytime="00:01:22.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" clubid="7289" name="Warsaw Masters Team">
          <CONTACT email="agnieszka.z.mazurkiewicz@gmail.com" name="Mazurkiewicz" phone="882185766" street="Agnieszka" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="7428">
              <RESULTS>
                <RESULT eventid="1476" points="388" reactiontime="+68" swimtime="00:00:32.94" resultid="7430" heatid="9455" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="5331" points="428" reactiontime="+76" swimtime="00:00:29.76" resultid="7431" heatid="9526" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="5399" points="389" swimtime="00:02:19.64" resultid="7432" heatid="9556" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="7433" heatid="9577" lane="8" entrytime="00:01:06.00" />
                <RESULT eventid="1280" points="381" swimtime="00:10:23.38" resultid="9435" heatid="9359" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:51.18" />
                    <SPLIT distance="200" swimtime="00:02:30.80" />
                    <SPLIT distance="250" swimtime="00:03:10.10" />
                    <SPLIT distance="300" swimtime="00:03:49.80" />
                    <SPLIT distance="350" swimtime="00:04:29.28" />
                    <SPLIT distance="400" swimtime="00:05:09.07" />
                    <SPLIT distance="450" swimtime="00:05:48.05" />
                    <SPLIT distance="500" swimtime="00:06:28.45" />
                    <SPLIT distance="550" swimtime="00:07:08.93" />
                    <SPLIT distance="600" swimtime="00:07:48.63" />
                    <SPLIT distance="650" swimtime="00:08:27.59" />
                    <SPLIT distance="700" swimtime="00:09:07.05" />
                    <SPLIT distance="750" swimtime="00:09:45.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-13" firstname="Justyna" gender="F" lastname="Dąbrowska-Bień" nation="POL" athleteid="7402">
              <RESULTS>
                <RESULT eventid="1493" points="262" reactiontime="+81" swimtime="00:03:37.19" resultid="7403" heatid="9459" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:44.58" />
                    <SPLIT distance="150" swimtime="00:02:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="270" reactiontime="+77" swimtime="00:01:39.17" resultid="7404" heatid="9502" lane="4" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="303" reactiontime="+75" swimtime="00:00:43.76" resultid="7405" heatid="9594" lane="1" entrytime="00:00:44.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="7354">
              <RESULTS>
                <RESULT eventid="1493" points="346" swimtime="00:03:18.04" resultid="7355" heatid="9461" lane="9" entrytime="00:03:13.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:34.85" />
                    <SPLIT distance="150" swimtime="00:02:25.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="336" reactiontime="+71" swimtime="00:01:32.24" resultid="7356" heatid="9503" lane="4" entrytime="00:01:28.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="260" reactiontime="+72" swimtime="00:02:56.80" resultid="7357" heatid="9546" lane="0" entrytime="00:02:47.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:00:30.08" />
                    <SPLIT distance="150" swimtime="00:02:12.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="348" reactiontime="+78" swimtime="00:00:41.77" resultid="7358" heatid="9595" lane="8" entrytime="00:00:40.47" />
                <RESULT eventid="5619" points="246" swimtime="00:06:17.08" resultid="7359" heatid="9609" lane="9" entrytime="00:05:54.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:16.82" />
                    <SPLIT distance="200" swimtime="00:03:05.76" />
                    <SPLIT distance="250" swimtime="00:03:53.99" />
                    <SPLIT distance="300" swimtime="00:04:42.11" />
                    <SPLIT distance="350" swimtime="00:05:30.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-07" firstname="Daniel" gender="M" lastname="Julian Aguilar" nation="POL" athleteid="7319">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="7320" heatid="9329" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1476" status="DNS" swimtime="00:00:00.00" resultid="7322" heatid="9456" lane="9" entrytime="00:00:31.50" />
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="7323" heatid="9488" lane="7" entrytime="00:00:59.50" />
                <RESULT eventid="5399" status="DNS" swimtime="00:00:00.00" resultid="7324" heatid="9557" lane="8" entrytime="00:02:15.00" />
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="7325" heatid="9567" lane="9" entrytime="00:06:00.00" />
                <RESULT eventid="5551" status="DNS" swimtime="00:00:00.00" resultid="7326" heatid="9589" lane="7" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-10-11" firstname="Grzegorz" gender="M" lastname="Matyszewski" nation="POL" athleteid="7340">
              <RESULTS>
                <RESULT eventid="1195" points="254" reactiontime="+83" swimtime="00:00:33.01" resultid="7341" heatid="9321" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1510" points="262" reactiontime="+65" swimtime="00:03:17.94" resultid="7342" heatid="9465" lane="7" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:31.13" />
                    <SPLIT distance="150" swimtime="00:02:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="210" reactiontime="+63" swimtime="00:01:18.91" resultid="7343" heatid="9481" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="280" swimtime="00:01:27.24" resultid="7344" heatid="9509" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="167" reactiontime="+64" swimtime="00:03:04.90" resultid="7345" heatid="9551" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                    <SPLIT distance="150" swimtime="00:02:18.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="304" reactiontime="+69" swimtime="00:00:38.58" resultid="7346" heatid="9600" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="5636" points="162" swimtime="00:06:43.15" resultid="7347" heatid="9618" lane="9" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:22.25" />
                    <SPLIT distance="200" swimtime="00:03:14.58" />
                    <SPLIT distance="250" swimtime="00:04:07.67" />
                    <SPLIT distance="300" swimtime="00:05:01.21" />
                    <SPLIT distance="350" swimtime="00:05:54.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="7411">
              <RESULTS>
                <RESULT eventid="1229" points="358" reactiontime="+79" swimtime="00:02:40.50" resultid="7412" heatid="9346" lane="5" entrytime="00:02:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:02:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="406" reactiontime="+77" swimtime="00:01:03.34" resultid="7414" heatid="9486" lane="0" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="417" reactiontime="+57" swimtime="00:02:16.45" resultid="7415" heatid="9556" lane="7" entrytime="00:02:18.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="411" swimtime="00:04:55.89" resultid="7416" heatid="9614" lane="1" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                    <SPLIT distance="150" swimtime="00:01:46.38" />
                    <SPLIT distance="200" swimtime="00:02:24.48" />
                    <SPLIT distance="250" swimtime="00:03:02.19" />
                    <SPLIT distance="300" swimtime="00:03:40.69" />
                    <SPLIT distance="350" swimtime="00:04:18.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="7422">
              <RESULTS>
                <RESULT eventid="1229" points="370" reactiontime="+93" swimtime="00:02:38.75" resultid="7423" heatid="9347" lane="3" entrytime="00:02:37.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:02.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="302" reactiontime="+104" swimtime="00:21:37.57" resultid="7424" heatid="9366" lane="4" entrytime="00:21:28.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                    <SPLIT distance="200" swimtime="00:02:47.85" />
                    <SPLIT distance="250" swimtime="00:03:32.16" />
                    <SPLIT distance="300" swimtime="00:04:15.54" />
                    <SPLIT distance="350" swimtime="00:04:59.51" />
                    <SPLIT distance="400" swimtime="00:05:42.40" />
                    <SPLIT distance="450" swimtime="00:06:26.81" />
                    <SPLIT distance="500" swimtime="00:07:09.82" />
                    <SPLIT distance="550" swimtime="00:07:53.11" />
                    <SPLIT distance="600" swimtime="00:08:36.03" />
                    <SPLIT distance="650" swimtime="00:09:19.07" />
                    <SPLIT distance="700" swimtime="00:10:01.89" />
                    <SPLIT distance="750" swimtime="00:10:45.56" />
                    <SPLIT distance="800" swimtime="00:11:28.58" />
                    <SPLIT distance="850" swimtime="00:12:12.31" />
                    <SPLIT distance="900" swimtime="00:12:55.55" />
                    <SPLIT distance="950" swimtime="00:13:40.19" />
                    <SPLIT distance="1000" swimtime="00:14:23.74" />
                    <SPLIT distance="1050" swimtime="00:15:08.03" />
                    <SPLIT distance="1100" swimtime="00:15:51.30" />
                    <SPLIT distance="1150" swimtime="00:16:36.04" />
                    <SPLIT distance="1200" swimtime="00:17:20.06" />
                    <SPLIT distance="1250" swimtime="00:18:04.22" />
                    <SPLIT distance="1300" swimtime="00:18:47.80" />
                    <SPLIT distance="1350" swimtime="00:19:31.97" />
                    <SPLIT distance="1400" swimtime="00:20:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="390" swimtime="00:02:53.27" resultid="7425" heatid="9467" lane="6" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="150" swimtime="00:02:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="290" reactiontime="+92" swimtime="00:02:48.34" resultid="7426" heatid="9495" lane="2" entrytime="00:02:49.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="150" swimtime="00:02:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" status="DNS" swimtime="00:00:00.00" resultid="7427" heatid="9567" lane="2" entrytime="00:05:42.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="7290">
              <RESULTS>
                <RESULT eventid="1212" points="218" reactiontime="+92" swimtime="00:03:29.24" resultid="7291" heatid="9338" lane="5" entrytime="00:03:20.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:43.93" />
                    <SPLIT distance="150" swimtime="00:02:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="201" reactiontime="+93" swimtime="00:13:46.48" resultid="7292" heatid="9356" lane="7" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                    <SPLIT distance="150" swimtime="00:02:26.59" />
                    <SPLIT distance="200" swimtime="00:03:18.35" />
                    <SPLIT distance="250" swimtime="00:04:10.38" />
                    <SPLIT distance="300" swimtime="00:05:02.53" />
                    <SPLIT distance="350" swimtime="00:05:55.14" />
                    <SPLIT distance="400" swimtime="00:06:47.84" />
                    <SPLIT distance="450" swimtime="00:07:39.89" />
                    <SPLIT distance="500" swimtime="00:08:32.18" />
                    <SPLIT distance="550" swimtime="00:09:25.06" />
                    <SPLIT distance="600" swimtime="00:10:17.89" />
                    <SPLIT distance="650" swimtime="00:11:10.95" />
                    <SPLIT distance="700" swimtime="00:12:04.29" />
                    <SPLIT distance="750" swimtime="00:12:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="267" reactiontime="+84" swimtime="00:03:35.89" resultid="7293" heatid="9460" lane="2" entrytime="00:03:26.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                    <SPLIT distance="100" swimtime="00:01:44.39" />
                    <SPLIT distance="150" swimtime="00:02:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1527" points="216" reactiontime="+95" swimtime="00:01:26.12" resultid="7294" heatid="9471" lane="5" entrytime="00:01:26.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="270" swimtime="00:01:39.15" resultid="7295" heatid="9503" lane="1" entrytime="00:01:33.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="226" reactiontime="+92" swimtime="00:03:05.35" resultid="7296" heatid="9544" lane="5" entrytime="00:03:02.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:30.68" />
                    <SPLIT distance="150" swimtime="00:02:19.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="7360">
              <RESULTS>
                <RESULT eventid="1195" points="420" reactiontime="+76" swimtime="00:00:27.91" resultid="7361" heatid="9327" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1229" points="409" reactiontime="+70" swimtime="00:02:33.48" resultid="7362" heatid="9348" lane="8" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="480" reactiontime="+67" swimtime="00:02:41.68" resultid="7363" heatid="9468" lane="2" entrytime="00:02:39.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="443" swimtime="00:01:14.91" resultid="7364" heatid="9512" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="483" reactiontime="+79" swimtime="00:00:33.07" resultid="7365" heatid="9603" lane="5" entrytime="00:00:33.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="7303">
              <RESULTS>
                <RESULT eventid="1133" points="424" reactiontime="+64" swimtime="00:00:31.49" resultid="7304" heatid="9313" lane="4" entrytime="00:00:31.84" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="7305" heatid="9460" lane="7" entrytime="00:03:29.07" />
                <RESULT eventid="1527" status="DNS" swimtime="00:00:00.00" resultid="7306" heatid="9473" lane="0" entrytime="00:01:18.00" />
                <RESULT eventid="5279" points="360" swimtime="00:01:30.12" resultid="7307" heatid="9503" lane="6" entrytime="00:01:31.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="400" reactiontime="+67" swimtime="00:00:39.88" resultid="7308" heatid="9595" lane="7" entrytime="00:00:40.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="7388">
              <RESULTS>
                <RESULT eventid="1195" points="157" reactiontime="+99" swimtime="00:00:38.71" resultid="7389" heatid="9319" lane="4" entrytime="00:00:39.10" />
                <RESULT eventid="1280" points="167" reactiontime="+101" swimtime="00:13:40.03" resultid="7390" heatid="9362" lane="5" entrytime="00:13:33.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                    <SPLIT distance="100" swimtime="00:03:21.16" />
                    <SPLIT distance="150" swimtime="00:02:28.03" />
                    <SPLIT distance="250" swimtime="00:04:14.31" />
                    <SPLIT distance="300" swimtime="00:05:06.41" />
                    <SPLIT distance="350" swimtime="00:05:59.30" />
                    <SPLIT distance="400" swimtime="00:06:51.32" />
                    <SPLIT distance="450" swimtime="00:07:43.71" />
                    <SPLIT distance="500" swimtime="00:10:19.96" />
                    <SPLIT distance="550" swimtime="00:09:28.53" />
                    <SPLIT distance="600" swimtime="00:13:40.11" />
                    <SPLIT distance="650" swimtime="00:12:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="73" reactiontime="+93" swimtime="00:00:57.48" resultid="7391" heatid="9449" lane="2" entrytime="00:00:51.20" />
                <RESULT eventid="1544" points="156" swimtime="00:01:27.05" resultid="7392" heatid="9480" lane="9" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="92" reactiontime="+108" swimtime="00:00:49.63" resultid="7393" heatid="9519" lane="6" entrytime="00:00:46.76" />
                <RESULT eventid="5399" points="152" reactiontime="+108" swimtime="00:03:10.97" resultid="7394" heatid="9551" lane="8" entrytime="00:03:05.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:32.78" />
                    <SPLIT distance="150" swimtime="00:02:22.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="166" reactiontime="+103" swimtime="00:06:39.95" resultid="7395" heatid="9618" lane="3" entrytime="00:06:41.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:36.53" />
                    <SPLIT distance="150" swimtime="00:02:27.42" />
                    <SPLIT distance="200" swimtime="00:03:19.23" />
                    <SPLIT distance="250" swimtime="00:04:11.23" />
                    <SPLIT distance="300" swimtime="00:05:02.55" />
                    <SPLIT distance="350" swimtime="00:05:52.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="7297">
              <RESULTS>
                <RESULT eventid="1229" points="362" reactiontime="+82" swimtime="00:02:39.88" resultid="7298" heatid="9347" lane="0" entrytime="00:02:39.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:02:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="366" reactiontime="+85" swimtime="00:10:31.67" resultid="7299" heatid="9359" lane="0" entrytime="00:10:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:51.47" />
                    <SPLIT distance="200" swimtime="00:02:31.29" />
                    <SPLIT distance="250" swimtime="00:03:11.08" />
                    <SPLIT distance="300" swimtime="00:03:51.12" />
                    <SPLIT distance="350" swimtime="00:04:31.31" />
                    <SPLIT distance="400" swimtime="00:05:11.95" />
                    <SPLIT distance="450" swimtime="00:05:53.12" />
                    <SPLIT distance="500" swimtime="00:06:33.29" />
                    <SPLIT distance="550" swimtime="00:07:13.57" />
                    <SPLIT distance="600" swimtime="00:07:54.19" />
                    <SPLIT distance="650" swimtime="00:08:34.46" />
                    <SPLIT distance="700" swimtime="00:09:15.06" />
                    <SPLIT distance="750" swimtime="00:09:54.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="404" reactiontime="+81" swimtime="00:01:03.45" resultid="7300" heatid="9486" lane="2" entrytime="00:01:02.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="392" reactiontime="+89" swimtime="00:02:19.35" resultid="7301" heatid="9556" lane="3" entrytime="00:02:17.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="397" reactiontime="+83" swimtime="00:04:59.22" resultid="7302" heatid="9614" lane="8" entrytime="00:05:00.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:49.33" />
                    <SPLIT distance="200" swimtime="00:02:28.24" />
                    <SPLIT distance="250" swimtime="00:03:07.29" />
                    <SPLIT distance="300" swimtime="00:03:45.84" />
                    <SPLIT distance="350" swimtime="00:04:23.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="7309">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1527" points="590" reactiontime="+71" swimtime="00:01:01.63" resultid="7310" heatid="9476" lane="7" entrytime="00:01:02.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="496" reactiontime="+75" swimtime="00:00:30.85" resultid="7311" heatid="9517" lane="3" entrytime="00:00:30.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5499" points="546" reactiontime="+74" swimtime="00:01:07.84" resultid="7312" heatid="9571" lane="4" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="578" reactiontime="+76" swimtime="00:00:35.28" resultid="7313" heatid="9596" lane="3" entrytime="00:00:35.81" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-23" firstname="Wojciech" gender="M" lastname="Janicki" nation="POL" athleteid="7314">
              <RESULTS>
                <RESULT eventid="1195" points="430" reactiontime="+75" swimtime="00:00:27.69" resultid="7315" heatid="9330" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1229" points="321" reactiontime="+75" swimtime="00:02:46.37" resultid="7316" heatid="9347" lane="8" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="450" swimtime="00:01:01.19" resultid="7317" heatid="9488" lane="1" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="467" reactiontime="+74" swimtime="00:00:28.91" resultid="7318" heatid="9527" lane="0" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="7334">
              <RESULTS>
                <RESULT eventid="1527" points="307" reactiontime="+72" swimtime="00:01:16.61" resultid="7335" heatid="9473" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="299" reactiontime="+86" swimtime="00:00:36.51" resultid="7336" heatid="9516" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="5382" points="324" reactiontime="+79" swimtime="00:02:44.48" resultid="7337" heatid="9545" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:02.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5499" points="248" reactiontime="+85" swimtime="00:01:28.22" resultid="7338" heatid="9570" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="299" reactiontime="+78" swimtime="00:05:53.47" resultid="7339" heatid="9610" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:05.18" />
                    <SPLIT distance="200" swimtime="00:02:51.15" />
                    <SPLIT distance="250" swimtime="00:03:36.93" />
                    <SPLIT distance="300" swimtime="00:04:23.29" />
                    <SPLIT distance="350" swimtime="00:05:09.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="277" reactiontime="+83" swimtime="00:12:23.26" resultid="9034" heatid="9356" lane="5" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                    <SPLIT distance="200" swimtime="00:02:57.07" />
                    <SPLIT distance="250" swimtime="00:03:43.52" />
                    <SPLIT distance="300" swimtime="00:04:30.77" />
                    <SPLIT distance="350" swimtime="00:05:17.74" />
                    <SPLIT distance="400" swimtime="00:06:04.89" />
                    <SPLIT distance="450" swimtime="00:06:52.42" />
                    <SPLIT distance="500" swimtime="00:07:40.63" />
                    <SPLIT distance="550" swimtime="00:08:28.16" />
                    <SPLIT distance="600" swimtime="00:09:16.82" />
                    <SPLIT distance="650" swimtime="00:10:04.82" />
                    <SPLIT distance="700" swimtime="00:10:51.55" />
                    <SPLIT distance="750" swimtime="00:11:38.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="7348">
              <RESULTS>
                <RESULT eventid="1229" points="207" swimtime="00:03:12.66" resultid="7349" heatid="9344" lane="6" entrytime="00:03:11.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="150" swimtime="00:02:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="240" reactiontime="+79" swimtime="00:03:23.83" resultid="7350" heatid="9465" lane="0" entrytime="00:03:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="265" reactiontime="+70" swimtime="00:01:28.93" resultid="7351" heatid="9509" lane="2" entrytime="00:01:27.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5467" points="173" swimtime="00:07:17.54" resultid="7352" heatid="9565" lane="6" entrytime="00:07:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.29" />
                    <SPLIT distance="100" swimtime="00:01:52.26" />
                    <SPLIT distance="150" swimtime="00:02:52.40" />
                    <SPLIT distance="200" swimtime="00:03:48.59" />
                    <SPLIT distance="250" swimtime="00:04:44.86" />
                    <SPLIT distance="300" swimtime="00:05:42.26" />
                    <SPLIT distance="350" swimtime="00:06:31.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="310" reactiontime="+82" swimtime="00:00:38.31" resultid="7353" heatid="9601" lane="4" entrytime="00:00:37.52" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="7434">
              <RESULTS>
                <RESULT eventid="1195" points="394" reactiontime="+75" swimtime="00:00:28.51" resultid="7435" heatid="9324" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1280" points="332" swimtime="00:10:52.37" resultid="7436" heatid="9359" lane="9" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:54.54" />
                    <SPLIT distance="200" swimtime="00:02:35.02" />
                    <SPLIT distance="250" swimtime="00:03:15.52" />
                    <SPLIT distance="300" swimtime="00:03:55.69" />
                    <SPLIT distance="350" swimtime="00:04:36.12" />
                    <SPLIT distance="400" swimtime="00:05:16.89" />
                    <SPLIT distance="450" swimtime="00:05:58.27" />
                    <SPLIT distance="500" swimtime="00:06:40.51" />
                    <SPLIT distance="550" swimtime="00:07:22.96" />
                    <SPLIT distance="600" swimtime="00:08:05.47" />
                    <SPLIT distance="650" swimtime="00:08:47.83" />
                    <SPLIT distance="700" swimtime="00:09:30.98" />
                    <SPLIT distance="750" swimtime="00:10:13.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="394" reactiontime="+72" swimtime="00:01:03.94" resultid="7437" heatid="9485" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="379" reactiontime="+71" swimtime="00:02:20.84" resultid="7438" heatid="9555" lane="5" entrytime="00:02:20.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="150" swimtime="00:01:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="362" reactiontime="+71" swimtime="00:05:08.67" resultid="7439" heatid="9615" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:52.23" />
                    <SPLIT distance="200" swimtime="00:02:31.85" />
                    <SPLIT distance="250" swimtime="00:03:11.87" />
                    <SPLIT distance="300" swimtime="00:03:52.34" />
                    <SPLIT distance="350" swimtime="00:04:31.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="7372">
              <RESULTS>
                <RESULT eventid="1510" points="214" swimtime="00:03:31.65" resultid="7373" heatid="9464" lane="6" entrytime="00:03:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                    <SPLIT distance="100" swimtime="00:01:40.11" />
                    <SPLIT distance="150" swimtime="00:02:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="112" reactiontime="+99" swimtime="00:03:51.17" resultid="7374" heatid="9494" lane="8" entrytime="00:03:45.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:44.37" />
                    <SPLIT distance="150" swimtime="00:02:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="211" reactiontime="+98" swimtime="00:01:35.94" resultid="7375" heatid="9508" lane="8" entrytime="00:01:34.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="150" reactiontime="+101" swimtime="00:03:11.88" resultid="7376" heatid="9548" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="142" reactiontime="+101" swimtime="00:01:35.48" resultid="7377" heatid="9573" lane="2" entrytime="00:01:36.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="219" reactiontime="+107" swimtime="00:00:43.05" resultid="7378" heatid="9599" lane="3" entrytime="00:00:41.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="7400">
              <RESULTS>
                <RESULT eventid="1195" points="521" reactiontime="+79" swimtime="00:00:25.98" resultid="7401" heatid="9331" lane="6" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="7417">
              <RESULTS>
                <RESULT eventid="1510" points="177" swimtime="00:03:45.23" resultid="7418" heatid="9463" lane="6" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.19" />
                    <SPLIT distance="100" swimtime="00:01:46.92" />
                    <SPLIT distance="150" swimtime="00:02:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="187" reactiontime="+99" swimtime="00:01:21.99" resultid="7419" heatid="9479" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="178" reactiontime="+108" swimtime="00:01:41.54" resultid="7420" heatid="9506" lane="7" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="129" reactiontime="+104" swimtime="00:00:44.35" resultid="7421" heatid="9518" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="7406">
              <RESULTS>
                <RESULT eventid="1212" points="335" swimtime="00:03:01.57" resultid="7407" heatid="9337" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:23.86" />
                    <SPLIT distance="150" swimtime="00:02:18.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="331" reactiontime="+74" swimtime="00:11:40.28" resultid="7408" heatid="9355" lane="8" entrytime="00:11:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                    <SPLIT distance="200" swimtime="00:02:48.30" />
                    <SPLIT distance="250" swimtime="00:03:32.72" />
                    <SPLIT distance="300" swimtime="00:04:16.68" />
                    <SPLIT distance="350" swimtime="00:05:01.39" />
                    <SPLIT distance="400" swimtime="00:05:45.80" />
                    <SPLIT distance="450" swimtime="00:06:30.63" />
                    <SPLIT distance="500" swimtime="00:07:15.52" />
                    <SPLIT distance="550" swimtime="00:08:00.16" />
                    <SPLIT distance="600" swimtime="00:08:44.96" />
                    <SPLIT distance="650" swimtime="00:09:29.67" />
                    <SPLIT distance="700" swimtime="00:10:14.14" />
                    <SPLIT distance="750" swimtime="00:10:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5314" points="372" reactiontime="+84" swimtime="00:00:33.94" resultid="7409" heatid="9516" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="5450" status="DNS" swimtime="00:00:00.00" resultid="7410" heatid="9562" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="7328">
              <RESULTS>
                <RESULT eventid="1195" points="361" reactiontime="+81" swimtime="00:00:29.35" resultid="7329" heatid="9324" lane="5" entrytime="00:00:29.56" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1544" points="370" reactiontime="+83" swimtime="00:01:05.29" resultid="7330" heatid="9482" lane="3" entrytime="00:01:09.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5365" points="318" reactiontime="+73" swimtime="00:01:15.91" resultid="7331" heatid="9534" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5399" points="338" swimtime="00:02:26.40" resultid="7332" heatid="9555" lane="9" entrytime="00:02:28.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5551" points="312" reactiontime="+72" swimtime="00:02:44.88" resultid="7333" heatid="9588" lane="8" entrytime="00:02:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="150" swimtime="00:02:02.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="7379">
              <RESULTS>
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="7380" heatid="9326" lane="5" entrytime="00:00:28.65" />
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="7381" heatid="9347" lane="6" entrytime="00:02:38.00" />
                <RESULT eventid="1476" points="381" reactiontime="+78" swimtime="00:00:33.15" resultid="7382" heatid="9455" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1544" points="455" swimtime="00:01:00.98" resultid="7383" heatid="9486" lane="6" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="423" reactiontime="+78" swimtime="00:00:29.86" resultid="7384" heatid="9523" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="5365" points="400" reactiontime="+72" swimtime="00:01:10.35" resultid="7385" heatid="9539" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="379" reactiontime="+82" swimtime="00:01:08.82" resultid="7386" heatid="9575" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="372" reactiontime="+74" swimtime="00:02:35.50" resultid="7387" heatid="9589" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:55.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="7366">
              <RESULTS>
                <RESULT eventid="1195" points="439" reactiontime="+77" swimtime="00:00:27.50" resultid="7367" heatid="9329" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="1544" points="589" reactiontime="+70" swimtime="00:00:55.95" resultid="7368" heatid="9490" lane="0" entrytime="00:00:55.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="558" reactiontime="+75" swimtime="00:00:27.23" resultid="7369" heatid="9528" lane="8" entrytime="00:00:26.57" />
                <RESULT eventid="5399" points="489" reactiontime="+78" swimtime="00:02:09.43" resultid="7370" heatid="9557" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                    <SPLIT distance="150" swimtime="00:01:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" status="DNS" swimtime="00:00:00.00" resultid="7371" heatid="9578" lane="0" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="7396">
              <RESULTS>
                <RESULT eventid="1297" points="92" swimtime="00:34:09.93" resultid="7397" heatid="9364" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.94" />
                    <SPLIT distance="100" swimtime="00:02:10.98" />
                    <SPLIT distance="150" swimtime="00:03:20.94" />
                    <SPLIT distance="200" swimtime="00:04:30.97" />
                    <SPLIT distance="250" swimtime="00:05:41.45" />
                    <SPLIT distance="300" swimtime="00:06:51.92" />
                    <SPLIT distance="350" swimtime="00:08:00.65" />
                    <SPLIT distance="400" swimtime="00:09:08.93" />
                    <SPLIT distance="450" swimtime="00:10:17.46" />
                    <SPLIT distance="500" swimtime="00:11:29.11" />
                    <SPLIT distance="550" swimtime="00:12:37.85" />
                    <SPLIT distance="600" swimtime="00:13:46.38" />
                    <SPLIT distance="650" swimtime="00:14:55.07" />
                    <SPLIT distance="700" swimtime="00:16:04.08" />
                    <SPLIT distance="750" swimtime="00:17:12.34" />
                    <SPLIT distance="800" swimtime="00:18:20.93" />
                    <SPLIT distance="850" swimtime="00:19:28.61" />
                    <SPLIT distance="900" swimtime="00:20:37.76" />
                    <SPLIT distance="950" swimtime="00:21:46.15" />
                    <SPLIT distance="1000" swimtime="00:22:53.78" />
                    <SPLIT distance="1050" swimtime="00:24:01.72" />
                    <SPLIT distance="1100" swimtime="00:25:10.00" />
                    <SPLIT distance="1150" swimtime="00:26:18.29" />
                    <SPLIT distance="1200" swimtime="00:27:26.10" />
                    <SPLIT distance="1250" swimtime="00:28:33.41" />
                    <SPLIT distance="1300" swimtime="00:29:40.34" />
                    <SPLIT distance="1350" swimtime="00:30:48.61" />
                    <SPLIT distance="1400" swimtime="00:31:56.60" />
                    <SPLIT distance="1450" swimtime="00:33:04.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="76" swimtime="00:04:26.02" resultid="7398" heatid="9542" lane="3" entrytime="00:04:16.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.88" />
                    <SPLIT distance="100" swimtime="00:02:07.99" />
                    <SPLIT distance="150" swimtime="00:03:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="82" swimtime="00:09:04.08" resultid="7399" heatid="9612" lane="6" entrytime="00:08:32.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.84" />
                    <SPLIT distance="100" swimtime="00:02:10.36" />
                    <SPLIT distance="150" swimtime="00:03:20.03" />
                    <SPLIT distance="200" swimtime="00:04:30.46" />
                    <SPLIT distance="250" swimtime="00:05:40.83" />
                    <SPLIT distance="300" swimtime="00:06:50.47" />
                    <SPLIT distance="350" swimtime="00:07:58.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WMT 2" number="2">
              <RESULTS>
                <RESULT eventid="5433" points="476" reactiontime="+74" swimtime="00:01:48.60" resultid="7441" heatid="9561" lane="5" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="100" swimtime="00:00:52.92" />
                    <SPLIT distance="150" swimtime="00:01:20.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7366" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="7314" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="7319" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7379" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WMT 4" number="4">
              <RESULTS>
                <RESULT eventid="1612" points="395" reactiontime="+72" swimtime="00:02:07.27" resultid="7443" heatid="9499" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:06.05" />
                    <SPLIT distance="150" swimtime="00:01:34.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7428" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="7360" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="7314" number="3" />
                    <RELAYPOSITION athleteid="7319" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WMT 5" number="5">
              <RESULTS>
                <RESULT eventid="1612" points="376" reactiontime="+68" swimtime="00:02:09.39" resultid="7444" heatid="9499" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:40.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7379" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="7297" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="7434" number="3" />
                    <RELAYPOSITION athleteid="7411" number="4" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WMT 1" number="1">
              <RESULTS>
                <RESULT eventid="1246" reactiontime="+71" swimtime="00:02:05.92" resultid="7440" heatid="9354" lane="0" entrytime="00:02:04.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                    <SPLIT distance="150" swimtime="00:01:35.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7400" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="7303" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="7290" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="7328" number="4" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WMT 3" number="3">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+65" swimtime="00:02:14.71" resultid="7442" heatid="9607" lane="1" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:43.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7319" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="7348" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="7309" number="3" />
                    <RELAYPOSITION athleteid="7303" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WZ" nation="POL" clubid="6874" name="Weteran Zabrze">
          <CONTACT city="Zabrze" name="Bosowski Włodzimierz" street="Św. Jana" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="102611600018" athleteid="6905">
              <RESULTS>
                <RESULT eventid="1510" points="172" reactiontime="+84" swimtime="00:03:47.39" resultid="6906" heatid="9463" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                    <SPLIT distance="100" swimtime="00:01:50.25" />
                    <SPLIT distance="150" swimtime="00:02:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="161" reactiontime="+104" swimtime="00:01:44.93" resultid="6907" heatid="9507" lane="8" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="168" reactiontime="+113" swimtime="00:00:47.02" resultid="6908" heatid="9598" lane="7" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="102611600022" athleteid="6915">
              <RESULTS>
                <RESULT eventid="1195" points="154" reactiontime="+107" swimtime="00:00:38.93" resultid="6916" heatid="9319" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1544" points="151" reactiontime="+107" swimtime="00:01:28.08" resultid="6917" heatid="9479" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="127" swimtime="00:03:22.58" resultid="6918" heatid="9550" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:37.35" />
                    <SPLIT distance="150" swimtime="00:02:31.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-20" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="102611600015" athleteid="6961">
              <RESULTS>
                <RESULT eventid="1195" points="245" reactiontime="+91" swimtime="00:00:33.41" resultid="6962" heatid="9321" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1476" points="104" reactiontime="+87" swimtime="00:00:51.11" resultid="6963" heatid="9450" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1544" points="187" reactiontime="+79" swimtime="00:01:21.94" resultid="6964" heatid="9480" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="169" reactiontime="+84" swimtime="00:00:40.56" resultid="6965" heatid="9521" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="102611600017" athleteid="6900">
              <RESULTS>
                <RESULT eventid="1133" points="172" reactiontime="+100" swimtime="00:00:42.54" resultid="6901" heatid="9310" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1527" points="144" reactiontime="+94" swimtime="00:01:38.45" resultid="6902" heatid="9471" lane="0" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" reactiontime="+96" status="DNF" swimtime="00:00:00.00" resultid="6903" heatid="9543" lane="8" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="6904" heatid="9579" lane="3" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="102611600023" athleteid="6919">
              <RESULTS>
                <RESULT eventid="1133" points="222" reactiontime="+83" swimtime="00:00:39.06" resultid="6920" heatid="9310" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1458" points="183" reactiontime="+80" swimtime="00:00:47.61" resultid="6921" heatid="9442" lane="8" entrytime="00:00:49.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1527" points="195" swimtime="00:01:29.04" resultid="6922" heatid="9471" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5348" points="161" reactiontime="+68" swimtime="00:01:46.70" resultid="6923" heatid="9530" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5534" points="152" reactiontime="+73" swimtime="00:03:51.99" resultid="6924" heatid="9580" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:01:53.49" />
                    <SPLIT distance="150" swimtime="00:02:54.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611100004" athleteid="6875">
              <RESULTS>
                <RESULT eventid="1476" points="170" reactiontime="+73" swimtime="00:00:43.35" resultid="6876" heatid="9450" lane="3" entrytime="00:00:44.11" />
                <RESULT eventid="5365" points="141" reactiontime="+73" swimtime="00:01:39.40" resultid="6877" heatid="9536" lane="0" entrytime="00:01:41.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="129" reactiontime="+72" swimtime="00:03:41.13" resultid="6878" heatid="9585" lane="1" entrytime="00:03:49.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                    <SPLIT distance="100" swimtime="00:01:43.93" />
                    <SPLIT distance="150" swimtime="00:02:43.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-27" firstname="Danuta" gender="F" lastname="Skorupa" nation="POL" license="102611600020" athleteid="6897">
              <RESULTS>
                <RESULT eventid="1458" points="48" reactiontime="+102" swimtime="00:01:14.35" resultid="6898" heatid="9441" lane="7" entrytime="00:00:59.50" />
                <RESULT eventid="5568" points="39" swimtime="00:01:26.55" resultid="6899" heatid="9591" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="102611600016" athleteid="6925">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1263" points="462" swimtime="00:10:27.00" resultid="6926" heatid="9355" lane="6" entrytime="00:10:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:54.62" />
                    <SPLIT distance="200" swimtime="00:02:34.23" />
                    <SPLIT distance="250" swimtime="00:03:14.00" />
                    <SPLIT distance="300" swimtime="00:03:53.57" />
                    <SPLIT distance="350" swimtime="00:04:33.27" />
                    <SPLIT distance="400" swimtime="00:05:12.70" />
                    <SPLIT distance="450" swimtime="00:05:52.35" />
                    <SPLIT distance="500" swimtime="00:06:31.69" />
                    <SPLIT distance="550" swimtime="00:07:11.44" />
                    <SPLIT distance="600" swimtime="00:07:50.76" />
                    <SPLIT distance="650" swimtime="00:08:30.36" />
                    <SPLIT distance="700" swimtime="00:09:09.65" />
                    <SPLIT distance="750" swimtime="00:09:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1493" points="423" swimtime="00:03:05.28" resultid="6927" heatid="9461" lane="1" entrytime="00:03:06.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5279" points="415" swimtime="00:01:25.91" resultid="6928" heatid="9504" lane="7" entrytime="00:01:24.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="449" reactiontime="+87" swimtime="00:02:27.47" resultid="6929" heatid="9547" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5568" points="411" reactiontime="+72" swimtime="00:00:39.53" resultid="6930" heatid="9595" lane="1" entrytime="00:00:40.05" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5619" points="456" swimtime="00:05:07.02" resultid="6931" heatid="9609" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                    <SPLIT distance="200" swimtime="00:02:32.39" />
                    <SPLIT distance="250" swimtime="00:03:11.76" />
                    <SPLIT distance="300" swimtime="00:03:50.74" />
                    <SPLIT distance="350" swimtime="00:04:29.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="102611600021" athleteid="6892">
              <RESULTS>
                <RESULT eventid="1476" points="207" reactiontime="+77" swimtime="00:00:40.61" resultid="6893" heatid="9451" lane="5" entrytime="00:00:40.24" />
                <RESULT eventid="1544" points="280" swimtime="00:01:11.67" resultid="6894" heatid="9482" lane="9" entrytime="00:01:12.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5365" points="200" reactiontime="+79" swimtime="00:01:28.56" resultid="6895" heatid="9537" lane="5" entrytime="00:01:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5551" points="187" reactiontime="+80" swimtime="00:03:15.64" resultid="6896" heatid="9586" lane="2" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="100" swimtime="00:01:35.17" />
                    <SPLIT distance="150" swimtime="00:02:25.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="102611600014" athleteid="6957">
              <RESULTS>
                <RESULT eventid="1195" points="107" reactiontime="+104" swimtime="00:00:43.91" resultid="6958" heatid="9319" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1476" points="66" reactiontime="+103" swimtime="00:00:59.34" resultid="6959" heatid="9449" lane="9" entrytime="00:00:58.00" />
                <RESULT eventid="5331" points="57" reactiontime="+111" swimtime="00:00:58.14" resultid="6960" heatid="9519" lane="2" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="102611600019" athleteid="6909">
              <RESULTS>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="1493" points="151" reactiontime="+93" swimtime="00:04:20.84" resultid="6910" heatid="9459" lane="0" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.88" />
                    <SPLIT distance="100" swimtime="00:02:04.13" />
                    <SPLIT distance="150" swimtime="00:03:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5279" points="168" swimtime="00:01:56.18" resultid="6911" heatid="9501" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5314" points="104" reactiontime="+93" swimtime="00:00:51.88" resultid="6912" heatid="9514" lane="6" entrytime="00:00:52.00" />
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5499" points="103" reactiontime="+93" swimtime="00:01:58.31" resultid="6913" heatid="9570" lane="0" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas lepszy od Rekordu Polski" eventid="5568" points="160" reactiontime="+93" swimtime="00:00:54.14" resultid="6914" heatid="9593" lane="0" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="102611600024" athleteid="6888">
              <RESULTS>
                <RESULT eventid="1133" points="110" reactiontime="+92" swimtime="00:00:49.39" resultid="6889" heatid="9309" lane="3" entrytime="00:00:49.50" />
                <RESULT eventid="1458" points="95" reactiontime="+81" swimtime="00:00:59.25" resultid="6890" heatid="9441" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="5568" points="127" reactiontime="+80" swimtime="00:00:58.36" resultid="6891" heatid="9592" lane="4" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1612" points="134" reactiontime="+76" swimtime="00:03:02.15" resultid="6939" heatid="9498" lane="7" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:34.53" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6875" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6905" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="6961" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="6957" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="5433" points="145" swimtime="00:02:41.49" resultid="6941" heatid="9560" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:02.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6875" number="1" />
                    <RELAYPOSITION athleteid="6957" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6905" number="3" />
                    <RELAYPOSITION athleteid="6961" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1595" points="151" reactiontime="+69" swimtime="00:03:19.24" resultid="6938" heatid="9497" lane="2" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:44.66" />
                    <SPLIT distance="150" swimtime="00:02:37.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6919" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="6888" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6909" number="3" />
                    <RELAYPOSITION athleteid="6900" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="5416" points="158" reactiontime="+80" swimtime="00:02:58.38" resultid="6940" heatid="9559" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:02:17.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6919" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6909" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="6888" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="6900" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1246" swimtime="00:02:32.26" resultid="6937" heatid="9353" lane="6" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:03.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6919" number="1" />
                    <RELAYPOSITION athleteid="6900" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="6915" number="3" />
                    <RELAYPOSITION athleteid="6892" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="400" agetotalmin="280" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="5602" reactiontime="+77" swimtime="00:03:00.05" resultid="6942" heatid="9607" lane="9" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:21.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6892" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6905" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="6909" number="3" />
                    <RELAYPOSITION athleteid="6919" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WSHS" nation="POL" clubid="7111" name="Wyższa Szkoła Humanitas w Sosnowcu">
          <ATHLETES>
            <ATHLETE birthdate="1996-03-24" firstname="Kinga" gender="F" lastname="Pluta" nation="POL" athleteid="7110">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="7113" heatid="9311" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="7114" heatid="9338" lane="3" entrytime="00:03:25.00" />
                <RESULT eventid="1458" points="314" reactiontime="+81" swimtime="00:00:39.79" resultid="7115" heatid="9445" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1493" points="342" swimtime="00:03:18.90" resultid="7116" heatid="9461" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="100" swimtime="00:01:33.64" />
                    <SPLIT distance="150" swimtime="00:02:25.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5279" points="379" reactiontime="+86" swimtime="00:01:28.54" resultid="7117" heatid="9501" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" status="DNS" swimtime="00:00:00.00" resultid="7118" heatid="9531" lane="8" entrytime="00:01:50.00" />
                <RESULT eventid="5534" status="DNS" swimtime="00:00:00.00" resultid="7119" heatid="9581" lane="4" entrytime="00:03:00.00" />
                <RESULT eventid="5568" points="404" reactiontime="+88" swimtime="00:00:39.75" resultid="7120" heatid="9593" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WAGR" nation="POL" region="WIE" clubid="6173" name="Wągrowiec">
          <CONTACT city="WĄGROWIEC" email="obywatel-ag @xl.wp.pl" name="GUZIAŁ ANDRZEJ" phone="508030407" state="WIELK" street="OS. NIEPODLEGŁOŚCI 9/4" zip="62-100" />
          <ATHLETES>
            <ATHLETE birthdate="1954-09-30" firstname="Andrzej" gender="M" lastname="Guział" nation="POL" athleteid="6174">
              <RESULTS>
                <RESULT eventid="1195" points="213" reactiontime="+98" swimtime="00:00:35.00" resultid="6175" heatid="9321" lane="9" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1280" points="130" reactiontime="+98" swimtime="00:14:50.34" resultid="6176" heatid="9362" lane="3" entrytime="00:13:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:30.44" />
                    <SPLIT distance="150" swimtime="00:02:23.60" />
                    <SPLIT distance="200" swimtime="00:03:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1510" points="210" swimtime="00:03:32.78" resultid="6177" heatid="9464" lane="1" entrytime="00:03:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="150" swimtime="00:02:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" points="207" swimtime="00:01:19.25" resultid="6178" heatid="9480" lane="6" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="206" reactiontime="+93" swimtime="00:01:36.71" resultid="6179" heatid="9507" lane="5" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5399" points="160" reactiontime="+91" swimtime="00:03:07.51" resultid="6180" heatid="9551" lane="2" entrytime="00:03:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:25.65" />
                    <SPLIT distance="150" swimtime="00:02:17.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="228" reactiontime="+88" swimtime="00:00:42.45" resultid="6181" heatid="9599" lane="2" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="5636" points="151" reactiontime="+98" swimtime="00:06:52.39" resultid="6182" heatid="9618" lane="4" entrytime="00:06:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:29.80" />
                    <SPLIT distance="150" swimtime="00:02:21.43" />
                    <SPLIT distance="200" swimtime="00:03:15.03" />
                    <SPLIT distance="250" swimtime="00:04:09.69" />
                    <SPLIT distance="300" swimtime="00:05:03.94" />
                    <SPLIT distance="350" swimtime="00:05:59.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="N" nation="POL" clubid="5822" name="Zawodnik Niezrzeszony">
          <CONTACT name="Karolina Szkudlarek" />
          <ATHLETES>
            <ATHLETE birthdate="1996-04-04" firstname="Karolina" gender="F" lastname="Szkudlarek" nation="POL" athleteid="5823">
              <RESULTS>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="5824" heatid="9314" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1458" points="431" reactiontime="+77" swimtime="00:00:35.82" resultid="5825" heatid="9446" lane="9" entrytime="00:00:34.50" />
                <RESULT eventid="1527" points="463" reactiontime="+82" swimtime="00:01:06.84" resultid="5826" heatid="9475" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5348" points="427" reactiontime="+69" swimtime="00:01:17.13" resultid="5827" heatid="9533" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5382" points="435" swimtime="00:02:29.02" resultid="5828" heatid="9547" lane="1" entrytime="00:02:24.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G2 - Pływak zanurzył się całkowicie w trakcie wyścigu (z wyjątkiem 15 m po starcie lub nawrocie)." eventid="5534" reactiontime="+75" status="DSQ" swimtime="00:02:50.56" resultid="5829" heatid="9582" lane="6" entrytime="00:02:42.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:07.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5619" points="394" reactiontime="+83" swimtime="00:05:22.38" resultid="5830" heatid="9609" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:01:56.80" />
                    <SPLIT distance="200" swimtime="00:02:37.82" />
                    <SPLIT distance="250" swimtime="00:03:19.14" />
                    <SPLIT distance="300" swimtime="00:04:00.82" />
                    <SPLIT distance="350" swimtime="00:04:41.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZUBR" nation="BLR" region="MINSK" clubid="6368" name="ZUBR Minsk">
          <CONTACT email="yauhenipuzan@gmail.com" name="Puzan Yauheni" phone="574504127" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-02" firstname="Aliaksandr" gender="M" lastname="Puzan" nation="BLR" athleteid="6369">
              <RESULTS>
                <RESULT eventid="1229" points="329" swimtime="00:02:45.01" resultid="6370" heatid="9346" lane="6" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:02:07.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1544" status="DNS" swimtime="00:00:00.00" resultid="6371" heatid="9487" lane="3" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1578" points="248" swimtime="00:02:57.45" resultid="6372" heatid="9495" lane="6" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5331" points="369" reactiontime="+73" swimtime="00:00:31.27" resultid="6373" heatid="9525" lane="0" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="5517" reactiontime="+60" status="DSQ" swimtime="00:01:11.77" resultid="6374" heatid="9576" lane="2" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-10" firstname="Siarhei" gender="M" lastname="Aliashkevich" nation="BLR" athleteid="6060">
              <RESULTS>
                <RESULT eventid="1229" points="440" reactiontime="+71" swimtime="00:02:29.86" resultid="6061" heatid="9348" lane="4" entrytime="00:02:28.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1476" points="437" reactiontime="+78" swimtime="00:00:31.66" resultid="6062" heatid="9456" lane="0" entrytime="00:00:31.38" entrycourse="LCM" />
                <RESULT eventid="5331" points="440" reactiontime="+78" swimtime="00:00:29.47" resultid="6063" heatid="9525" lane="3" entrytime="00:00:29.61" entrycourse="LCM" />
                <RESULT eventid="5399" points="418" reactiontime="+70" swimtime="00:02:16.39" resultid="6064" heatid="9557" lane="7" entrytime="00:02:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:07.90" />
                    <SPLIT distance="150" swimtime="00:01:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5517" points="434" swimtime="00:01:05.80" resultid="6065" heatid="9577" lane="9" entrytime="00:01:06.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5636" points="439" reactiontime="+73" swimtime="00:04:49.41" resultid="6066" heatid="9614" lane="2" entrytime="00:04:55.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:46.75" />
                    <SPLIT distance="200" swimtime="00:02:23.71" />
                    <SPLIT distance="250" swimtime="00:03:01.00" />
                    <SPLIT distance="300" swimtime="00:03:37.93" />
                    <SPLIT distance="350" swimtime="00:04:14.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-12" firstname="Roman" gender="M" lastname="Kostitsin" nation="BLR" athleteid="6067">
              <RESULTS>
                <RESULT eventid="1195" points="328" reactiontime="+89" swimtime="00:00:30.31" resultid="6068" heatid="9323" lane="4" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1510" points="307" swimtime="00:03:07.67" resultid="6069" heatid="9466" lane="6" entrytime="00:03:02.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:02:20.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5297" points="317" reactiontime="+79" swimtime="00:01:23.75" resultid="6070" heatid="9510" lane="2" entrytime="00:01:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5585" points="353" reactiontime="+73" swimtime="00:00:36.70" resultid="6071" heatid="9602" lane="5" entrytime="00:00:35.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KS Warszawianka" version="Build 21215">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Warszawa" name="Letnie Otwarte Mistrzostwa Polski w pływaniu w kat. MASTERS" course="LCM" nation="POL" timing="AUTOMATIC">
      <AGEDATE value="2012-05-26" type="YEAR" />
      <POOL lanemax="9" />
      <POINTTABLE pointtableid="3005" name="FINA Point Scoring" version="2012" />
      <SESSIONS>
        <SESSION date="2012-05-26" daytime="09:00" name="I  BLOK" number="1" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="1058" daytime="09:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1103" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4142" />
                    <RANKING order="2" place="2" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5156" />
                    <RANKING order="2" place="2" resultid="2414" />
                    <RANKING order="3" place="3" resultid="3236" />
                    <RANKING order="4" place="4" resultid="5140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3533" />
                    <RANKING order="2" place="2" resultid="3107" />
                    <RANKING order="3" place="3" resultid="4128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3130" />
                    <RANKING order="2" place="2" resultid="3912" />
                    <RANKING order="3" place="3" resultid="4012" />
                    <RANKING order="4" place="4" resultid="2625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                    <RANKING order="2" place="2" resultid="2459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3836" />
                    <RANKING order="2" place="2" resultid="3193" />
                    <RANKING order="3" place="3" resultid="3486" />
                    <RANKING order="4" place="4" resultid="4817" />
                    <RANKING order="5" place="5" resultid="5107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2448" />
                    <RANKING order="2" place="2" resultid="4054" />
                    <RANKING order="3" place="3" resultid="2265" />
                    <RANKING order="4" place="4" resultid="3956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4083" />
                    <RANKING order="2" place="2" resultid="4047" />
                    <RANKING order="3" place="3" resultid="3962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2402" />
                    <RANKING order="2" place="2" resultid="5682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1903" />
                    <RANKING order="2" place="2" resultid="1946" />
                    <RANKING order="3" place="3" resultid="4158" />
                    <RANKING order="4" place="4" resultid="3981" />
                    <RANKING order="5" place="5" resultid="2425" />
                    <RANKING order="6" place="-1" resultid="4941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="1101" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6970" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6971" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6972" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6973" daytime="09:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="09:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot;/20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2321" />
                    <RANKING order="2" place="2" resultid="4330" />
                    <RANKING order="3" place="3" resultid="3135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot;/25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3077" />
                    <RANKING order="2" place="2" resultid="4301" />
                    <RANKING order="3" place="3" resultid="4314" />
                    <RANKING order="4" place="4" resultid="4249" />
                    <RANKING order="5" place="5" resultid="3581" />
                    <RANKING order="6" place="6" resultid="4310" />
                    <RANKING order="7" place="7" resultid="2752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3876" />
                    <RANKING order="2" place="2" resultid="3451" />
                    <RANKING order="3" place="3" resultid="4206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3587" />
                    <RANKING order="2" place="2" resultid="3500" />
                    <RANKING order="3" place="3" resultid="3472" />
                    <RANKING order="4" place="4" resultid="2530" />
                    <RANKING order="5" place="5" resultid="2391" />
                    <RANKING order="6" place="6" resultid="3506" />
                    <RANKING order="7" place="7" resultid="3479" />
                    <RANKING order="8" place="8" resultid="3162" />
                    <RANKING order="9" place="9" resultid="2044" />
                    <RANKING order="10" place="10" resultid="4920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                    <RANKING order="2" place="2" resultid="2506" />
                    <RANKING order="3" place="3" resultid="2368" />
                    <RANKING order="4" place="4" resultid="2519" />
                    <RANKING order="5" place="5" resultid="3739" />
                    <RANKING order="6" place="6" resultid="3114" />
                    <RANKING order="7" place="-1" resultid="3743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;/45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4102" />
                    <RANKING order="2" place="2" resultid="2995" />
                    <RANKING order="3" place="3" resultid="1653" />
                    <RANKING order="4" place="4" resultid="3050" />
                    <RANKING order="5" place="-1" resultid="2307" />
                    <RANKING order="6" place="-1" resultid="3025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4236" />
                    <RANKING order="2" place="2" resultid="2831" />
                    <RANKING order="3" place="3" resultid="3002" />
                    <RANKING order="4" place="4" resultid="2853" />
                    <RANKING order="5" place="5" resultid="2345" />
                    <RANKING order="6" place="6" resultid="3142" />
                    <RANKING order="7" place="-1" resultid="2878" />
                    <RANKING order="8" place="-1" resultid="2746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1802" />
                    <RANKING order="2" place="2" resultid="2586" />
                    <RANKING order="3" place="3" resultid="2059" />
                    <RANKING order="4" place="4" resultid="2609" />
                    <RANKING order="5" place="5" resultid="2514" />
                    <RANKING order="6" place="6" resultid="3944" />
                    <RANKING order="7" place="-1" resultid="2051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5119" />
                    <RANKING order="2" place="2" resultid="1814" />
                    <RANKING order="3" place="3" resultid="3709" />
                    <RANKING order="4" place="4" resultid="3890" />
                    <RANKING order="5" place="5" resultid="1624" />
                    <RANKING order="6" place="6" resultid="3574" />
                    <RANKING order="7" place="7" resultid="4885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2687" />
                    <RANKING order="2" place="2" resultid="3902" />
                    <RANKING order="3" place="3" resultid="2784" />
                    <RANKING order="4" place="4" resultid="1742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1899" />
                    <RANKING order="2" place="2" resultid="3998" />
                    <RANKING order="3" place="3" resultid="3937" />
                    <RANKING order="4" place="4" resultid="4293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4031" />
                    <RANKING order="2" place="2" resultid="2981" />
                    <RANKING order="3" place="3" resultid="2682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6974" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6975" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6976" daytime="09:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6977" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6978" daytime="09:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6979" daytime="09:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6980" daytime="09:50" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="09:55" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7225" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1767" />
                    <RANKING order="2" place="2" resultid="1758" />
                    <RANKING order="3" place="3" resultid="3855" />
                    <RANKING order="4" place="-1" resultid="4060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7226" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2432" />
                    <RANKING order="2" place="2" resultid="3635" />
                    <RANKING order="3" place="3" resultid="4162" />
                    <RANKING order="4" place="4" resultid="2827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7227" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3674" />
                    <RANKING order="2" place="2" resultid="2300" />
                    <RANKING order="3" place="3" resultid="4224" />
                    <RANKING order="4" place="4" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7228" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                    <RANKING order="2" place="2" resultid="3913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7229" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3544" />
                    <RANKING order="2" place="2" resultid="2395" />
                    <RANKING order="3" place="3" resultid="2460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7230" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2407" />
                    <RANKING order="2" place="2" resultid="2553" />
                    <RANKING order="3" place="3" resultid="3551" />
                    <RANKING order="4" place="4" resultid="2915" />
                    <RANKING order="5" place="5" resultid="2802" />
                    <RANKING order="6" place="6" resultid="5100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7231" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1818" />
                    <RANKING order="2" place="2" resultid="1825" />
                    <RANKING order="3" place="3" resultid="4112" />
                    <RANKING order="4" place="4" resultid="3756" />
                    <RANKING order="5" place="5" resultid="3991" />
                    <RANKING order="6" place="6" resultid="2454" />
                    <RANKING order="7" place="7" resultid="2266" />
                    <RANKING order="8" place="-1" resultid="3957" />
                    <RANKING order="9" place="-1" resultid="4035" />
                    <RANKING order="10" place="-1" resultid="4055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7232" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1661" />
                    <RANKING order="2" place="2" resultid="2418" />
                    <RANKING order="3" place="3" resultid="1832" />
                    <RANKING order="4" place="4" resultid="3963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7233" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1929" />
                    <RANKING order="2" place="2" resultid="2935" />
                    <RANKING order="3" place="3" resultid="4017" />
                    <RANKING order="4" place="4" resultid="1664" />
                    <RANKING order="5" place="5" resultid="2773" />
                    <RANKING order="6" place="6" resultid="3969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7234" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1959" />
                    <RANKING order="2" place="2" resultid="4846" />
                    <RANKING order="3" place="3" resultid="3988" />
                    <RANKING order="4" place="4" resultid="3179" />
                    <RANKING order="5" place="5" resultid="1978" />
                    <RANKING order="6" place="6" resultid="4213" />
                    <RANKING order="7" place="7" resultid="2912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7235" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7236" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7237" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4190" />
                    <RANKING order="2" place="2" resultid="4901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7238" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3951" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6981" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6982" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6983" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6984" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6985" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6986" daytime="10:05" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1134" daytime="10:05" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7239" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5685" />
                    <RANKING order="2" place="2" resultid="4255" />
                    <RANKING order="3" place="3" resultid="3919" />
                    <RANKING order="4" place="4" resultid="4325" />
                    <RANKING order="5" place="5" resultid="4153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7240" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5067" />
                    <RANKING order="2" place="2" resultid="3820" />
                    <RANKING order="3" place="3" resultid="1618" />
                    <RANKING order="4" place="4" resultid="3172" />
                    <RANKING order="5" place="5" resultid="2560" />
                    <RANKING order="6" place="6" resultid="2872" />
                    <RANKING order="7" place="-1" resultid="4321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7241" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3070" />
                    <RANKING order="2" place="2" resultid="4207" />
                    <RANKING order="3" place="3" resultid="2939" />
                    <RANKING order="4" place="4" resultid="3862" />
                    <RANKING order="5" place="5" resultid="4125" />
                    <RANKING order="6" place="6" resultid="3897" />
                    <RANKING order="7" place="7" resultid="3155" />
                    <RANKING order="8" place="8" resultid="3883" />
                    <RANKING order="9" place="-1" resultid="2814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7242" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3020" />
                    <RANKING order="2" place="2" resultid="3438" />
                    <RANKING order="3" place="3" resultid="3040" />
                    <RANKING order="4" place="4" resultid="2632" />
                    <RANKING order="5" place="5" resultid="2292" />
                    <RANKING order="6" place="6" resultid="4859" />
                    <RANKING order="7" place="7" resultid="4972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7243" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3123" />
                    <RANKING order="2" place="2" resultid="3168" />
                    <RANKING order="3" place="3" resultid="1919" />
                    <RANKING order="4" place="4" resultid="1924" />
                    <RANKING order="5" place="5" resultid="2356" />
                    <RANKING order="6" place="6" resultid="2921" />
                    <RANKING order="7" place="7" resultid="4967" />
                    <RANKING order="8" place="8" resultid="3726" />
                    <RANKING order="9" place="9" resultid="3431" />
                    <RANKING order="10" place="10" resultid="2780" />
                    <RANKING order="11" place="11" resultid="1690" />
                    <RANKING order="12" place="12" resultid="3210" />
                    <RANKING order="13" place="13" resultid="4924" />
                    <RANKING order="14" place="14" resultid="5125" />
                    <RANKING order="15" place="15" resultid="3115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7244" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3045" />
                    <RANKING order="2" place="2" resultid="1634" />
                    <RANKING order="3" place="3" resultid="4824" />
                    <RANKING order="4" place="4" resultid="4217" />
                    <RANKING order="5" place="5" resultid="2821" />
                    <RANKING order="6" place="6" resultid="2574" />
                    <RANKING order="7" place="7" resultid="3493" />
                    <RANKING order="8" place="8" resultid="3702" />
                    <RANKING order="9" place="9" resultid="2338" />
                    <RANKING order="10" place="10" resultid="3051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7245" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3064" />
                    <RANKING order="2" place="2" resultid="2380" />
                    <RANKING order="3" place="3" resultid="2832" />
                    <RANKING order="4" place="4" resultid="5585" />
                    <RANKING order="5" place="5" resultid="2523" />
                    <RANKING order="6" place="6" resultid="2616" />
                    <RANKING order="7" place="7" resultid="1750" />
                    <RANKING order="8" place="-1" resultid="1726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7246" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1797" />
                    <RANKING order="2" place="2" resultid="3032" />
                    <RANKING order="3" place="3" resultid="5675" />
                    <RANKING order="4" place="4" resultid="4097" />
                    <RANKING order="5" place="5" resultid="3593" />
                    <RANKING order="6" place="6" resultid="2673" />
                    <RANKING order="7" place="7" resultid="1893" />
                    <RANKING order="8" place="8" resultid="4913" />
                    <RANKING order="9" place="-1" resultid="3695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7247" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4834" />
                    <RANKING order="2" place="2" resultid="2661" />
                    <RANKING order="3" place="3" resultid="3869" />
                    <RANKING order="4" place="4" resultid="4088" />
                    <RANKING order="5" place="5" resultid="3458" />
                    <RANKING order="6" place="6" resultid="1935" />
                    <RANKING order="7" place="7" resultid="1698" />
                    <RANKING order="8" place="8" resultid="2037" />
                    <RANKING order="9" place="9" resultid="4005" />
                    <RANKING order="10" place="10" resultid="2990" />
                    <RANKING order="11" place="11" resultid="3891" />
                    <RANKING order="12" place="12" resultid="2668" />
                    <RANKING order="13" place="13" resultid="1982" />
                    <RANKING order="14" place="14" resultid="3083" />
                    <RANKING order="15" place="15" resultid="1849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7248" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2951" />
                    <RANKING order="2" place="2" resultid="1942" />
                    <RANKING order="3" place="3" resultid="3057" />
                    <RANKING order="4" place="4" resultid="3903" />
                    <RANKING order="5" place="5" resultid="1701" />
                    <RANKING order="6" place="6" resultid="1743" />
                    <RANKING order="7" place="7" resultid="2362" />
                    <RANKING order="8" place="8" resultid="1888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7249" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1952" />
                    <RANKING order="2" place="2" resultid="2847" />
                    <RANKING order="3" place="3" resultid="3681" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="5" resultid="4294" />
                    <RANKING order="6" place="-1" resultid="3688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7250" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2654" />
                    <RANKING order="2" place="2" resultid="1880" />
                    <RANKING order="3" place="3" resultid="3649" />
                    <RANKING order="4" place="4" resultid="2329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7251" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                    <RANKING order="2" place="2" resultid="3568" />
                    <RANKING order="3" place="3" resultid="3826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7252" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2896" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6987" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6988" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6989" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6990" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6991" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6992" daytime="10:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6993" daytime="10:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6994" daytime="10:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6995" daytime="10:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6996" daytime="10:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6997" daytime="10:20" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1149" daytime="10:20" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1151" agemax="119" agemin="100" name="KATEGORIA: &quot;A&quot;/100-119/" calculate="TOTAL" />
                <AGEGROUP agegroupid="1152" agemax="159" agemin="120" name="KATEGORIA: &quot;B&quot;/120-159/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="7218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="199" agemin="160" name="KATEGORIA: &quot;C&quot;/160-199/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="239" agemin="200" name="KATEGORIA: &quot;D&quot;/200-239/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2469" />
                    <RANKING order="2" place="2" resultid="7220" />
                    <RANKING order="3" place="3" resultid="7591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="279" agemin="240" name="KATEGORIA: &quot;E&quot;/240-279/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1989" />
                    <RANKING order="2" place="2" resultid="3975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="-1" agemin="280" name="KATEGORIA: &quot;F&quot;/280 i starsi/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4945" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6998" daytime="10:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1164" daytime="10:30" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1588" agemax="119" agemin="100" name="KATEGORIA: &quot;A&quot;/100-119/" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6967" />
                    <RANKING order="2" place="2" resultid="4466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="159" agemin="120" name="KATEGORIA: &quot;B&quot;/120-159/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4269" />
                    <RANKING order="2" place="2" resultid="3512" />
                    <RANKING order="3" place="3" resultid="1991" />
                    <RANKING order="4" place="4" resultid="7224" />
                    <RANKING order="5" place="5" resultid="6966" />
                    <RANKING order="6" place="6" resultid="6965" />
                    <RANKING order="7" place="-1" resultid="7216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="199" agemin="160" name="KATEGORIA: &quot;C&quot;/160-199/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7215" />
                    <RANKING order="2" place="2" resultid="2467" />
                    <RANKING order="3" place="3" resultid="7221" />
                    <RANKING order="4" place="4" resultid="7212" />
                    <RANKING order="5" place="5" resultid="4984" />
                    <RANKING order="6" place="-1" resultid="2837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="239" agemin="200" name="KATEGORIA: &quot;D&quot;/200-239/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3513" />
                    <RANKING order="2" place="2" resultid="2472" />
                    <RANKING order="3" place="3" resultid="4106" />
                    <RANKING order="4" place="-1" resultid="7217" />
                    <RANKING order="5" place="-1" resultid="3715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1592" agemax="279" agemin="240" name="KATEGORIA: &quot;E&quot;/240-279/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1990" />
                    <RANKING order="2" place="2" resultid="1838" />
                    <RANKING order="3" place="3" resultid="7176" />
                    <RANKING order="4" place="-1" resultid="3925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1593" agemax="-1" agemin="280" name="KATEGORIA: &quot;F&quot;/280 i starsi/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7223" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6999" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7000" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7001" daytime="10:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="10:40" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7253" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1773" />
                    <RANKING order="2" place="2" resultid="1759" />
                    <RANKING order="3" place="3" resultid="3856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7254" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3636" />
                    <RANKING order="2" place="2" resultid="5141" />
                    <RANKING order="3" place="3" resultid="4842" />
                    <RANKING order="4" place="4" resultid="3666" />
                    <RANKING order="5" place="5" resultid="4163" />
                    <RANKING order="6" place="6" resultid="5482" />
                    <RANKING order="7" place="7" resultid="1649" />
                    <RANKING order="8" place="-1" resultid="3814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7255" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3417" />
                    <RANKING order="2" place="2" resultid="2570" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="4" resultid="5582" />
                    <RANKING order="5" place="5" resultid="2301" />
                    <RANKING order="6" place="6" resultid="3108" />
                    <RANKING order="7" place="7" resultid="4129" />
                    <RANKING order="8" place="8" resultid="3091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7256" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4290" />
                    <RANKING order="2" place="2" resultid="1791" />
                    <RANKING order="3" place="3" resultid="2626" />
                    <RANKING order="4" place="4" resultid="3010" />
                    <RANKING order="5" place="5" resultid="4849" />
                    <RANKING order="6" place="6" resultid="2437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7257" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1914" />
                    <RANKING order="2" place="2" resultid="5136" />
                    <RANKING order="3" place="3" resultid="3545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7258" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2868" />
                    <RANKING order="2" place="2" resultid="2408" />
                    <RANKING order="3" place="3" resultid="2554" />
                    <RANKING order="4" place="4" resultid="4818" />
                    <RANKING order="5" place="5" resultid="2442" />
                    <RANKING order="6" place="6" resultid="3487" />
                    <RANKING order="7" place="7" resultid="2803" />
                    <RANKING order="8" place="8" resultid="2947" />
                    <RANKING order="9" place="9" resultid="5108" />
                    <RANKING order="10" place="10" resultid="5101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7259" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1826" />
                    <RANKING order="2" place="2" resultid="4113" />
                    <RANKING order="3" place="3" resultid="1819" />
                    <RANKING order="4" place="4" resultid="2449" />
                    <RANKING order="5" place="5" resultid="4036" />
                    <RANKING order="6" place="6" resultid="2603" />
                    <RANKING order="7" place="7" resultid="2455" />
                    <RANKING order="8" place="8" resultid="3992" />
                    <RANKING order="9" place="9" resultid="2581" />
                    <RANKING order="10" place="10" resultid="2272" />
                    <RANKING order="11" place="-1" resultid="4024" />
                    <RANKING order="12" place="-1" resultid="4042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7260" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1833" />
                    <RANKING order="2" place="2" resultid="5114" />
                    <RANKING order="3" place="3" resultid="4048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7261" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4077" />
                    <RANKING order="2" place="2" resultid="1938" />
                    <RANKING order="3" place="3" resultid="2774" />
                    <RANKING order="4" place="4" resultid="3217" />
                    <RANKING order="5" place="5" resultid="3970" />
                    <RANKING order="6" place="-1" resultid="4895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7262" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3180" />
                    <RANKING order="2" place="2" resultid="2908" />
                    <RANKING order="3" place="3" resultid="2426" />
                    <RANKING order="4" place="4" resultid="3982" />
                    <RANKING order="5" place="5" resultid="4942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7263" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4932" />
                    <RANKING order="2" place="2" resultid="3807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7264" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7265" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7266" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3952" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7002" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7003" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7004" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7005" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7006" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7007" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7008" daytime="10:50" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1194" daytime="10:55" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7267" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5037" />
                    <RANKING order="2" place="2" resultid="3677" />
                    <RANKING order="3" place="3" resultid="3559" />
                    <RANKING order="4" place="4" resultid="3136" />
                    <RANKING order="5" place="5" resultid="3920" />
                    <RANKING order="6" place="6" resultid="2332" />
                    <RANKING order="7" place="7" resultid="4256" />
                    <RANKING order="8" place="-1" resultid="5062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7268" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2546" />
                    <RANKING order="2" place="2" resultid="1857" />
                    <RANKING order="3" place="3" resultid="3771" />
                    <RANKING order="4" place="4" resultid="4200" />
                    <RANKING order="5" place="5" resultid="4230" />
                    <RANKING order="6" place="6" resultid="4306" />
                    <RANKING order="7" place="7" resultid="3149" />
                    <RANKING order="8" place="8" resultid="3790" />
                    <RANKING order="9" place="9" resultid="4315" />
                    <RANKING order="10" place="10" resultid="3173" />
                    <RANKING order="11" place="11" resultid="1777" />
                    <RANKING order="12" place="12" resultid="4250" />
                    <RANKING order="13" place="13" resultid="4135" />
                    <RANKING order="14" place="14" resultid="1986" />
                    <RANKING order="15" place="15" resultid="1867" />
                    <RANKING order="16" place="16" resultid="5056" />
                    <RANKING order="17" place="17" resultid="3582" />
                    <RANKING order="18" place="18" resultid="1630" />
                    <RANKING order="19" place="19" resultid="4260" />
                    <RANKING order="20" place="-1" resultid="4182" />
                    <RANKING order="21" place="-1" resultid="2873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7269" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1862" />
                    <RANKING order="2" place="2" resultid="5034" />
                    <RANKING order="3" place="3" resultid="3877" />
                    <RANKING order="4" place="4" resultid="3844" />
                    <RANKING order="5" place="5" resultid="3071" />
                    <RANKING order="6" place="6" resultid="3863" />
                    <RANKING order="7" place="7" resultid="3608" />
                    <RANKING order="8" place="8" resultid="2973" />
                    <RANKING order="9" place="9" resultid="3537" />
                    <RANKING order="10" place="10" resultid="3156" />
                    <RANKING order="11" place="11" resultid="5653" />
                    <RANKING order="12" place="-1" resultid="1873" />
                    <RANKING order="13" place="-1" resultid="2815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7270" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2864" />
                    <RANKING order="2" place="2" resultid="3439" />
                    <RANKING order="3" place="3" resultid="3473" />
                    <RANKING order="4" place="4" resultid="2633" />
                    <RANKING order="5" place="5" resultid="3611" />
                    <RANKING order="6" place="6" resultid="2293" />
                    <RANKING order="7" place="7" resultid="2564" />
                    <RANKING order="8" place="8" resultid="5584" />
                    <RANKING order="9" place="9" resultid="5073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7271" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2357" />
                    <RANKING order="2" place="2" resultid="4961" />
                    <RANKING order="3" place="3" resultid="3432" />
                    <RANKING order="4" place="4" resultid="5126" />
                    <RANKING order="5" place="5" resultid="3727" />
                    <RANKING order="6" place="6" resultid="1704" />
                    <RANKING order="7" place="7" resultid="3211" />
                    <RANKING order="8" place="8" resultid="5047" />
                    <RANKING order="9" place="9" resultid="3186" />
                    <RANKING order="10" place="10" resultid="4925" />
                    <RANKING order="11" place="11" resultid="1974" />
                    <RANKING order="12" place="12" resultid="3744" />
                    <RANKING order="13" place="13" resultid="3116" />
                    <RANKING order="14" place="-1" resultid="3782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7272" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3642" />
                    <RANKING order="2" place="2" resultid="2592" />
                    <RANKING order="3" place="3" resultid="4218" />
                    <RANKING order="4" place="4" resultid="1635" />
                    <RANKING order="5" place="5" resultid="4285" />
                    <RANKING order="6" place="6" resultid="1654" />
                    <RANKING order="7" place="7" resultid="2822" />
                    <RANKING order="8" place="8" resultid="2996" />
                    <RANKING order="9" place="9" resultid="3703" />
                    <RANKING order="10" place="10" resultid="2339" />
                    <RANKING order="11" place="11" resultid="2575" />
                    <RANKING order="12" place="12" resultid="3052" />
                    <RANKING order="13" place="13" resultid="3015" />
                    <RANKING order="14" place="-1" resultid="2308" />
                    <RANKING order="15" place="-1" resultid="1683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7273" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3065" />
                    <RANKING order="2" place="2" resultid="2809" />
                    <RANKING order="3" place="3" resultid="3465" />
                    <RANKING order="4" place="4" resultid="1786" />
                    <RANKING order="5" place="5" resultid="4237" />
                    <RANKING order="6" place="6" resultid="2931" />
                    <RANKING order="7" place="7" resultid="6419" />
                    <RANKING order="8" place="8" resultid="1751" />
                    <RANKING order="9" place="9" resultid="2346" />
                    <RANKING order="10" place="10" resultid="3143" />
                    <RANKING order="11" place="-1" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7274" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3033" />
                    <RANKING order="2" place="2" resultid="1894" />
                    <RANKING order="3" place="3" resultid="2674" />
                    <RANKING order="4" place="4" resultid="4168" />
                    <RANKING order="5" place="5" resultid="3594" />
                    <RANKING order="6" place="6" resultid="1722" />
                    <RANKING order="7" place="7" resultid="3795" />
                    <RANKING order="8" place="8" resultid="2610" />
                    <RANKING order="9" place="9" resultid="4914" />
                    <RANKING order="10" place="10" resultid="6691" />
                    <RANKING order="11" place="11" resultid="3945" />
                    <RANKING order="12" place="-1" resultid="4910" />
                    <RANKING order="13" place="-1" resultid="3696" />
                    <RANKING order="14" place="-1" resultid="5478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7275" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4835" />
                    <RANKING order="2" place="2" resultid="2662" />
                    <RANKING order="3" place="3" resultid="3870" />
                    <RANKING order="4" place="4" resultid="4175" />
                    <RANKING order="5" place="5" resultid="4242" />
                    <RANKING order="6" place="6" resultid="1909" />
                    <RANKING order="7" place="7" resultid="3459" />
                    <RANKING order="8" place="8" resultid="3084" />
                    <RANKING order="9" place="9" resultid="4006" />
                    <RANKING order="10" place="10" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7276" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2952" />
                    <RANKING order="2" place="2" resultid="1809" />
                    <RANKING order="3" place="3" resultid="2688" />
                    <RANKING order="4" place="4" resultid="2373" />
                    <RANKING order="5" place="5" resultid="3058" />
                    <RANKING order="6" place="6" resultid="2901" />
                    <RANKING order="7" place="7" resultid="2785" />
                    <RANKING order="8" place="8" resultid="2363" />
                    <RANKING order="9" place="9" resultid="1889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7277" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                    <RANKING order="2" place="2" resultid="3999" />
                    <RANKING order="3" place="3" resultid="3849" />
                    <RANKING order="4" place="-1" resultid="3689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7278" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2655" />
                    <RANKING order="2" place="2" resultid="1881" />
                    <RANKING order="3" place="3" resultid="3650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7279" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3658" />
                    <RANKING order="2" place="2" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7280" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2897" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7009" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7010" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7011" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7012" daytime="11:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7013" daytime="11:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7014" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7015" daytime="11:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7016" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7017" daytime="11:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7018" daytime="11:15" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7019" daytime="11:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7020" daytime="11:20" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7021" daytime="11:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7022" daytime="11:20" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1209" daytime="11:25" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7281" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/" />
                <AGEGROUP agegroupid="7282" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7283" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2622" />
                    <RANKING order="2" place="2" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7284" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/" />
                <AGEGROUP agegroupid="7285" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/" />
                <AGEGROUP agegroupid="7286" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3837" />
                    <RANKING order="2" place="2" resultid="3552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7287" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4025" />
                    <RANKING order="2" place="2" resultid="1643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7288" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7289" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1930" />
                    <RANKING order="2" place="2" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7290" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7291" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/" />
                <AGEGROUP agegroupid="7292" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7293" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7294" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7023" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7024" daytime="11:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="11:35" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7295" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3762" />
                    <RANKING order="2" place="2" resultid="2322" />
                    <RANKING order="3" place="3" resultid="3560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7296" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5030" />
                    <RANKING order="2" place="2" resultid="1968" />
                    <RANKING order="3" place="-1" resultid="4183" />
                    <RANKING order="4" place="-1" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7297" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1963" />
                    <RANKING order="2" place="2" resultid="3884" />
                    <RANKING order="3" place="3" resultid="4854" />
                    <RANKING order="4" place="4" resultid="3452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7298" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3445" />
                    <RANKING order="2" place="2" resultid="2386" />
                    <RANKING order="3" place="3" resultid="4973" />
                    <RANKING order="4" place="4" resultid="3507" />
                    <RANKING order="5" place="5" resultid="2045" />
                    <RANKING order="6" place="-1" resultid="3480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7299" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3124" />
                    <RANKING order="2" place="2" resultid="2352" />
                    <RANKING order="3" place="3" resultid="1733" />
                    <RANKING order="4" place="4" resultid="2892" />
                    <RANKING order="5" place="5" resultid="2507" />
                    <RANKING order="6" place="6" resultid="4979" />
                    <RANKING order="7" place="7" resultid="5048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7300" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1641" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="3494" />
                    <RANKING order="4" place="-1" resultid="3026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7301" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2888" />
                    <RANKING order="2" place="2" resultid="2854" />
                    <RANKING order="3" place="3" resultid="3466" />
                    <RANKING order="4" place="-1" resultid="6422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7302" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5676" />
                    <RANKING order="2" place="2" resultid="4120" />
                    <RANKING order="3" place="3" resultid="2060" />
                    <RANKING order="4" place="4" resultid="4092" />
                    <RANKING order="5" place="-1" resultid="2052" />
                    <RANKING order="6" place="-1" resultid="1803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7303" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4243" />
                    <RANKING order="2" place="2" resultid="3710" />
                    <RANKING order="3" place="3" resultid="2038" />
                    <RANKING order="4" place="4" resultid="4886" />
                    <RANKING order="5" place="5" resultid="1850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7304" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7305" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3682" />
                    <RANKING order="2" place="2" resultid="3938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7306" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7307" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7308" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7025" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7026" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7027" daytime="11:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7028" daytime="11:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7029" daytime="11:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2012-05-26" daytime="16:00" name="II BLOK" number="2" warmupfrom="15:00" warmupuntil="15:45">
          <EVENTS>
            <EVENT eventid="1240" daytime="16:00" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7309" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7310" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5485" />
                    <RANKING order="2" place="2" resultid="4843" />
                    <RANKING order="3" place="3" resultid="3103" />
                    <RANKING order="4" place="4" resultid="3637" />
                    <RANKING order="5" place="5" resultid="3237" />
                    <RANKING order="6" place="6" resultid="5483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7311" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3418" />
                    <RANKING order="2" place="2" resultid="4266" />
                    <RANKING order="3" place="3" resultid="2302" />
                    <RANKING order="4" place="4" resultid="2280" />
                    <RANKING order="5" place="5" resultid="3205" />
                    <RANKING order="6" place="6" resultid="3092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7312" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                    <RANKING order="2" place="2" resultid="2925" />
                    <RANKING order="3" place="3" resultid="3914" />
                    <RANKING order="4" place="4" resultid="4850" />
                    <RANKING order="5" place="5" resultid="2928" />
                    <RANKING order="6" place="6" resultid="2627" />
                    <RANKING order="7" place="7" resultid="2438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7313" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3190" />
                    <RANKING order="2" place="2" resultid="4138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7314" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3838" />
                    <RANKING order="2" place="2" resultid="2443" />
                    <RANKING order="3" place="3" resultid="3488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7315" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1820" />
                    <RANKING order="2" place="2" resultid="4037" />
                    <RANKING order="3" place="3" resultid="3757" />
                    <RANKING order="4" place="4" resultid="2456" />
                    <RANKING order="5" place="5" resultid="3993" />
                    <RANKING order="6" place="6" resultid="1675" />
                    <RANKING order="7" place="7" resultid="2604" />
                    <RANKING order="8" place="8" resultid="2273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7316" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2420" />
                    <RANKING order="2" place="2" resultid="1834" />
                    <RANKING order="3" place="3" resultid="4049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7317" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1931" />
                    <RANKING order="2" place="2" resultid="4078" />
                    <RANKING order="3" place="3" resultid="2775" />
                    <RANKING order="4" place="4" resultid="4019" />
                    <RANKING order="5" place="-1" resultid="4896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7318" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1960" />
                    <RANKING order="2" place="2" resultid="3181" />
                    <RANKING order="3" place="3" resultid="3983" />
                    <RANKING order="4" place="4" resultid="2427" />
                    <RANKING order="5" place="-1" resultid="1948" />
                    <RANKING order="6" place="-1" resultid="4943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7319" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7320" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7321" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7322" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7030" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7031" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7032" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7033" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7034" daytime="16:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="16:10" gender="M" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7323" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5097" />
                    <RANKING order="2" place="2" resultid="3678" />
                    <RANKING order="3" place="3" resultid="3561" />
                    <RANKING order="4" place="4" resultid="3137" />
                    <RANKING order="5" place="5" resultid="3921" />
                    <RANKING order="6" place="-1" resultid="5063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7324" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2547" />
                    <RANKING order="2" place="2" resultid="3671" />
                    <RANKING order="3" place="3" resultid="1858" />
                    <RANKING order="4" place="4" resultid="2296" />
                    <RANKING order="5" place="5" resultid="5031" />
                    <RANKING order="6" place="6" resultid="4874" />
                    <RANKING order="7" place="7" resultid="5068" />
                    <RANKING order="8" place="8" resultid="4201" />
                    <RANKING order="9" place="9" resultid="4231" />
                    <RANKING order="10" place="10" resultid="4307" />
                    <RANKING order="11" place="11" resultid="3150" />
                    <RANKING order="12" place="12" resultid="3791" />
                    <RANKING order="13" place="13" resultid="4184" />
                    <RANKING order="14" place="14" resultid="1868" />
                    <RANKING order="15" place="15" resultid="5057" />
                    <RANKING order="16" place="16" resultid="5092" />
                    <RANKING order="17" place="17" resultid="1987" />
                    <RANKING order="18" place="18" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7325" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4208" />
                    <RANKING order="2" place="2" resultid="2940" />
                    <RANKING order="3" place="3" resultid="3609" />
                    <RANKING order="4" place="4" resultid="1874" />
                    <RANKING order="5" place="5" resultid="3538" />
                    <RANKING order="6" place="6" resultid="3898" />
                    <RANKING order="7" place="7" resultid="3885" />
                    <RANKING order="8" place="8" resultid="2974" />
                    <RANKING order="9" place="9" resultid="5654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7326" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3021" />
                    <RANKING order="2" place="2" resultid="3446" />
                    <RANKING order="3" place="3" resultid="5490" />
                    <RANKING order="4" place="4" resultid="3750" />
                    <RANKING order="5" place="5" resultid="3612" />
                    <RANKING order="6" place="6" resultid="2634" />
                    <RANKING order="7" place="7" resultid="2387" />
                    <RANKING order="8" place="8" resultid="4974" />
                    <RANKING order="9" place="9" resultid="3440" />
                    <RANKING order="10" place="10" resultid="4514" />
                    <RANKING order="11" place="11" resultid="3163" />
                    <RANKING order="12" place="-1" resultid="3631" />
                    <RANKING order="13" place="-1" resultid="2944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7327" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3125" />
                    <RANKING order="2" place="2" resultid="1920" />
                    <RANKING order="3" place="3" resultid="1734" />
                    <RANKING order="4" place="4" resultid="2353" />
                    <RANKING order="5" place="5" resultid="2369" />
                    <RANKING order="6" place="6" resultid="2893" />
                    <RANKING order="7" place="7" resultid="3728" />
                    <RANKING order="8" place="8" resultid="4980" />
                    <RANKING order="9" place="9" resultid="5127" />
                    <RANKING order="10" place="10" resultid="5049" />
                    <RANKING order="11" place="11" resultid="3187" />
                    <RANKING order="12" place="12" resultid="1975" />
                    <RANKING order="13" place="13" resultid="3745" />
                    <RANKING order="14" place="-1" resultid="3212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7328" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1636" />
                    <RANKING order="2" place="2" resultid="2593" />
                    <RANKING order="3" place="3" resultid="4825" />
                    <RANKING order="4" place="4" resultid="3495" />
                    <RANKING order="5" place="5" resultid="3704" />
                    <RANKING order="6" place="6" resultid="2796" />
                    <RANKING order="7" place="-1" resultid="3027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7329" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3066" />
                    <RANKING order="2" place="2" resultid="2381" />
                    <RANKING order="3" place="3" resultid="4828" />
                    <RANKING order="4" place="4" resultid="2855" />
                    <RANKING order="5" place="5" resultid="1752" />
                    <RANKING order="6" place="6" resultid="5161" />
                    <RANKING order="7" place="7" resultid="3003" />
                    <RANKING order="8" place="8" resultid="3776" />
                    <RANKING order="9" place="9" resultid="3144" />
                    <RANKING order="10" place="10" resultid="2617" />
                    <RANKING order="11" place="-1" resultid="2747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7330" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1798" />
                    <RANKING order="2" place="2" resultid="1781" />
                    <RANKING order="3" place="3" resultid="2587" />
                    <RANKING order="4" place="4" resultid="1729" />
                    <RANKING order="5" place="5" resultid="2675" />
                    <RANKING order="6" place="6" resultid="4169" />
                    <RANKING order="7" place="7" resultid="3595" />
                    <RANKING order="8" place="8" resultid="1723" />
                    <RANKING order="9" place="9" resultid="2515" />
                    <RANKING order="10" place="10" resultid="3946" />
                    <RANKING order="11" place="-1" resultid="5479" />
                    <RANKING order="12" place="-1" resultid="3697" />
                    <RANKING order="13" place="-1" resultid="6692" />
                    <RANKING order="14" place="-1" resultid="3796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7331" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4244" />
                    <RANKING order="2" place="2" resultid="4836" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="3871" />
                    <RANKING order="5" place="5" resultid="1910" />
                    <RANKING order="6" place="6" resultid="3085" />
                    <RANKING order="7" place="7" resultid="1983" />
                    <RANKING order="8" place="8" resultid="2669" />
                    <RANKING order="9" place="9" resultid="1851" />
                    <RANKING order="10" place="-1" resultid="4007" />
                    <RANKING order="11" place="-1" resultid="4176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7332" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2689" />
                    <RANKING order="2" place="2" resultid="1810" />
                    <RANKING order="3" place="3" resultid="2905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7333" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2884" />
                    <RANKING order="2" place="2" resultid="3939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7334" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7335" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7336" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7035" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7036" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7037" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7038" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7039" daytime="16:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7040" daytime="16:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7041" daytime="16:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7042" daytime="16:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7043" daytime="16:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7044" daytime="16:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7045" daytime="16:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7046" daytime="16:25" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1271" daytime="16:25" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7337" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4143" />
                    <RANKING order="2" place="2" resultid="1768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7338" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2433" />
                    <RANKING order="2" place="2" resultid="5157" />
                    <RANKING order="3" place="3" resultid="2415" />
                    <RANKING order="4" place="4" resultid="4164" />
                    <RANKING order="5" place="5" resultid="5142" />
                    <RANKING order="6" place="-1" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7339" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3534" />
                    <RANKING order="2" place="2" resultid="3109" />
                    <RANKING order="3" place="3" resultid="3591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7340" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3131" />
                    <RANKING order="2" place="2" resultid="3915" />
                    <RANKING order="3" place="3" resultid="4013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7341" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3191" />
                    <RANKING order="2" place="2" resultid="1915" />
                    <RANKING order="3" place="3" resultid="2461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7342" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2410" />
                    <RANKING order="2" place="2" resultid="3194" />
                    <RANKING order="3" place="3" resultid="5109" />
                    <RANKING order="4" place="4" resultid="4879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7343" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1827" />
                    <RANKING order="2" place="2" resultid="2450" />
                    <RANKING order="3" place="3" resultid="4038" />
                    <RANKING order="4" place="4" resultid="1667" />
                    <RANKING order="5" place="5" resultid="2267" />
                    <RANKING order="6" place="6" resultid="4917" />
                    <RANKING order="7" place="7" resultid="3958" />
                    <RANKING order="8" place="8" resultid="4043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7344" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4084" />
                    <RANKING order="2" place="2" resultid="3964" />
                    <RANKING order="3" place="3" resultid="3600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7345" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2403" />
                    <RANKING order="2" place="2" resultid="3006" />
                    <RANKING order="3" place="3" resultid="3971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7346" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1949" />
                    <RANKING order="2" place="2" resultid="1979" />
                    <RANKING order="3" place="3" resultid="4159" />
                    <RANKING order="4" place="4" resultid="1905" />
                    <RANKING order="5" place="5" resultid="4214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7347" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7348" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7349" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7350" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7047" daytime="16:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7048" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7049" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7050" daytime="16:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7051" daytime="16:35" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="16:35" gender="M" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7351" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2323" />
                    <RANKING order="2" place="2" resultid="5088" />
                    <RANKING order="3" place="3" resultid="4331" />
                    <RANKING order="4" place="4" resultid="3922" />
                    <RANKING order="5" place="5" resultid="2333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7352" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4875" />
                    <RANKING order="2" place="2" resultid="3078" />
                    <RANKING order="3" place="3" resultid="4302" />
                    <RANKING order="4" place="4" resultid="5474" />
                    <RANKING order="5" place="5" resultid="3583" />
                    <RANKING order="6" place="6" resultid="4311" />
                    <RANKING order="7" place="7" resultid="5093" />
                    <RANKING order="8" place="8" resultid="2754" />
                    <RANKING order="9" place="9" resultid="4261" />
                    <RANKING order="10" place="-1" resultid="4316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7353" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4209" />
                    <RANKING order="2" place="2" resultid="1695" />
                    <RANKING order="3" place="3" resultid="3864" />
                    <RANKING order="4" place="4" resultid="3453" />
                    <RANKING order="5" place="5" resultid="3626" />
                    <RANKING order="6" place="6" resultid="5501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7354" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3501" />
                    <RANKING order="2" place="2" resultid="3588" />
                    <RANKING order="3" place="3" resultid="1707" />
                    <RANKING order="4" place="4" resultid="3474" />
                    <RANKING order="5" place="5" resultid="1716" />
                    <RANKING order="6" place="6" resultid="4860" />
                    <RANKING order="7" place="7" resultid="3481" />
                    <RANKING order="8" place="8" resultid="2565" />
                    <RANKING order="9" place="8" resultid="5074" />
                    <RANKING order="10" place="10" resultid="3508" />
                    <RANKING order="11" place="11" resultid="4921" />
                    <RANKING order="12" place="-1" resultid="2294" />
                    <RANKING order="13" place="-1" resultid="2531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7355" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4938" />
                    <RANKING order="2" place="2" resultid="3425" />
                    <RANKING order="3" place="3" resultid="1921" />
                    <RANKING order="4" place="4" resultid="2508" />
                    <RANKING order="5" place="5" resultid="2370" />
                    <RANKING order="6" place="6" resultid="3213" />
                    <RANKING order="7" place="7" resultid="2520" />
                    <RANKING order="8" place="8" resultid="1691" />
                    <RANKING order="9" place="-1" resultid="3746" />
                    <RANKING order="10" place="-1" resultid="3740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7356" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2958" />
                    <RANKING order="2" place="2" resultid="4103" />
                    <RANKING order="3" place="3" resultid="2997" />
                    <RANKING order="4" place="4" resultid="5085" />
                    <RANKING order="5" place="5" resultid="1719" />
                    <RANKING order="6" place="6" resultid="2340" />
                    <RANKING order="7" place="7" resultid="3053" />
                    <RANKING order="8" place="-1" resultid="2309" />
                    <RANKING order="9" place="-1" resultid="1687" />
                    <RANKING order="10" place="-1" resultid="3028" />
                    <RANKING order="11" place="-1" resultid="1684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7357" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4238" />
                    <RANKING order="2" place="2" resultid="2879" />
                    <RANKING order="3" place="3" resultid="2833" />
                    <RANKING order="4" place="4" resultid="1753" />
                    <RANKING order="5" place="5" resultid="2347" />
                    <RANKING order="6" place="6" resultid="3734" />
                    <RANKING order="7" place="-1" resultid="2748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7358" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2588" />
                    <RANKING order="2" place="2" resultid="5677" />
                    <RANKING order="3" place="3" resultid="1804" />
                    <RANKING order="4" place="4" resultid="4093" />
                    <RANKING order="5" place="5" resultid="2061" />
                    <RANKING order="6" place="6" resultid="2611" />
                    <RANKING order="7" place="7" resultid="2516" />
                    <RANKING order="8" place="8" resultid="3947" />
                    <RANKING order="9" place="9" resultid="5045" />
                    <RANKING order="10" place="10" resultid="6424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7359" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5120" />
                    <RANKING order="2" place="2" resultid="1815" />
                    <RANKING order="3" place="3" resultid="3576" />
                    <RANKING order="4" place="4" resultid="7597" />
                    <RANKING order="5" place="5" resultid="3892" />
                    <RANKING order="6" place="6" resultid="1625" />
                    <RANKING order="7" place="7" resultid="2991" />
                    <RANKING order="8" place="-1" resultid="3086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7360" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3904" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="1702" />
                    <RANKING order="4" place="4" resultid="1744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7361" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1954" />
                    <RANKING order="2" place="2" resultid="4000" />
                    <RANKING order="3" place="3" resultid="5131" />
                    <RANKING order="4" place="4" resultid="1900" />
                    <RANKING order="5" place="5" resultid="3940" />
                    <RANKING order="6" place="6" resultid="2885" />
                    <RANKING order="7" place="7" resultid="4295" />
                    <RANKING order="8" place="-1" resultid="3690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7362" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4032" />
                    <RANKING order="2" place="2" resultid="2656" />
                    <RANKING order="3" place="3" resultid="2683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7363" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7364" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7052" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7053" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7054" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7055" daytime="16:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7056" daytime="16:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7057" daytime="16:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7058" daytime="16:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7059" daytime="16:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7060" daytime="16:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7061" daytime="16:50" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1301" daytime="16:50" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7365" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7366" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2434" />
                    <RANKING order="2" place="2" resultid="2828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7367" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3675" />
                    <RANKING order="2" place="2" resultid="4225" />
                    <RANKING order="3" place="3" resultid="2303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7368" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1792" />
                    <RANKING order="2" place="2" resultid="1672" />
                    <RANKING order="3" place="3" resultid="3011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7369" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4139" />
                    <RANKING order="2" place="2" resultid="3546" />
                    <RANKING order="3" place="3" resultid="2396" />
                    <RANKING order="4" place="4" resultid="2462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7370" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5651" />
                    <RANKING order="2" place="2" resultid="2555" />
                    <RANKING order="3" place="3" resultid="2916" />
                    <RANKING order="4" place="4" resultid="3553" />
                    <RANKING order="5" place="5" resultid="2804" />
                    <RANKING order="6" place="6" resultid="5102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7371" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="3758" />
                    <RANKING order="3" place="3" resultid="4026" />
                    <RANKING order="4" place="4" resultid="3994" />
                    <RANKING order="5" place="5" resultid="4056" />
                    <RANKING order="6" place="-1" resultid="3959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7372" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7373" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1932" />
                    <RANKING order="2" place="2" resultid="2936" />
                    <RANKING order="3" place="3" resultid="3972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7374" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/" />
                <AGEGROUP agegroupid="7375" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4934" />
                    <RANKING order="2" place="2" resultid="3809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7376" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7377" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4191" />
                    <RANKING order="2" place="2" resultid="4902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7378" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3953" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7062" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7063" daytime="16:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7064" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7065" daytime="17:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1316" daytime="17:05" gender="M" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7379" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4257" />
                    <RANKING order="2" place="2" resultid="4326" />
                    <RANKING order="3" place="3" resultid="5686" />
                    <RANKING order="4" place="4" resultid="4154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7380" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2548" />
                    <RANKING order="2" place="2" resultid="5069" />
                    <RANKING order="3" place="3" resultid="3821" />
                    <RANKING order="4" place="4" resultid="1619" />
                    <RANKING order="5" place="5" resultid="2561" />
                    <RANKING order="6" place="6" resultid="3174" />
                    <RANKING order="7" place="-1" resultid="1969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7381" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3072" />
                    <RANKING order="2" place="2" resultid="4126" />
                    <RANKING order="3" place="3" resultid="3899" />
                    <RANKING order="4" place="4" resultid="3157" />
                    <RANKING order="5" place="-1" resultid="2816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7382" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3022" />
                    <RANKING order="2" place="2" resultid="3441" />
                    <RANKING order="3" place="3" resultid="3041" />
                    <RANKING order="4" place="4" resultid="2635" />
                    <RANKING order="5" place="5" resultid="2392" />
                    <RANKING order="6" place="6" resultid="3616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7383" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1925" />
                    <RANKING order="2" place="2" resultid="2922" />
                    <RANKING order="3" place="3" resultid="3169" />
                    <RANKING order="4" place="4" resultid="2358" />
                    <RANKING order="5" place="5" resultid="4968" />
                    <RANKING order="6" place="6" resultid="2781" />
                    <RANKING order="7" place="7" resultid="4926" />
                    <RANKING order="8" place="8" resultid="3117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7384" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3046" />
                    <RANKING order="2" place="2" resultid="4826" />
                    <RANKING order="3" place="3" resultid="4219" />
                    <RANKING order="4" place="4" resultid="2823" />
                    <RANKING order="5" place="5" resultid="3496" />
                    <RANKING order="6" place="6" resultid="2576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7385" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2382" />
                    <RANKING order="2" place="2" resultid="2834" />
                    <RANKING order="3" place="3" resultid="2526" />
                    <RANKING order="4" place="4" resultid="2618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7386" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3034" />
                    <RANKING order="2" place="2" resultid="4098" />
                    <RANKING order="3" place="3" resultid="3596" />
                    <RANKING order="4" place="4" resultid="2676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7387" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2663" />
                    <RANKING order="2" place="2" resultid="3460" />
                    <RANKING order="3" place="3" resultid="4089" />
                    <RANKING order="4" place="4" resultid="2039" />
                    <RANKING order="5" place="5" resultid="3893" />
                    <RANKING order="6" place="6" resultid="4887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7388" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2953" />
                    <RANKING order="2" place="2" resultid="1943" />
                    <RANKING order="3" place="3" resultid="3059" />
                    <RANKING order="4" place="4" resultid="2364" />
                    <RANKING order="5" place="5" resultid="1745" />
                    <RANKING order="6" place="-1" resultid="1890" />
                    <RANKING order="7" place="-1" resultid="3905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7389" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1955" />
                    <RANKING order="2" place="2" resultid="3683" />
                    <RANKING order="3" place="3" resultid="2848" />
                    <RANKING order="4" place="4" resultid="4296" />
                    <RANKING order="5" place="-1" resultid="3850" />
                    <RANKING order="6" place="-1" resultid="3691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7390" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2657" />
                    <RANKING order="2" place="2" resultid="3651" />
                    <RANKING order="3" place="3" resultid="2983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7391" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3570" />
                    <RANKING order="2" place="2" resultid="3828" />
                    <RANKING order="3" place="3" resultid="2679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7392" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2898" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7066" daytime="17:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7067" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7068" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7069" daytime="17:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7070" daytime="17:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7071" daytime="17:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7072" daytime="17:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1331" daytime="17:25" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1594" agemax="119" agemin="100" name="KATEGORIA: &quot;A&quot;/100-119/" calculate="TOTAL" />
                <AGEGROUP agegroupid="1595" agemax="159" agemin="120" name="KATEGORIA: &quot;B&quot;/120-159/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7603" />
                    <RANKING order="2" place="2" resultid="2471" />
                    <RANKING order="3" place="3" resultid="7604" />
                    <RANKING order="4" place="4" resultid="7592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1596" agemax="199" agemin="160" name="KATEGORIA: &quot;C&quot;/160-199/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4864" />
                    <RANKING order="2" place="2" resultid="7610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="239" agemin="200" name="KATEGORIA: &quot;D&quot;/200-239/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2468" />
                    <RANKING order="2" place="2" resultid="7605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="279" agemin="240" name="KATEGORIA: &quot;E&quot;/240-279/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1992" />
                    <RANKING order="2" place="2" resultid="4063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="-1" agemin="280" name="KATEGORIA: &quot;F&quot;/280 i starsi/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4946" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7073" daytime="17:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7608" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1346" daytime="17:30" gender="M" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1600" agemax="119" agemin="100" name="KATEGORIA: &quot;A&quot;/100-119/" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5149" />
                    <RANKING order="2" place="2" resultid="6968" />
                    <RANKING order="3" place="3" resultid="4467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="159" agemin="120" name="KATEGORIA: &quot;B&quot;/120-159/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4352" />
                    <RANKING order="2" place="2" resultid="3800" />
                    <RANKING order="3" place="3" resultid="7600" />
                    <RANKING order="4" place="4" resultid="1993" />
                    <RANKING order="5" place="5" resultid="6969" />
                    <RANKING order="6" place="6" resultid="3926" />
                    <RANKING order="7" place="7" resultid="7599" />
                    <RANKING order="8" place="8" resultid="3514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="199" agemin="160" name="KATEGORIA: &quot;C&quot;/160-199/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4985" />
                    <RANKING order="2" place="2" resultid="2466" />
                    <RANKING order="3" place="3" resultid="7601" />
                    <RANKING order="4" place="4" resultid="7595" />
                    <RANKING order="5" place="-1" resultid="2836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="239" agemin="200" name="KATEGORIA: &quot;D&quot;/200-239/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7607" />
                    <RANKING order="2" place="2" resultid="3515" />
                    <RANKING order="3" place="3" resultid="7602" />
                    <RANKING order="4" place="-1" resultid="3716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="279" agemin="240" name="KATEGORIA: &quot;E&quot;/240-279/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1994" />
                    <RANKING order="2" place="2" resultid="1839" />
                    <RANKING order="3" place="3" resultid="7177" />
                    <RANKING order="4" place="4" resultid="2476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="-1" agemin="280" name="KATEGORIA: &quot;F&quot;/280 i starsi/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7606" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7074" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7075" daytime="17:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7076" daytime="17:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1361" daytime="17:40" gender="F" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7393" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="3857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7394" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3638" />
                    <RANKING order="2" place="2" resultid="1738" />
                    <RANKING order="3" place="3" resultid="5143" />
                    <RANKING order="4" place="4" resultid="3667" />
                    <RANKING order="5" place="5" resultid="1650" />
                    <RANKING order="6" place="-1" resultid="3815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7395" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3419" />
                    <RANKING order="2" place="2" resultid="2571" />
                    <RANKING order="3" place="3" resultid="4226" />
                    <RANKING order="4" place="4" resultid="3110" />
                    <RANKING order="5" place="5" resultid="2281" />
                    <RANKING order="6" place="6" resultid="3206" />
                    <RANKING order="7" place="7" resultid="4130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7396" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1614" />
                    <RANKING order="2" place="2" resultid="2628" />
                    <RANKING order="3" place="3" resultid="3012" />
                    <RANKING order="4" place="4" resultid="2439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7397" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3198" />
                    <RANKING order="2" place="2" resultid="2397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7398" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2869" />
                    <RANKING order="2" place="2" resultid="2556" />
                    <RANKING order="3" place="3" resultid="3195" />
                    <RANKING order="4" place="4" resultid="2917" />
                    <RANKING order="5" place="5" resultid="4819" />
                    <RANKING order="6" place="6" resultid="5103" />
                    <RANKING order="7" place="-1" resultid="5110" />
                    <RANKING order="8" place="-1" resultid="2805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7399" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4115" />
                    <RANKING order="2" place="2" resultid="1828" />
                    <RANKING order="3" place="3" resultid="1821" />
                    <RANKING order="4" place="4" resultid="2582" />
                    <RANKING order="5" place="5" resultid="1644" />
                    <RANKING order="6" place="6" resultid="2605" />
                    <RANKING order="7" place="7" resultid="1676" />
                    <RANKING order="8" place="8" resultid="4918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7400" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7401" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2776" />
                    <RANKING order="2" place="2" resultid="1939" />
                    <RANKING order="3" place="3" resultid="3218" />
                    <RANKING order="4" place="4" resultid="3007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7402" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3182" />
                    <RANKING order="2" place="2" resultid="2909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7403" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/" />
                <AGEGROUP agegroupid="7404" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7405" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7406" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7077" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7078" daytime="17:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7079" daytime="17:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7080" daytime="17:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7081" daytime="17:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1376" daytime="18:00" gender="M" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7407" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5038" />
                    <RANKING order="2" place="2" resultid="3763" />
                    <RANKING order="3" place="3" resultid="2334" />
                    <RANKING order="4" place="4" resultid="3138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7408" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4202" />
                    <RANKING order="2" place="2" resultid="3151" />
                    <RANKING order="3" place="3" resultid="4232" />
                    <RANKING order="4" place="4" resultid="4317" />
                    <RANKING order="5" place="5" resultid="4185" />
                    <RANKING order="6" place="6" resultid="4251" />
                    <RANKING order="7" place="7" resultid="3175" />
                    <RANKING order="8" place="8" resultid="1778" />
                    <RANKING order="9" place="9" resultid="1869" />
                    <RANKING order="10" place="10" resultid="2874" />
                    <RANKING order="11" place="-1" resultid="1620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7409" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3878" />
                    <RANKING order="2" place="2" resultid="1863" />
                    <RANKING order="3" place="3" resultid="3845" />
                    <RANKING order="4" place="4" resultid="3865" />
                    <RANKING order="5" place="5" resultid="1875" />
                    <RANKING order="6" place="6" resultid="5493" />
                    <RANKING order="7" place="7" resultid="5655" />
                    <RANKING order="8" place="-1" resultid="3539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7410" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3447" />
                    <RANKING order="2" place="2" resultid="3768" />
                    <RANKING order="3" place="3" resultid="2865" />
                    <RANKING order="4" place="4" resultid="3475" />
                    <RANKING order="5" place="5" resultid="3751" />
                    <RANKING order="6" place="6" resultid="2046" />
                    <RANKING order="7" place="7" resultid="3737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7411" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3126" />
                    <RANKING order="2" place="2" resultid="1926" />
                    <RANKING order="3" place="3" resultid="4962" />
                    <RANKING order="4" place="4" resultid="3433" />
                    <RANKING order="5" place="5" resultid="2509" />
                    <RANKING order="6" place="6" resultid="5128" />
                    <RANKING order="7" place="7" resultid="4927" />
                    <RANKING order="8" place="8" resultid="3118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7412" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3643" />
                    <RANKING order="2" place="2" resultid="3047" />
                    <RANKING order="3" place="3" resultid="4286" />
                    <RANKING order="4" place="4" resultid="4220" />
                    <RANKING order="5" place="5" resultid="4104" />
                    <RANKING order="6" place="6" resultid="2577" />
                    <RANKING order="7" place="7" resultid="3016" />
                    <RANKING order="8" place="-1" resultid="2797" />
                    <RANKING order="9" place="-1" resultid="1655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7413" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3067" />
                    <RANKING order="2" place="2" resultid="4829" />
                    <RANKING order="3" place="3" resultid="2810" />
                    <RANKING order="4" place="4" resultid="1787" />
                    <RANKING order="5" place="5" resultid="1712" />
                    <RANKING order="6" place="6" resultid="4239" />
                    <RANKING order="7" place="7" resultid="2932" />
                    <RANKING order="8" place="8" resultid="4892" />
                    <RANKING order="9" place="9" resultid="3145" />
                    <RANKING order="10" place="-1" resultid="6420" />
                    <RANKING order="11" place="-1" resultid="3467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7414" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1782" />
                    <RANKING order="2" place="2" resultid="4121" />
                    <RANKING order="3" place="3" resultid="1895" />
                    <RANKING order="4" place="4" resultid="4170" />
                    <RANKING order="5" place="5" resultid="4882" />
                    <RANKING order="6" place="6" resultid="2612" />
                    <RANKING order="7" place="7" resultid="3797" />
                    <RANKING order="8" place="-1" resultid="3698" />
                    <RANKING order="9" place="-1" resultid="1799" />
                    <RANKING order="10" place="-1" resultid="2053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7415" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4837" />
                    <RANKING order="2" place="2" resultid="2664" />
                    <RANKING order="3" place="3" resultid="3577" />
                    <RANKING order="4" place="4" resultid="3711" />
                    <RANKING order="5" place="5" resultid="1852" />
                    <RANKING order="6" place="-1" resultid="4177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7416" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2375" />
                    <RANKING order="2" place="2" resultid="2954" />
                    <RANKING order="3" place="3" resultid="3060" />
                    <RANKING order="4" place="-1" resultid="2902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7417" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7418" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                    <RANKING order="2" place="2" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7419" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3660" />
                    <RANKING order="2" place="2" resultid="3829" />
                    <RANKING order="3" place="3" resultid="2680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7420" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7082" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7083" daytime="18:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7084" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7085" daytime="18:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7086" daytime="18:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7087" daytime="18:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7088" daytime="18:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7089" daytime="18:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7090" daytime="18:30" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1391" daytime="18:35" gender="F" number="21" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7421" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4144" />
                    <RANKING order="2" place="2" resultid="1769" />
                    <RANKING order="3" place="3" resultid="3858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7422" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3238" />
                    <RANKING order="2" place="2" resultid="3104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7423" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4267" />
                    <RANKING order="2" place="2" resultid="3093" />
                    <RANKING order="3" place="3" resultid="4131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7424" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                    <RANKING order="2" place="2" resultid="4014" />
                    <RANKING order="3" place="-1" resultid="4851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7425" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1916" />
                    <RANKING order="2" place="2" resultid="3547" />
                    <RANKING order="3" place="3" resultid="2398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7426" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3839" />
                    <RANKING order="2" place="2" resultid="2444" />
                    <RANKING order="3" place="3" resultid="3489" />
                    <RANKING order="4" place="4" resultid="4820" />
                    <RANKING order="5" place="5" resultid="3554" />
                    <RANKING order="6" place="6" resultid="2948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7427" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5650" />
                    <RANKING order="2" place="2" resultid="2268" />
                    <RANKING order="3" place="3" resultid="1645" />
                    <RANKING order="4" place="4" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7428" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4085" />
                    <RANKING order="2" place="2" resultid="2421" />
                    <RANKING order="3" place="3" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7429" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4079" />
                    <RANKING order="2" place="2" resultid="2404" />
                    <RANKING order="3" place="3" resultid="4020" />
                    <RANKING order="4" place="-1" resultid="4897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7430" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3984" />
                    <RANKING order="2" place="2" resultid="2428" />
                    <RANKING order="3" place="3" resultid="4944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7431" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/" />
                <AGEGROUP agegroupid="7432" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7433" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7434" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7091" daytime="18:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7092" daytime="18:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7093" daytime="18:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7094" daytime="18:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="18:55" gender="M" number="22" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7435" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2324" />
                    <RANKING order="2" place="2" resultid="3562" />
                    <RANKING order="3" place="3" resultid="3764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7436" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1970" />
                    <RANKING order="2" place="2" resultid="3792" />
                    <RANKING order="3" place="3" resultid="4150" />
                    <RANKING order="4" place="4" resultid="4252" />
                    <RANKING order="5" place="5" resultid="3079" />
                    <RANKING order="6" place="6" resultid="4147" />
                    <RANKING order="7" place="7" resultid="5587" />
                    <RANKING order="8" place="8" resultid="2755" />
                    <RANKING order="9" place="-1" resultid="6963" />
                    <RANKING order="10" place="-1" resultid="4303" />
                    <RANKING order="11" place="-1" resultid="3822" />
                    <RANKING order="12" place="-1" resultid="5094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7437" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2941" />
                    <RANKING order="2" place="2" resultid="3879" />
                    <RANKING order="3" place="3" resultid="3073" />
                    <RANKING order="4" place="4" resultid="1964" />
                    <RANKING order="5" place="5" resultid="3454" />
                    <RANKING order="6" place="-1" resultid="2817" />
                    <RANKING order="7" place="-1" resultid="2959" />
                    <RANKING order="8" place="-1" resultid="3886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7438" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3502" />
                    <RANKING order="2" place="2" resultid="5491" />
                    <RANKING order="3" place="3" resultid="4975" />
                    <RANKING order="4" place="4" resultid="3482" />
                    <RANKING order="5" place="5" resultid="3164" />
                    <RANKING order="6" place="6" resultid="2566" />
                    <RANKING order="7" place="7" resultid="2047" />
                    <RANKING order="8" place="8" resultid="3752" />
                    <RANKING order="9" place="9" resultid="3617" />
                    <RANKING order="10" place="-1" resultid="3509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7439" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="4963" />
                    <RANKING order="3" place="3" resultid="3729" />
                    <RANKING order="4" place="4" resultid="3434" />
                    <RANKING order="5" place="5" resultid="4969" />
                    <RANKING order="6" place="6" resultid="4981" />
                    <RANKING order="7" place="7" resultid="3119" />
                    <RANKING order="8" place="-1" resultid="5050" />
                    <RANKING order="9" place="-1" resultid="2359" />
                    <RANKING order="10" place="-1" resultid="1692" />
                    <RANKING order="11" place="-1" resultid="3784" />
                    <RANKING order="12" place="-1" resultid="3170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7440" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3644" />
                    <RANKING order="2" place="2" resultid="1637" />
                    <RANKING order="3" place="3" resultid="2977" />
                    <RANKING order="4" place="4" resultid="2594" />
                    <RANKING order="5" place="5" resultid="2998" />
                    <RANKING order="6" place="6" resultid="3705" />
                    <RANKING order="7" place="7" resultid="2341" />
                    <RANKING order="8" place="-1" resultid="2310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7441" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2889" />
                    <RANKING order="2" place="2" resultid="2880" />
                    <RANKING order="3" place="3" resultid="2856" />
                    <RANKING order="4" place="4" resultid="3468" />
                    <RANKING order="5" place="5" resultid="2348" />
                    <RANKING order="6" place="6" resultid="3777" />
                    <RANKING order="7" place="-1" resultid="1713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7442" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3035" />
                    <RANKING order="2" place="2" resultid="5678" />
                    <RANKING order="3" place="3" resultid="4094" />
                    <RANKING order="4" place="4" resultid="4883" />
                    <RANKING order="5" place="-1" resultid="2062" />
                    <RANKING order="6" place="-1" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7443" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5121" />
                    <RANKING order="2" place="2" resultid="1680" />
                    <RANKING order="3" place="3" resultid="3872" />
                    <RANKING order="4" place="4" resultid="4245" />
                    <RANKING order="5" place="5" resultid="3461" />
                    <RANKING order="6" place="6" resultid="2040" />
                    <RANKING order="7" place="7" resultid="3712" />
                    <RANKING order="8" place="8" resultid="2670" />
                    <RANKING order="9" place="9" resultid="4888" />
                    <RANKING order="10" place="-1" resultid="4008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7444" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2690" />
                    <RANKING order="2" place="2" resultid="2376" />
                    <RANKING order="3" place="3" resultid="2787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7445" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4001" />
                    <RANKING order="2" place="2" resultid="3684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7446" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7447" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7448" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7095" daytime="18:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7096" daytime="19:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7097" daytime="19:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7098" daytime="19:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7099" daytime="19:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7100" daytime="19:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7101" daytime="19:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7102" daytime="19:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7103" daytime="19:25" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2012-05-27" daytime="09:00" name="III BLOK" number="3" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="1422" daytime="09:00" gender="F" number="23" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7449" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/" />
                <AGEGROUP agegroupid="7450" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3603" />
                    <RANKING order="2" place="2" resultid="3105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7451" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3420" />
                    <RANKING order="2" place="2" resultid="2304" />
                    <RANKING order="3" place="3" resultid="2623" />
                    <RANKING order="4" place="4" resultid="2282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7452" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4852" />
                    <RANKING order="2" place="2" resultid="2440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7453" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/" />
                <AGEGROUP agegroupid="7454" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3840" />
                    <RANKING order="2" place="2" resultid="2445" />
                    <RANKING order="3" place="3" resultid="2949" />
                    <RANKING order="4" place="4" resultid="3555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7455" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1822" />
                    <RANKING order="2" place="2" resultid="4039" />
                    <RANKING order="3" place="3" resultid="1646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7456" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2422" />
                    <RANKING order="2" place="2" resultid="4051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7457" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4021" />
                    <RANKING order="2" place="-1" resultid="4898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7458" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7459" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/" />
                <AGEGROUP agegroupid="7460" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7461" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7462" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7104" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7105" daytime="09:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1438" daytime="09:05" gender="M" number="24" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7463" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3563" />
                    <RANKING order="2" place="2" resultid="3765" />
                    <RANKING order="3" place="-1" resultid="5064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7464" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2549" />
                    <RANKING order="2" place="2" resultid="5071" />
                    <RANKING order="3" place="3" resultid="4203" />
                    <RANKING order="4" place="4" resultid="5032" />
                    <RANKING order="5" place="5" resultid="3773" />
                    <RANKING order="6" place="6" resultid="4151" />
                    <RANKING order="7" place="7" resultid="5588" />
                    <RANKING order="8" place="8" resultid="4186" />
                    <RANKING order="9" place="9" resultid="1870" />
                    <RANKING order="10" place="-1" resultid="4148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7465" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1965" />
                    <RANKING order="2" place="2" resultid="1876" />
                    <RANKING order="3" place="3" resultid="3455" />
                    <RANKING order="4" place="-1" resultid="3887" />
                    <RANKING order="5" place="-1" resultid="3540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7466" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3023" />
                    <RANKING order="2" place="2" resultid="3448" />
                    <RANKING order="3" place="3" resultid="2388" />
                    <RANKING order="4" place="4" resultid="3503" />
                    <RANKING order="5" place="5" resultid="4976" />
                    <RANKING order="6" place="6" resultid="3165" />
                    <RANKING order="7" place="7" resultid="4515" />
                    <RANKING order="8" place="8" resultid="3510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7467" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3127" />
                    <RANKING order="2" place="2" resultid="1735" />
                    <RANKING order="3" place="3" resultid="3730" />
                    <RANKING order="4" place="4" resultid="2894" />
                    <RANKING order="5" place="5" resultid="5051" />
                    <RANKING order="6" place="-1" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7468" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                    <RANKING order="2" place="2" resultid="2595" />
                    <RANKING order="3" place="3" resultid="2978" />
                    <RANKING order="4" place="4" resultid="3497" />
                    <RANKING order="5" place="5" resultid="2798" />
                    <RANKING order="6" place="-1" resultid="3029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7469" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4830" />
                    <RANKING order="2" place="2" resultid="2890" />
                    <RANKING order="3" place="3" resultid="2857" />
                    <RANKING order="4" place="-1" resultid="2383" />
                    <RANKING order="5" place="-1" resultid="3469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7470" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1800" />
                    <RANKING order="2" place="2" resultid="5679" />
                    <RANKING order="3" place="3" resultid="4122" />
                    <RANKING order="4" place="4" resultid="2517" />
                    <RANKING order="5" place="-1" resultid="1806" />
                    <RANKING order="6" place="-1" resultid="3699" />
                    <RANKING order="7" place="-1" resultid="6693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7471" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4246" />
                    <RANKING order="2" place="2" resultid="3873" />
                    <RANKING order="3" place="3" resultid="4838" />
                    <RANKING order="4" place="4" resultid="5122" />
                    <RANKING order="5" place="5" resultid="3894" />
                    <RANKING order="6" place="6" resultid="2671" />
                    <RANKING order="7" place="7" resultid="3713" />
                    <RANKING order="8" place="8" resultid="2041" />
                    <RANKING order="9" place="9" resultid="1853" />
                    <RANKING order="10" place="10" resultid="4889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7472" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="1811" />
                    <RANKING order="3" place="3" resultid="2377" />
                    <RANKING order="4" place="4" resultid="6417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7473" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7474" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7475" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7476" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7106" daytime="09:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7107" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7108" daytime="09:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7109" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7110" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7111" daytime="09:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7112" daytime="09:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1453" daytime="09:20" gender="F" number="25" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7477" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7618" />
                    <RANKING order="2" place="2" resultid="1770" />
                    <RANKING order="3" place="3" resultid="1762" />
                    <RANKING order="4" place="4" resultid="4061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7478" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5060" />
                    <RANKING order="2" place="2" resultid="3604" />
                    <RANKING order="3" place="3" resultid="3639" />
                    <RANKING order="4" place="4" resultid="5487" />
                    <RANKING order="5" place="5" resultid="4165" />
                    <RANKING order="6" place="6" resultid="4844" />
                    <RANKING order="7" place="7" resultid="5144" />
                    <RANKING order="8" place="8" resultid="3668" />
                    <RANKING order="9" place="-1" resultid="3816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7479" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3421" />
                    <RANKING order="2" place="2" resultid="4268" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="3111" />
                    <RANKING order="5" place="5" resultid="4132" />
                    <RANKING order="6" place="6" resultid="3207" />
                    <RANKING order="7" place="7" resultid="3094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7480" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3132" />
                    <RANKING order="2" place="2" resultid="4291" />
                    <RANKING order="3" place="3" resultid="3088" />
                    <RANKING order="4" place="4" resultid="3916" />
                    <RANKING order="5" place="5" resultid="2629" />
                    <RANKING order="6" place="6" resultid="2926" />
                    <RANKING order="7" place="7" resultid="2929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7481" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="3199" />
                    <RANKING order="3" place="3" resultid="5137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7482" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2411" />
                    <RANKING order="2" place="2" resultid="2557" />
                    <RANKING order="3" place="3" resultid="3490" />
                    <RANKING order="4" place="4" resultid="4821" />
                    <RANKING order="5" place="5" resultid="5111" />
                    <RANKING order="6" place="6" resultid="5104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7483" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1829" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="3" resultid="2457" />
                    <RANKING order="4" place="4" resultid="2606" />
                    <RANKING order="5" place="5" resultid="2451" />
                    <RANKING order="6" place="6" resultid="3995" />
                    <RANKING order="7" place="7" resultid="2269" />
                    <RANKING order="8" place="8" resultid="2275" />
                    <RANKING order="9" place="9" resultid="4044" />
                    <RANKING order="10" place="10" resultid="3960" />
                    <RANKING order="11" place="-1" resultid="2583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7484" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1662" />
                    <RANKING order="2" place="2" resultid="1836" />
                    <RANKING order="3" place="3" resultid="5116" />
                    <RANKING order="4" place="4" resultid="3601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7485" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4080" />
                    <RANKING order="2" place="2" resultid="2777" />
                    <RANKING order="3" place="3" resultid="1940" />
                    <RANKING order="4" place="4" resultid="1665" />
                    <RANKING order="5" place="5" resultid="3219" />
                    <RANKING order="6" place="6" resultid="3973" />
                    <RANKING order="7" place="-1" resultid="4899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7486" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1961" />
                    <RANKING order="2" place="2" resultid="4847" />
                    <RANKING order="3" place="3" resultid="3989" />
                    <RANKING order="4" place="4" resultid="1980" />
                    <RANKING order="5" place="5" resultid="3183" />
                    <RANKING order="6" place="6" resultid="2910" />
                    <RANKING order="7" place="7" resultid="3985" />
                    <RANKING order="8" place="8" resultid="2429" />
                    <RANKING order="9" place="9" resultid="4215" />
                    <RANKING order="10" place="10" resultid="2913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7487" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7488" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7489" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4192" />
                    <RANKING order="2" place="-1" resultid="4906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7490" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3954" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7113" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7114" daytime="09:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7115" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7116" daytime="09:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7117" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7118" daytime="09:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7119" daytime="09:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7120" daytime="09:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1468" daytime="09:35" gender="M" number="26" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7491" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2335" />
                    <RANKING order="2" place="2" resultid="3139" />
                    <RANKING order="3" place="3" resultid="4258" />
                    <RANKING order="4" place="4" resultid="3923" />
                    <RANKING order="5" place="5" resultid="4327" />
                    <RANKING order="6" place="6" resultid="4155" />
                    <RANKING order="7" place="-1" resultid="5065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7492" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3672" />
                    <RANKING order="2" place="2" resultid="2550" />
                    <RANKING order="3" place="3" resultid="1859" />
                    <RANKING order="4" place="4" resultid="2297" />
                    <RANKING order="5" place="5" resultid="4308" />
                    <RANKING order="6" place="6" resultid="1779" />
                    <RANKING order="7" place="7" resultid="5078" />
                    <RANKING order="8" place="8" resultid="3774" />
                    <RANKING order="9" place="9" resultid="3152" />
                    <RANKING order="10" place="10" resultid="4233" />
                    <RANKING order="11" place="11" resultid="3176" />
                    <RANKING order="12" place="12" resultid="3788" />
                    <RANKING order="13" place="13" resultid="5475" />
                    <RANKING order="14" place="14" resultid="4318" />
                    <RANKING order="15" place="15" resultid="1988" />
                    <RANKING order="16" place="16" resultid="4136" />
                    <RANKING order="17" place="17" resultid="4322" />
                    <RANKING order="18" place="18" resultid="5058" />
                    <RANKING order="19" place="19" resultid="3584" />
                    <RANKING order="20" place="20" resultid="1871" />
                    <RANKING order="21" place="21" resultid="4262" />
                    <RANKING order="22" place="22" resultid="3620" />
                    <RANKING order="23" place="23" resultid="2875" />
                    <RANKING order="24" place="-1" resultid="1631" />
                    <RANKING order="25" place="-1" resultid="3793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7493" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1864" />
                    <RANKING order="2" place="2" resultid="4210" />
                    <RANKING order="3" place="3" resultid="3121" />
                    <RANKING order="4" place="4" resultid="2988" />
                    <RANKING order="5" place="5" resultid="2942" />
                    <RANKING order="6" place="6" resultid="5035" />
                    <RANKING order="7" place="7" resultid="5054" />
                    <RANKING order="8" place="8" resultid="3846" />
                    <RANKING order="9" place="9" resultid="3866" />
                    <RANKING order="10" place="10" resultid="5041" />
                    <RANKING order="11" place="11" resultid="1877" />
                    <RANKING order="12" place="12" resultid="3541" />
                    <RANKING order="13" place="13" resultid="2975" />
                    <RANKING order="14" place="14" resultid="4855" />
                    <RANKING order="15" place="15" resultid="3159" />
                    <RANKING order="16" place="16" resultid="5656" />
                    <RANKING order="17" place="17" resultid="5043" />
                    <RANKING order="18" place="18" resultid="3624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7494" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                    <RANKING order="2" place="2" resultid="3042" />
                    <RANKING order="3" place="3" resultid="2636" />
                    <RANKING order="4" place="4" resultid="4861" />
                    <RANKING order="5" place="5" resultid="3613" />
                    <RANKING order="6" place="6" resultid="3753" />
                    <RANKING order="7" place="7" resultid="2567" />
                    <RANKING order="8" place="8" resultid="1710" />
                    <RANKING order="9" place="9" resultid="5075" />
                    <RANKING order="10" place="-1" resultid="3632" />
                    <RANKING order="11" place="-1" resultid="2945" />
                    <RANKING order="12" place="-1" resultid="7594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7495" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3785" />
                    <RANKING order="2" place="2" resultid="1736" />
                    <RANKING order="3" place="3" resultid="3435" />
                    <RANKING order="4" place="4" resultid="2360" />
                    <RANKING order="5" place="5" resultid="4964" />
                    <RANKING order="6" place="6" resultid="4970" />
                    <RANKING order="7" place="7" resultid="3833" />
                    <RANKING order="8" place="8" resultid="5129" />
                    <RANKING order="9" place="9" resultid="4982" />
                    <RANKING order="10" place="10" resultid="1705" />
                    <RANKING order="11" place="11" resultid="3188" />
                    <RANKING order="12" place="12" resultid="5052" />
                    <RANKING order="13" place="13" resultid="4928" />
                    <RANKING order="14" place="14" resultid="3747" />
                    <RANKING order="15" place="-1" resultid="3214" />
                    <RANKING order="16" place="-1" resultid="1976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7496" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3645" />
                    <RANKING order="2" place="2" resultid="2596" />
                    <RANKING order="3" place="3" resultid="1639" />
                    <RANKING order="4" place="4" resultid="4287" />
                    <RANKING order="5" place="5" resultid="2824" />
                    <RANKING order="6" place="6" resultid="2999" />
                    <RANKING order="7" place="7" resultid="3706" />
                    <RANKING order="8" place="8" resultid="2342" />
                    <RANKING order="9" place="9" resultid="2578" />
                    <RANKING order="10" place="10" resultid="3054" />
                    <RANKING order="11" place="11" resultid="3017" />
                    <RANKING order="12" place="-1" resultid="1656" />
                    <RANKING order="13" place="-1" resultid="1685" />
                    <RANKING order="14" place="-1" resultid="5134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7497" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3068" />
                    <RANKING order="2" place="2" resultid="2811" />
                    <RANKING order="3" place="3" resultid="2881" />
                    <RANKING order="4" place="4" resultid="1714" />
                    <RANKING order="5" place="5" resultid="2933" />
                    <RANKING order="6" place="6" resultid="3004" />
                    <RANKING order="7" place="7" resultid="1754" />
                    <RANKING order="8" place="8" resultid="3778" />
                    <RANKING order="9" place="9" resultid="3146" />
                    <RANKING order="10" place="10" resultid="3735" />
                    <RANKING order="11" place="-1" resultid="6421" />
                    <RANKING order="12" place="-1" resultid="1727" />
                    <RANKING order="13" place="-1" resultid="2527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7498" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1783" />
                    <RANKING order="2" place="2" resultid="1730" />
                    <RANKING order="3" place="3" resultid="1896" />
                    <RANKING order="4" place="4" resultid="2677" />
                    <RANKING order="5" place="5" resultid="4171" />
                    <RANKING order="6" place="6" resultid="4911" />
                    <RANKING order="7" place="7" resultid="3597" />
                    <RANKING order="8" place="8" resultid="2589" />
                    <RANKING order="9" place="9" resultid="4099" />
                    <RANKING order="10" place="10" resultid="1724" />
                    <RANKING order="11" place="11" resultid="7619" />
                    <RANKING order="12" place="12" resultid="2613" />
                    <RANKING order="13" place="13" resultid="3948" />
                    <RANKING order="14" place="14" resultid="6425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7499" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2665" />
                    <RANKING order="2" place="2" resultid="4839" />
                    <RANKING order="3" place="3" resultid="1681" />
                    <RANKING order="4" place="4" resultid="3874" />
                    <RANKING order="5" place="5" resultid="3462" />
                    <RANKING order="6" place="6" resultid="1911" />
                    <RANKING order="7" place="7" resultid="4247" />
                    <RANKING order="8" place="8" resultid="1936" />
                    <RANKING order="9" place="9" resultid="5499" />
                    <RANKING order="10" place="10" resultid="4009" />
                    <RANKING order="11" place="11" resultid="3578" />
                    <RANKING order="12" place="12" resultid="1699" />
                    <RANKING order="13" place="13" resultid="1984" />
                    <RANKING order="14" place="14" resultid="7620" />
                    <RANKING order="15" place="15" resultid="1626" />
                    <RANKING order="16" place="16" resultid="2992" />
                    <RANKING order="17" place="-1" resultid="4178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7500" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="2955" />
                    <RANKING order="3" place="3" resultid="1812" />
                    <RANKING order="4" place="4" resultid="3061" />
                    <RANKING order="5" place="5" resultid="2903" />
                    <RANKING order="6" place="6" resultid="2365" />
                    <RANKING order="7" place="7" resultid="5583" />
                    <RANKING order="8" place="8" resultid="1746" />
                    <RANKING order="9" place="9" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7501" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1956" />
                    <RANKING order="2" place="2" resultid="2886" />
                    <RANKING order="3" place="3" resultid="4002" />
                    <RANKING order="4" place="4" resultid="5132" />
                    <RANKING order="5" place="5" resultid="3038" />
                    <RANKING order="6" place="6" resultid="3852" />
                    <RANKING order="7" place="-1" resultid="3692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7502" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2658" />
                    <RANKING order="2" place="2" resultid="2330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7503" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3662" />
                    <RANKING order="2" place="2" resultid="3830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7504" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2899" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7121" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7122" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7123" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7124" daytime="09:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7125" daytime="09:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7126" daytime="09:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7127" daytime="09:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7128" daytime="09:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7129" daytime="09:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7130" daytime="09:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7131" daytime="09:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7132" daytime="09:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7133" daytime="09:50" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7134" daytime="09:55" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7135" daytime="09:55" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7136" daytime="09:55" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1483" daytime="09:55" gender="F" number="27" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7505" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7506" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2435" />
                    <RANKING order="2" place="2" resultid="2829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7507" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4227" />
                    <RANKING order="2" place="2" resultid="2305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7508" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3089" />
                    <RANKING order="2" place="2" resultid="1794" />
                    <RANKING order="3" place="3" resultid="3013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7509" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3549" />
                    <RANKING order="2" place="2" resultid="2399" />
                    <RANKING order="3" place="3" resultid="2463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7510" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2918" />
                    <RANKING order="2" place="2" resultid="2558" />
                    <RANKING order="3" place="3" resultid="3556" />
                    <RANKING order="4" place="4" resultid="5105" />
                    <RANKING order="5" place="-1" resultid="2806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7511" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4116" />
                    <RANKING order="2" place="2" resultid="3759" />
                    <RANKING order="3" place="3" resultid="4028" />
                    <RANKING order="4" place="4" resultid="3996" />
                    <RANKING order="5" place="5" resultid="4057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7512" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2423" />
                    <RANKING order="2" place="2" resultid="3966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7513" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1933" />
                    <RANKING order="2" place="2" resultid="2937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7514" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7515" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7516" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7517" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7518" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7137" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7138" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7139" daytime="10:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1498" daytime="10:10" gender="M" number="28" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7519" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5687" />
                    <RANKING order="2" place="-1" resultid="4328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7520" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5492" />
                    <RANKING order="2" place="2" resultid="1971" />
                    <RANKING order="3" place="3" resultid="1621" />
                    <RANKING order="4" place="4" resultid="2562" />
                    <RANKING order="5" place="5" resultid="3177" />
                    <RANKING order="6" place="6" resultid="4323" />
                    <RANKING order="7" place="-1" resultid="2756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7521" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3074" />
                    <RANKING order="2" place="2" resultid="3880" />
                    <RANKING order="3" place="3" resultid="1966" />
                    <RANKING order="4" place="4" resultid="3900" />
                    <RANKING order="5" place="-1" resultid="2818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7522" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3443" />
                    <RANKING order="2" place="2" resultid="2637" />
                    <RANKING order="3" place="3" resultid="3483" />
                    <RANKING order="4" place="-1" resultid="2048" />
                    <RANKING order="5" place="-1" resultid="3043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7523" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1927" />
                    <RANKING order="2" place="2" resultid="2923" />
                    <RANKING order="3" place="3" resultid="3128" />
                    <RANKING order="4" place="4" resultid="2782" />
                    <RANKING order="5" place="5" resultid="4929" />
                    <RANKING order="6" place="-1" resultid="2510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7524" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2597" />
                    <RANKING order="2" place="2" resultid="4221" />
                    <RANKING order="3" place="3" resultid="2825" />
                    <RANKING order="4" place="4" resultid="3498" />
                    <RANKING order="5" place="5" resultid="2579" />
                    <RANKING order="6" place="6" resultid="2799" />
                    <RANKING order="7" place="-1" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7525" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2384" />
                    <RANKING order="2" place="2" resultid="3470" />
                    <RANKING order="3" place="3" resultid="2619" />
                    <RANKING order="4" place="4" resultid="2528" />
                    <RANKING order="5" place="5" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7526" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3036" />
                    <RANKING order="2" place="2" resultid="4095" />
                    <RANKING order="3" place="3" resultid="3598" />
                    <RANKING order="4" place="-1" resultid="2063" />
                    <RANKING order="5" place="-1" resultid="2055" />
                    <RANKING order="6" place="-1" resultid="4100" />
                    <RANKING order="7" place="-1" resultid="3700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7527" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2666" />
                    <RANKING order="2" place="2" resultid="3463" />
                    <RANKING order="3" place="3" resultid="4090" />
                    <RANKING order="4" place="4" resultid="2042" />
                    <RANKING order="5" place="5" resultid="4890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7528" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2956" />
                    <RANKING order="2" place="2" resultid="1944" />
                    <RANKING order="3" place="3" resultid="2788" />
                    <RANKING order="4" place="-1" resultid="2366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7529" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3685" />
                    <RANKING order="2" place="2" resultid="2849" />
                    <RANKING order="3" place="3" resultid="4297" />
                    <RANKING order="4" place="4" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7530" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2659" />
                    <RANKING order="2" place="2" resultid="2985" />
                    <RANKING order="3" place="3" resultid="3653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7531" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3571" />
                    <RANKING order="2" place="2" resultid="3831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7532" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7140" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7141" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7142" daytime="10:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7143" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7144" daytime="10:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7145" daytime="10:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7146" daytime="10:40" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1513" daytime="10:45" gender="X" number="29" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1606" agemax="119" agemin="100" name="KATEGORIA: &quot;A&quot;/100-119/" calculate="TOTAL" />
                <AGEGROUP agegroupid="1607" agemax="159" agemin="120" name="KATEGORIA: &quot;B&quot;/120-159/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="7612" />
                    <RANKING order="3" place="3" resultid="7613" />
                    <RANKING order="4" place="4" resultid="2475" />
                    <RANKING order="5" place="5" resultid="7615" />
                    <RANKING order="6" place="6" resultid="3627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="199" agemin="160" name="KATEGORIA: &quot;C&quot;/160-199/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2473" />
                    <RANKING order="2" place="2" resultid="4863" />
                    <RANKING order="3" place="3" resultid="7617" />
                    <RANKING order="4" place="4" resultid="7622" />
                    <RANKING order="5" place="5" resultid="7614" />
                    <RANKING order="6" place="6" resultid="2838" />
                    <RANKING order="7" place="7" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="239" agemin="200" name="KATEGORIA: &quot;D&quot;/200-239/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="1840" />
                    <RANKING order="3" place="3" resultid="7623" />
                    <RANKING order="4" place="4" resultid="7621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1610" agemax="279" agemin="240" name="KATEGORIA: &quot;E&quot;/240-279/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2465" />
                    <RANKING order="2" place="2" resultid="3976" />
                    <RANKING order="3" place="-1" resultid="7616" />
                    <RANKING order="4" place="-1" resultid="1995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1611" agemax="-1" agemin="280" name="KATEGORIA: &quot;F&quot;/280 i starsi/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1996" />
                    <RANKING order="2" place="2" resultid="4062" />
                    <RANKING order="3" place="3" resultid="4947" />
                    <RANKING order="4" place="-1" resultid="3283" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7147" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7148" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7149" daytime="10:55" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1528" daytime="11:00" gender="F" number="30" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7533" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4145" />
                    <RANKING order="2" place="-1" resultid="1771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7534" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5159" />
                    <RANKING order="2" place="2" resultid="3239" />
                    <RANKING order="3" place="3" resultid="2416" />
                    <RANKING order="4" place="4" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7535" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3535" />
                    <RANKING order="2" place="2" resultid="3112" />
                    <RANKING order="3" place="3" resultid="3622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7536" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3133" />
                    <RANKING order="2" place="2" resultid="3917" />
                    <RANKING order="3" place="3" resultid="1673" />
                    <RANKING order="4" place="4" resultid="4015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7537" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1917" />
                    <RANKING order="2" place="2" resultid="2464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7538" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3841" />
                    <RANKING order="2" place="2" resultid="3196" />
                    <RANKING order="3" place="3" resultid="3491" />
                    <RANKING order="4" place="4" resultid="5112" />
                    <RANKING order="5" place="5" resultid="4880" />
                    <RANKING order="6" place="-1" resultid="2412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7539" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2452" />
                    <RANKING order="2" place="2" resultid="1830" />
                    <RANKING order="3" place="3" resultid="4040" />
                    <RANKING order="4" place="4" resultid="1668" />
                    <RANKING order="5" place="5" resultid="4058" />
                    <RANKING order="6" place="6" resultid="7625" />
                    <RANKING order="7" place="7" resultid="4045" />
                    <RANKING order="8" place="-1" resultid="2270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7540" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4086" />
                    <RANKING order="2" place="2" resultid="4052" />
                    <RANKING order="3" place="3" resultid="3967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7541" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2405" />
                    <RANKING order="2" place="2" resultid="3008" />
                    <RANKING order="3" place="3" resultid="4022" />
                    <RANKING order="4" place="4" resultid="3974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7542" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1950" />
                    <RANKING order="2" place="2" resultid="1907" />
                    <RANKING order="3" place="3" resultid="3986" />
                    <RANKING order="4" place="4" resultid="2430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7543" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4936" />
                    <RANKING order="2" place="2" resultid="3811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7544" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7545" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7546" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7150" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7151" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7152" daytime="11:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7153" daytime="11:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7154" daytime="11:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1543" daytime="11:15" gender="M" number="31" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7547" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2325" />
                    <RANKING order="2" place="2" resultid="5089" />
                    <RANKING order="3" place="3" resultid="4332" />
                    <RANKING order="4" place="4" resultid="3140" />
                    <RANKING order="5" place="5" resultid="3924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7548" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4876" />
                    <RANKING order="2" place="2" resultid="3081" />
                    <RANKING order="3" place="3" resultid="4304" />
                    <RANKING order="4" place="4" resultid="5476" />
                    <RANKING order="5" place="5" resultid="4319" />
                    <RANKING order="6" place="6" resultid="3585" />
                    <RANKING order="7" place="7" resultid="4312" />
                    <RANKING order="8" place="8" resultid="2757" />
                    <RANKING order="9" place="9" resultid="4263" />
                    <RANKING order="10" place="-1" resultid="4253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7549" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4211" />
                    <RANKING order="2" place="2" resultid="1696" />
                    <RANKING order="3" place="3" resultid="3456" />
                    <RANKING order="4" place="4" resultid="3867" />
                    <RANKING order="5" place="-1" resultid="5502" />
                    <RANKING order="6" place="-1" resultid="3542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7550" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3589" />
                    <RANKING order="2" place="2" resultid="3504" />
                    <RANKING order="3" place="3" resultid="3476" />
                    <RANKING order="4" place="4" resultid="1708" />
                    <RANKING order="5" place="5" resultid="4862" />
                    <RANKING order="6" place="6" resultid="1717" />
                    <RANKING order="7" place="7" resultid="3511" />
                    <RANKING order="8" place="8" resultid="5076" />
                    <RANKING order="9" place="9" resultid="2393" />
                    <RANKING order="10" place="-1" resultid="4922" />
                    <RANKING order="11" place="-1" resultid="3484" />
                    <RANKING order="12" place="-1" resultid="2568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7551" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3427" />
                    <RANKING order="2" place="2" resultid="4939" />
                    <RANKING order="3" place="3" resultid="2511" />
                    <RANKING order="4" place="4" resultid="1922" />
                    <RANKING order="5" place="5" resultid="2371" />
                    <RANKING order="6" place="6" resultid="3215" />
                    <RANKING order="7" place="7" resultid="1693" />
                    <RANKING order="8" place="8" resultid="2521" />
                    <RANKING order="9" place="9" resultid="4983" />
                    <RANKING order="10" place="10" resultid="3741" />
                    <RANKING order="11" place="11" resultid="3748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7552" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4105" />
                    <RANKING order="2" place="2" resultid="3000" />
                    <RANKING order="3" place="3" resultid="1720" />
                    <RANKING order="4" place="4" resultid="3707" />
                    <RANKING order="5" place="5" resultid="3055" />
                    <RANKING order="6" place="-1" resultid="2311" />
                    <RANKING order="7" place="-1" resultid="3030" />
                    <RANKING order="8" place="-1" resultid="1688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7553" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4240" />
                    <RANKING order="2" place="2" resultid="2882" />
                    <RANKING order="3" place="3" resultid="2835" />
                    <RANKING order="4" place="4" resultid="5162" />
                    <RANKING order="5" place="5" resultid="1755" />
                    <RANKING order="6" place="6" resultid="2349" />
                    <RANKING order="7" place="7" resultid="2620" />
                    <RANKING order="8" place="-1" resultid="2749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7554" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2590" />
                    <RANKING order="2" place="2" resultid="1807" />
                    <RANKING order="3" place="3" resultid="5680" />
                    <RANKING order="4" place="4" resultid="3949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7555" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5123" />
                    <RANKING order="2" place="2" resultid="1816" />
                    <RANKING order="3" place="3" resultid="4010" />
                    <RANKING order="4" place="4" resultid="3579" />
                    <RANKING order="5" place="5" resultid="7598" />
                    <RANKING order="6" place="6" resultid="3895" />
                    <RANKING order="7" place="7" resultid="3714" />
                    <RANKING order="8" place="8" resultid="1627" />
                    <RANKING order="9" place="9" resultid="1854" />
                    <RANKING order="10" place="10" resultid="2993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7556" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3906" />
                    <RANKING order="2" place="2" resultid="2789" />
                    <RANKING order="3" place="3" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7557" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1957" />
                    <RANKING order="2" place="2" resultid="1901" />
                    <RANKING order="3" place="3" resultid="4003" />
                    <RANKING order="4" place="4" resultid="3942" />
                    <RANKING order="5" place="5" resultid="4298" />
                    <RANKING order="6" place="-1" resultid="3693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7558" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4033" />
                    <RANKING order="2" place="2" resultid="2986" />
                    <RANKING order="3" place="3" resultid="2684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7559" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7560" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7155" daytime="11:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7156" daytime="11:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7157" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7158" daytime="11:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7159" daytime="11:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7160" daytime="11:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7161" daytime="11:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7162" daytime="11:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7163" daytime="11:35" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1558" daytime="11:35" gender="F" number="32" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7561" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1763" />
                    <RANKING order="2" place="2" resultid="3860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7562" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                    <RANKING order="2" place="2" resultid="5145" />
                    <RANKING order="3" place="3" resultid="1651" />
                    <RANKING order="4" place="-1" resultid="3817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7563" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2572" />
                    <RANKING order="2" place="2" resultid="4228" />
                    <RANKING order="3" place="3" resultid="4857" />
                    <RANKING order="4" place="4" resultid="2283" />
                    <RANKING order="5" place="5" resultid="3095" />
                    <RANKING order="6" place="6" resultid="4133" />
                    <RANKING order="7" place="7" resultid="3208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7564" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1615" />
                    <RANKING order="2" place="2" resultid="2630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7565" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5138" />
                    <RANKING order="2" place="2" resultid="3200" />
                    <RANKING order="3" place="3" resultid="2400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7566" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2870" />
                    <RANKING order="2" place="2" resultid="2446" />
                    <RANKING order="3" place="3" resultid="2919" />
                    <RANKING order="4" place="4" resultid="4822" />
                    <RANKING order="5" place="5" resultid="2807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7567" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4117" />
                    <RANKING order="2" place="2" resultid="4029" />
                    <RANKING order="3" place="3" resultid="2584" />
                    <RANKING order="4" place="4" resultid="1647" />
                    <RANKING order="5" place="5" resultid="2276" />
                    <RANKING order="6" place="6" resultid="2607" />
                    <RANKING order="7" place="7" resultid="7626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7568" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1837" />
                    <RANKING order="2" place="2" resultid="5117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7569" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4081" />
                    <RANKING order="2" place="2" resultid="2778" />
                    <RANKING order="3" place="3" resultid="3220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7570" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7571" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/" />
                <AGEGROUP agegroupid="7572" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/" />
                <AGEGROUP agegroupid="7573" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7574" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7164" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7165" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7166" daytime="12:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7167" daytime="12:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1573" daytime="12:10" gender="M" number="33" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7575" agemax="24" agemin="20" name="KATEGORIA  WIEKOWA: &quot;0&quot; /20-24/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2326" />
                    <RANKING order="2" place="2" resultid="3766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7576" agemax="29" agemin="25" name="KATEGORIA  WIEKOWA: &quot;A&quot; /25-29/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4204" />
                    <RANKING order="2" place="2" resultid="1972" />
                    <RANKING order="3" place="3" resultid="3153" />
                    <RANKING order="4" place="4" resultid="4234" />
                    <RANKING order="5" place="5" resultid="3823" />
                    <RANKING order="6" place="6" resultid="4187" />
                    <RANKING order="7" place="7" resultid="5095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7577" agemax="34" agemin="30" name="KATEGORIA  WIEKOWA: &quot;B&quot;/30-34/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3881" />
                    <RANKING order="2" place="2" resultid="3075" />
                    <RANKING order="3" place="3" resultid="5657" />
                    <RANKING order="4" place="4" resultid="3160" />
                    <RANKING order="5" place="5" resultid="3888" />
                    <RANKING order="6" place="-1" resultid="2819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7578" agemax="39" agemin="35" name="KATEGORIA  WIEKOWA: &quot;C&quot;/35-39/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3449" />
                    <RANKING order="2" place="2" resultid="3769" />
                    <RANKING order="3" place="3" resultid="2866" />
                    <RANKING order="4" place="4" resultid="2389" />
                    <RANKING order="5" place="5" resultid="3477" />
                    <RANKING order="6" place="6" resultid="2533" />
                    <RANKING order="7" place="7" resultid="3754" />
                    <RANKING order="8" place="8" resultid="4977" />
                    <RANKING order="9" place="9" resultid="3614" />
                    <RANKING order="10" place="10" resultid="3166" />
                    <RANKING order="11" place="11" resultid="2049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7579" agemax="44" agemin="40" name="KATEGORIA  WIEKOWA: &quot;D&quot;/40-44/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3428" />
                    <RANKING order="2" place="2" resultid="4965" />
                    <RANKING order="3" place="3" resultid="3436" />
                    <RANKING order="4" place="4" resultid="3731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7580" agemax="49" agemin="45" name="KATEGORIA  WIEKOWA: &quot;E&quot;45-49/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3646" />
                    <RANKING order="2" place="2" resultid="2979" />
                    <RANKING order="3" place="3" resultid="4288" />
                    <RANKING order="4" place="4" resultid="4222" />
                    <RANKING order="5" place="5" resultid="2343" />
                    <RANKING order="6" place="6" resultid="3018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7581" agemax="54" agemin="50" name="KATEGORIA  WIEKOWA: &quot;F&quot;/50-54/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2812" />
                    <RANKING order="2" place="2" resultid="2858" />
                    <RANKING order="3" place="3" resultid="1789" />
                    <RANKING order="4" place="4" resultid="2350" />
                    <RANKING order="5" place="5" resultid="3779" />
                    <RANKING order="6" place="6" resultid="3147" />
                    <RANKING order="7" place="-1" resultid="4831" />
                    <RANKING order="8" place="-1" resultid="4893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7582" agemax="59" agemin="55" name="KATEGORIA  WIEKOWA: &quot;G&quot;/55-59/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4123" />
                    <RANKING order="2" place="2" resultid="4172" />
                    <RANKING order="3" place="3" resultid="2614" />
                    <RANKING order="4" place="4" resultid="3799" />
                    <RANKING order="5" place="5" resultid="4915" />
                    <RANKING order="6" place="-1" resultid="2064" />
                    <RANKING order="7" place="-1" resultid="1897" />
                    <RANKING order="8" place="-1" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7583" agemax="64" agemin="60" name="KATEGORIA  WIEKOWA: &quot;H&quot;/60-64/">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7584" agemax="69" agemin="65" name="KATEGORIA  WIEKOWA: &quot;I&quot;/65-69/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2378" />
                    <RANKING order="2" place="2" resultid="3062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7585" agemax="74" agemin="70" name="KATEGORIA  WIEKOWA: &quot;J&quot;/70-74/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2850" />
                    <RANKING order="2" place="2" resultid="3686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7586" agemax="79" agemin="75" name="KATEGORIA  WIEKOWA: &quot;K&quot;/75-79/">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1885" />
                    <RANKING order="2" place="2" resultid="3654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7587" agemax="84" agemin="80" name="KATEGORIA  WIEKOWA: &quot;L&quot;/80-84/" />
                <AGEGROUP agegroupid="7588" agemax="89" agemin="85" name="KATEGORIA  WIEKOWA: &quot;M&quot;/85-89/" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7168" daytime="12:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7169" daytime="12:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7170" daytime="12:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7171" daytime="12:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7172" daytime="12:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7173" daytime="12:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7174" daytime="12:55" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="AZALM" name="AZS Almamer" nation="POL">
          <CONTACT name="sołtyk judyta" />
          <ATHLETES>
            <ATHLETE birthdate="1974-11-19" firstname="judyta" gender="F" lastname="sołtyk" nation="POL" athleteid="1613">
              <RESULTS>
                <RESULT eventid="1361" points="412" swimtime="00:02:31.81" resultid="1614" heatid="7081" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:52.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="419" swimtime="00:05:19.54" resultid="1615" heatid="7167" lane="2" entrytime="00:05:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                    <SPLIT distance="200" swimtime="00:02:35.36" />
                    <SPLIT distance="250" swimtime="00:03:16.52" />
                    <SPLIT distance="300" swimtime="00:03:58.24" />
                    <SPLIT distance="350" swimtime="00:04:39.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01511" name="MTP Delfin Cieszyn" nation="POL" region="SLA">
          <CONTACT name="Widzik" />
          <ATHLETES>
            <ATHLETE birthdate="1986-05-25" firstname="Łukasz" gender="M" lastname="Widzik" nation="POL" athleteid="1617">
              <RESULTS>
                <RESULT eventid="1134" points="421" swimtime="00:00:32.07" resultid="1618" heatid="6996" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1316" points="415" swimtime="00:01:09.58" resultid="1619" heatid="7072" lane="0" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="1620" heatid="7089" lane="6" entrytime="00:02:13.00" />
                <RESULT eventid="1498" points="427" swimtime="00:02:28.55" resultid="1621" heatid="7146" lane="7" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Ryszard" gender="M" lastname="Jabłecki" nation="POL" athleteid="1623">
              <RESULTS>
                <RESULT eventid="1104" points="150" swimtime="00:03:59.52" resultid="1624" heatid="6975" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.61" />
                    <SPLIT distance="100" swimtime="00:01:57.59" />
                    <SPLIT distance="150" swimtime="00:03:00.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="149" swimtime="00:00:50.23" resultid="1625" heatid="7053" lane="4" entrytime="00:00:47.00" />
                <RESULT eventid="1468" points="124" swimtime="00:00:41.85" resultid="1626" heatid="7122" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1543" points="145" swimtime="00:01:51.31" resultid="1627" heatid="7156" lane="6" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEZR" name="niezrzeszony" nation="POL" region="LU">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1984-08-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" license="1" athleteid="1629">
              <RESULTS>
                <RESULT eventid="1194" points="322" swimtime="00:01:08.44" resultid="1630" heatid="7016" lane="3" entrytime="00:01:07.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="1631" heatid="7129" lane="3" entrytime="00:00:29.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-03-18" firstname="Tomasz" gender="M" lastname="Najderek" nation="POL" athleteid="1776">
              <RESULTS>
                <RESULT eventid="1194" points="482" swimtime="00:00:59.82" resultid="1777" heatid="7020" lane="8" entrytime="00:01:01.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="342" swimtime="00:02:25.79" resultid="1778" heatid="7089" lane="8" entrytime="00:02:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="150" swimtime="00:01:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="502" swimtime="00:00:26.30" resultid="1779" heatid="7135" lane="6" entrytime="00:00:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="SINICKI" nation="POL" athleteid="1780">
              <RESULTS>
                <RESULT eventid="1256" points="306" swimtime="00:00:33.27" resultid="1781" heatid="7041" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1376" points="283" swimtime="00:02:35.26" resultid="1782" heatid="7086" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="331" swimtime="00:00:30.22" resultid="1783" heatid="7130" lane="0" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="1848">
              <RESULTS>
                <RESULT eventid="1134" points="72" swimtime="00:00:57.74" resultid="1849" heatid="6988" lane="8" entrytime="00:00:58.00" />
                <RESULT eventid="1224" points="46" swimtime="00:05:10.21" resultid="1850" heatid="7025" lane="2" entrytime="00:05:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.22" />
                    <SPLIT distance="100" swimtime="00:02:30.68" />
                    <SPLIT distance="150" swimtime="00:03:54.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="63" swimtime="00:00:56.20" resultid="1851" heatid="7036" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1376" points="61" swimtime="00:04:18.06" resultid="1852" heatid="7082" lane="5" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.61" />
                    <SPLIT distance="100" swimtime="00:02:02.61" />
                    <SPLIT distance="150" swimtime="00:03:12.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="51" swimtime="00:02:13.52" resultid="1853" heatid="7106" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="90" swimtime="00:02:10.36" resultid="1854" heatid="7156" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-30" firstname="Krzysztof" gender="M" lastname="Krzak" nation="POL" athleteid="2529">
              <RESULTS>
                <RESULT eventid="1104" points="329" swimtime="00:03:04.28" resultid="2530" heatid="6978" lane="8" entrytime="00:03:11.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:29.30" />
                    <SPLIT distance="150" swimtime="00:02:17.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2531" heatid="7057" lane="6" entrytime="00:00:37.71" entrycourse="LCM" />
                <RESULT eventid="1573" points="325" swimtime="00:05:20.03" resultid="2533" heatid="7172" lane="8" entrytime="00:05:16.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="150" swimtime="00:01:53.54" />
                    <SPLIT distance="200" swimtime="00:02:34.21" />
                    <SPLIT distance="250" swimtime="00:03:15.59" />
                    <SPLIT distance="300" swimtime="00:03:57.34" />
                    <SPLIT distance="350" swimtime="00:04:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="340" swimtime="00:02:43.28" resultid="5491" heatid="7100" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Andrzej" gender="M" lastname="Michałkowski" nation="POL" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1104" points="149" swimtime="00:03:59.79" resultid="3574" heatid="6975" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.42" />
                    <SPLIT distance="100" swimtime="00:01:51.73" />
                    <SPLIT distance="150" swimtime="00:02:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="126" swimtime="00:01:33.42" resultid="3575" heatid="7011" lane="7" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="231" swimtime="00:00:43.43" resultid="3576" heatid="7055" lane="7" entrytime="00:00:43.50" />
                <RESULT eventid="1376" points="95" swimtime="00:03:42.94" resultid="3577" heatid="7083" lane="0" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:43.81" />
                    <SPLIT distance="150" swimtime="00:02:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="161" swimtime="00:00:38.43" resultid="3578" heatid="7123" lane="3" entrytime="00:00:37.50" />
                <RESULT eventid="1543" points="180" swimtime="00:01:43.65" resultid="3579" heatid="7157" lane="7" entrytime="00:01:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="3580">
              <RESULTS>
                <RESULT eventid="1104" points="355" swimtime="00:02:59.69" resultid="3581" heatid="6979" lane="7" entrytime="00:03:03.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:02:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="374" swimtime="00:01:05.10" resultid="3582" heatid="7017" lane="6" entrytime="00:01:05.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="445" swimtime="00:00:34.93" resultid="3583" heatid="7060" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1468" points="368" swimtime="00:00:29.16" resultid="3584" heatid="7130" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1543" points="378" swimtime="00:01:20.95" resultid="3585" heatid="7162" lane="8" entrytime="00:01:18.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Arkadiusz" gender="M" lastname="Bilski" nation="POL" athleteid="3586">
              <RESULTS>
                <RESULT eventid="1104" points="424" swimtime="00:02:49.33" resultid="3587" heatid="6980" lane="1" entrytime="00:02:45.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="448" swimtime="00:00:34.83" resultid="3588" heatid="7061" lane="9" entrytime="00:00:32.60" />
                <RESULT eventid="1543" points="447" swimtime="00:01:16.59" resultid="3589" heatid="7163" lane="8" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Ewa" gender="F" lastname="Balcewicz" nation="POL" athleteid="3590">
              <RESULTS>
                <RESULT eventid="1271" points="289" swimtime="00:00:45.06" resultid="3591" heatid="7051" lane="6" entrytime="00:00:36.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="3592">
              <RESULTS>
                <RESULT eventid="1134" points="237" swimtime="00:00:38.81" resultid="3593" heatid="6992" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1194" points="268" swimtime="00:01:12.67" resultid="3594" heatid="7014" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="170" swimtime="00:00:40.42" resultid="3595" heatid="7038" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1316" points="185" swimtime="00:01:31.13" resultid="3596" heatid="7069" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="263" swimtime="00:00:32.63" resultid="3597" heatid="7127" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1498" points="156" swimtime="00:03:27.85" resultid="3598" heatid="7143" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                    <SPLIT distance="100" swimtime="00:01:43.69" />
                    <SPLIT distance="150" swimtime="00:02:37.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="3599">
              <RESULTS>
                <RESULT eventid="1271" points="85" swimtime="00:01:07.70" resultid="3600" heatid="7048" lane="7" entrytime="00:01:13.85" />
                <RESULT eventid="1453" points="115" swimtime="00:00:48.72" resultid="3601" heatid="7115" lane="0" entrytime="00:00:53.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Karolina" gender="F" lastname="Szczuka" nation="POL" athleteid="3602">
              <RESULTS>
                <RESULT eventid="1422" points="336" swimtime="00:01:20.57" resultid="3603" heatid="7105" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="456" swimtime="00:00:30.83" resultid="3604" heatid="7120" lane="9" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Michał" gender="M" lastname="Mandes" nation="POL" athleteid="3607">
              <RESULTS>
                <RESULT eventid="1194" points="389" swimtime="00:01:04.24" resultid="3608" heatid="7017" lane="0" entrytime="00:01:06.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="393" swimtime="00:00:30.60" resultid="3609" heatid="7041" lane="6" entrytime="00:00:32.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Marek" gender="M" lastname="Żuber" nation="POL" athleteid="3610">
              <RESULTS>
                <RESULT eventid="1194" points="390" swimtime="00:01:04.16" resultid="3611" heatid="7020" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="372" swimtime="00:00:31.16" resultid="3612" heatid="7043" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1468" points="395" swimtime="00:00:28.48" resultid="3613" heatid="7132" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1573" points="296" swimtime="00:05:30.11" resultid="3614" heatid="7171" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:18.61" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                    <SPLIT distance="200" swimtime="00:02:44.41" />
                    <SPLIT distance="250" swimtime="00:03:27.34" />
                    <SPLIT distance="300" swimtime="00:04:11.02" />
                    <SPLIT distance="350" swimtime="00:04:53.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Robert" gender="M" lastname="Budek" nation="POL" athleteid="3615">
              <RESULTS>
                <RESULT eventid="1316" points="100" swimtime="00:01:51.57" resultid="3616" heatid="7066" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="109" swimtime="00:03:58.17" resultid="3617" heatid="7095" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                    <SPLIT distance="100" swimtime="00:01:59.08" />
                    <SPLIT distance="150" swimtime="00:03:09.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Rafał" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3618">
              <RESULTS>
                <RESULT eventid="1256" points="98" swimtime="00:00:48.57" resultid="3619" heatid="7037" lane="2" />
                <RESULT eventid="1468" points="203" swimtime="00:00:35.55" resultid="3620" heatid="7121" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Magda" gender="F" lastname="Konieczkowska" nation="POL" athleteid="3621">
              <RESULTS>
                <RESULT eventid="1528" points="237" swimtime="00:01:44.00" resultid="3622" heatid="7150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Paweł" gender="M" lastname="Sadowski" nation="POL" athleteid="3623">
              <RESULTS>
                <RESULT eventid="1468" points="79" swimtime="00:00:48.70" resultid="3624" heatid="7121" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Andrzej" gender="M" lastname="Gadaś" nation="POL" athleteid="3625">
              <RESULTS>
                <RESULT eventid="1286" points="367" swimtime="00:00:37.24" resultid="3626" heatid="7052" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="Cieplucha" nation="POL" athleteid="3673">
              <RESULTS>
                <RESULT eventid="1119" points="423" swimtime="00:00:36.02" resultid="3674" heatid="6986" lane="8" entrytime="00:00:37.13" />
                <RESULT comment="Rekord Polski Masters w kat. E /30-34/" eventid="1301" points="408" swimtime="00:01:18.30" resultid="3675" heatid="7065" lane="7" entrytime="00:01:19.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-14" firstname="Przemysław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="3676">
              <RESULTS>
                <RESULT eventid="1194" points="540" swimtime="00:00:57.60" resultid="3677" heatid="7020" lane="1" entrytime="00:01:00.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="505" swimtime="00:00:28.15" resultid="3678" heatid="7044" lane="5" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Piotr" gender="M" lastname="Capała" nation="POL" athleteid="3767">
              <RESULTS>
                <RESULT eventid="1376" points="437" swimtime="00:02:14.33" resultid="3768" heatid="7090" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="150" swimtime="00:01:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="424" swimtime="00:04:52.79" resultid="3769" heatid="7174" lane="3" entrytime="00:04:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                    <SPLIT distance="200" swimtime="00:02:20.43" />
                    <SPLIT distance="250" swimtime="00:02:57.85" />
                    <SPLIT distance="300" swimtime="00:03:36.27" />
                    <SPLIT distance="350" swimtime="00:04:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Piotr" gender="M" lastname="Słotwiński" nation="POL" athleteid="3770">
              <RESULTS>
                <RESULT eventid="1194" points="626" swimtime="00:00:54.83" resultid="3771" heatid="7022" lane="3" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Piotr" gender="M" lastname="Szczuka" nation="POL" athleteid="3772">
              <RESULTS>
                <RESULT eventid="1438" points="492" swimtime="00:01:03.10" resultid="3773" heatid="7112" lane="1" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="492" swimtime="00:00:26.48" resultid="3774" heatid="7136" lane="7" entrytime="00:00:25.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Leszek" gender="M" lastname="Rąpała" nation="POL" athleteid="3775">
              <RESULTS>
                <RESULT eventid="1256" points="145" swimtime="00:00:42.68" resultid="3776" heatid="7036" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1406" points="115" swimtime="00:03:53.77" resultid="3777" heatid="7096" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:59.81" />
                    <SPLIT distance="150" swimtime="00:03:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="226" swimtime="00:00:34.28" resultid="3778" heatid="7126" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1573" points="160" swimtime="00:06:45.08" resultid="3779" heatid="7169" lane="1" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:33.87" />
                    <SPLIT distance="150" swimtime="00:02:25.39" />
                    <SPLIT distance="200" swimtime="00:03:20.38" />
                    <SPLIT distance="250" swimtime="00:04:13.52" />
                    <SPLIT distance="300" swimtime="00:05:07.82" />
                    <SPLIT distance="350" swimtime="00:06:00.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Tomasz" gender="M" lastname="Rozmysłowski" nation="POL" athleteid="3780">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="3782" heatid="7020" lane="0" entrytime="00:01:01.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3784" heatid="7102" lane="9" entrytime="00:02:40.00" />
                <RESULT eventid="1468" points="439" swimtime="00:00:27.51" resultid="3785" heatid="7133" lane="0" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Paweł" gender="M" lastname="Rumin" nation="POL" athleteid="3787">
              <RESULTS>
                <RESULT eventid="1468" points="446" swimtime="00:00:27.35" resultid="3788" heatid="7133" lane="7" entrytime="00:00:27.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Michał" gender="M" lastname="Skrzyński" nation="POL" athleteid="3789">
              <RESULTS>
                <RESULT eventid="1194" points="510" swimtime="00:00:58.70" resultid="3790" heatid="7021" lane="1" entrytime="00:00:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="479" swimtime="00:00:28.65" resultid="3791" heatid="7044" lane="2" entrytime="00:00:28.90" />
                <RESULT eventid="1406" points="479" swimtime="00:02:25.61" resultid="3792" heatid="7102" lane="5" entrytime="00:02:31.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="3793" heatid="7134" lane="7" entrytime="00:00:26.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Wojciech" gender="M" lastname="Szcześniak" nation="POL" athleteid="3794">
              <RESULTS>
                <RESULT eventid="1194" points="199" swimtime="00:01:20.25" resultid="3795" heatid="7012" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3796" heatid="7039" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1376" points="156" swimtime="00:03:09.27" resultid="3797" heatid="7084" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="160" swimtime="00:06:45.24" resultid="3799" heatid="7169" lane="2" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:33.67" />
                    <SPLIT distance="150" swimtime="00:02:25.47" />
                    <SPLIT distance="200" swimtime="00:03:19.53" />
                    <SPLIT distance="250" swimtime="00:04:14.19" />
                    <SPLIT distance="300" swimtime="00:05:08.41" />
                    <SPLIT distance="350" swimtime="00:06:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="222" swimtime="00:00:34.50" resultid="7619" heatid="7128" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Igor" gender="M" lastname="Zbrzeski" nation="POL" athleteid="3832">
              <RESULTS>
                <RESULT eventid="1468" points="377" swimtime="00:00:28.92" resultid="3833" heatid="7132" lane="1" entrytime="00:00:27.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Arkadiusz" gender="M" lastname="Doliński" nation="POL" athleteid="4124">
              <RESULTS>
                <RESULT eventid="1134" points="308" swimtime="00:00:35.57" resultid="4125" heatid="6993" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1316" points="303" swimtime="00:01:17.32" resultid="4126" heatid="7069" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Emilia" gender="F" lastname="Sopolińska" nation="POL" athleteid="4127">
              <RESULTS>
                <RESULT eventid="1058" points="188" swimtime="00:04:04.45" resultid="4128" heatid="6971" lane="3" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.81" />
                    <SPLIT distance="100" swimtime="00:01:57.14" />
                    <SPLIT distance="150" swimtime="00:03:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="235" swimtime="00:01:24.28" resultid="4129" heatid="7006" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="210" swimtime="00:03:10.06" resultid="4130" heatid="7079" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                    <SPLIT distance="150" swimtime="00:02:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="184" swimtime="00:03:41.62" resultid="4131" heatid="7092" lane="6" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.52" />
                    <SPLIT distance="100" swimtime="00:01:51.90" />
                    <SPLIT distance="150" swimtime="00:02:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="248" swimtime="00:00:37.74" resultid="4132" heatid="7117" lane="0" entrytime="00:00:37.60" />
                <RESULT eventid="1558" points="203" swimtime="00:06:46.35" resultid="4133" heatid="7165" lane="4" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:34.26" />
                    <SPLIT distance="150" swimtime="00:02:26.07" />
                    <SPLIT distance="200" swimtime="00:03:17.50" />
                    <SPLIT distance="250" swimtime="00:04:10.16" />
                    <SPLIT distance="300" swimtime="00:05:03.44" />
                    <SPLIT distance="350" swimtime="00:05:56.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Krzysztof" gender="M" lastname="Nowogrodzki" nation="POL" athleteid="4134">
              <RESULTS>
                <RESULT eventid="1194" points="443" swimtime="00:01:01.52" resultid="4135" heatid="7019" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="409" swimtime="00:00:28.16" resultid="4136" heatid="7130" lane="7" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" athleteid="4137">
              <RESULTS>
                <RESULT eventid="1240" points="417" swimtime="00:00:33.55" resultid="4138" heatid="7034" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1301" points="360" swimtime="00:01:21.65" resultid="4139" heatid="7065" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-16" firstname="Monika" gender="F" lastname="Winogrodzka" nation="POL" athleteid="4161">
              <RESULTS>
                <RESULT eventid="1119" points="373" swimtime="00:00:37.59" resultid="4162" heatid="6986" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1179" points="319" swimtime="00:01:16.19" resultid="4163" heatid="7008" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="309" swimtime="00:00:44.07" resultid="4164" heatid="7051" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1453" points="385" swimtime="00:00:32.61" resultid="4165" heatid="7120" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Małgorzata" gender="F" lastname="Michałkiewicz" nation="POL" athleteid="5155">
              <RESULTS>
                <RESULT eventid="1058" points="356" swimtime="00:03:17.58" resultid="5156" heatid="6973" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:34.29" />
                    <SPLIT distance="150" swimtime="00:02:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="335" swimtime="00:00:42.89" resultid="5157" heatid="7051" lane="0" entrytime="00:00:39.50" />
                <RESULT eventid="1528" points="345" swimtime="00:01:31.88" resultid="5159" heatid="7154" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Witold" gender="M" lastname="Szczechla" nation="POL" athleteid="5160">
              <RESULTS>
                <RESULT eventid="1256" points="213" swimtime="00:00:37.52" resultid="5161" heatid="7038" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1543" points="223" swimtime="00:01:36.57" resultid="5162" heatid="7157" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Michał " gender="M" lastname="Rożalski" nation="POL" athleteid="5473">
              <RESULTS>
                <RESULT eventid="1286" points="500" swimtime="00:00:33.59" resultid="5474" heatid="7060" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="1468" points="432" swimtime="00:00:27.65" resultid="5475" heatid="7133" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1543" points="439" swimtime="00:01:17.07" resultid="5476" heatid="7161" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="F" lastname="Kotusińska " nation="POL" athleteid="5481">
              <RESULTS>
                <RESULT eventid="1179" points="255" swimtime="00:01:22.09" resultid="5482" heatid="7006" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="224" swimtime="00:00:41.26" resultid="5483" heatid="7033" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Ewa" gender="F" lastname="Galica" nation="POL" athleteid="5484">
              <RESULTS>
                <RESULT eventid="1240" points="410" swimtime="00:00:33.73" resultid="5485" heatid="7034" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1453" points="414" swimtime="00:00:31.82" resultid="5487" heatid="7120" lane="2" entrytime="00:00:29.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="5674">
              <RESULTS>
                <RESULT eventid="1134" points="248" swimtime="00:00:38.24" resultid="5675" heatid="6993" lane="2" entrytime="00:00:36.70" />
                <RESULT eventid="1224" points="201" swimtime="00:03:10.11" resultid="5676" heatid="7027" lane="4" entrytime="00:03:06.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:26.33" />
                    <SPLIT distance="150" swimtime="00:02:18.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="335" swimtime="00:00:38.39" resultid="5677" heatid="7057" lane="4" entrytime="00:00:37.45" />
                <RESULT eventid="1406" points="231" swimtime="00:03:05.55" resultid="5678" heatid="7099" lane="9" entrytime="00:02:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:22.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="205" swimtime="00:01:24.38" resultid="5679" heatid="7109" lane="8" entrytime="00:01:21.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="285" swimtime="00:01:28.99" resultid="5680" heatid="7159" lane="6" entrytime="00:01:26.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Emil" gender="M" lastname="Paciorkowski" nation="POL" athleteid="6418">
              <RESULTS>
                <RESULT eventid="1194" points="231" swimtime="00:01:16.39" resultid="6419" heatid="7013" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="6420" heatid="7085" lane="0" entrytime="00:02:50.00" />
                <RESULT comment="O-4 - Przedwczwsny start" eventid="1468" status="DSQ" swimtime="00:00:33.50" resultid="6421" heatid="7127" lane="0" entrytime="00:00:31.70" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="6422" heatid="7025" lane="5" entrytime="00:04:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Volodymyr" gender="M" lastname="Timofeyev" nation="POL" athleteid="7596">
              <RESULTS>
                <RESULT eventid="1286" points="183" swimtime="00:00:46.97" resultid="7597" heatid="7052" lane="1" />
                <RESULT eventid="1543" points="163" swimtime="00:01:47.14" resultid="7598" heatid="7155" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Krzysztof" gender="M" lastname="Klepko" nation="POL" athleteid="7611" />
            <ATHLETE birthdate="1987-01-01" firstname="sEWERYN" gender="M" lastname="aFANSJEW" nation="POL" athleteid="7624" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1346" points="497" swimtime="00:01:47.08" resultid="3800" heatid="7076" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="100" swimtime="00:00:55.01" />
                    <SPLIT distance="150" swimtime="00:01:19.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3772" number="1" />
                    <RELAYPOSITION athleteid="7611" number="2" />
                    <RELAYPOSITION athleteid="3770" number="3" />
                    <RELAYPOSITION athleteid="3767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1513" points="114" swimtime="00:03:12.38" resultid="3627" heatid="7147" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.70" />
                    <SPLIT distance="100" swimtime="00:01:56.95" />
                    <SPLIT distance="150" swimtime="00:02:39.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3615" number="1" />
                    <RELAYPOSITION athleteid="3618" number="2" />
                    <RELAYPOSITION athleteid="3621" number="3" />
                    <RELAYPOSITION athleteid="7624" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAELB" name="Victory Masters Elbląg" nation="POL" region="WAR">
          <CONTACT name="LATECKI GRZEGORZ" phone="606147184" />
          <ATHLETES>
            <ATHLETE birthdate="1965-03-12" firstname="GRZEGORZ" gender="M" lastname="LATECKI" nation="POL" athleteid="1633">
              <RESULTS>
                <RESULT eventid="1134" points="386" swimtime="00:00:32.99" resultid="1634" heatid="6995" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1194" points="409" swimtime="00:01:03.18" resultid="1635" heatid="7019" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="419" swimtime="00:00:29.97" resultid="1636" heatid="7043" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1406" points="375" swimtime="00:02:38.06" resultid="1637" heatid="7102" lane="8" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:15.53" />
                    <SPLIT distance="150" swimtime="00:02:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="379" swimtime="00:01:08.79" resultid="1638" heatid="7111" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="377" swimtime="00:00:28.93" resultid="1639" heatid="7133" lane="9" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="ANDRZEJ" gender="M" lastname="PASIECZNY" nation="POL" athleteid="1640">
              <RESULTS>
                <RESULT eventid="1224" points="429" swimtime="00:02:27.79" resultid="1641" heatid="7029" lane="7" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:09.42" />
                    <SPLIT distance="150" swimtime="00:01:47.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="BEATA" gender="F" lastname="KARAŚ" nation="POL" athleteid="1642">
              <RESULTS>
                <RESULT eventid="1209" points="117" swimtime="00:04:08.65" resultid="1643" heatid="7023" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                    <SPLIT distance="100" swimtime="00:01:55.30" />
                    <SPLIT distance="150" swimtime="00:03:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="162" swimtime="00:03:27.00" resultid="1644" heatid="7078" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:40.91" />
                    <SPLIT distance="150" swimtime="00:02:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="128" swimtime="00:04:09.97" resultid="1645" heatid="7092" lane="0" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.53" />
                    <SPLIT distance="100" swimtime="00:02:01.58" />
                    <SPLIT distance="150" swimtime="00:03:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="116" swimtime="00:01:54.85" resultid="1646" heatid="7104" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="150" swimtime="00:07:29.72" resultid="1647" heatid="7165" lane="0" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.19" />
                    <SPLIT distance="100" swimtime="00:01:48.84" />
                    <SPLIT distance="150" swimtime="00:02:45.31" />
                    <SPLIT distance="200" swimtime="00:03:42.96" />
                    <SPLIT distance="250" swimtime="00:04:40.11" />
                    <SPLIT distance="300" swimtime="00:05:37.96" />
                    <SPLIT distance="350" swimtime="00:06:34.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-30" firstname="KAROLINA" gender="F" lastname="KARAŚ" nation="POL" athleteid="1648">
              <RESULTS>
                <RESULT eventid="1179" points="130" swimtime="00:01:42.70" resultid="1649" heatid="7003" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="129" swimtime="00:03:43.27" resultid="1650" heatid="7078" lane="1" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                    <SPLIT distance="100" swimtime="00:01:46.95" />
                    <SPLIT distance="150" swimtime="00:02:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="128" swimtime="00:07:54.47" resultid="1651" heatid="7164" lane="4" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:50.52" />
                    <SPLIT distance="150" swimtime="00:02:50.91" />
                    <SPLIT distance="200" swimtime="00:03:52.92" />
                    <SPLIT distance="250" swimtime="00:04:54.95" />
                    <SPLIT distance="300" swimtime="00:05:55.69" />
                    <SPLIT distance="350" swimtime="00:06:56.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-18" firstname="TOMASZ" gender="M" lastname="GLEB" nation="POL" athleteid="1652">
              <RESULTS>
                <RESULT eventid="1104" points="267" swimtime="00:03:17.61" resultid="1653" heatid="6976" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:34.03" />
                    <SPLIT distance="150" swimtime="00:02:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="355" swimtime="00:01:06.20" resultid="1654" heatid="7017" lane="8" entrytime="00:01:06.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="1655" heatid="7087" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="1656" heatid="7131" lane="0" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EULVI" name="Euro-Lviv" nation="UKR">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+38 032 2430304" name="Masters Swimming Club &quot;Euro-Lviv&quot;" phone="+38 067 6734796" street="Karpincya Str. 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1978-05-16" firstname="Iryna" gender="F" lastname="Bura" nation="UKR" athleteid="1658">
              <RESULTS>
                <RESULT eventid="1453" points="350" swimtime="00:00:33.66" resultid="1659" heatid="7119" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1179" points="312" swimtime="00:01:16.73" resultid="5582" heatid="7007" lane="7" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-06" firstname="Lyudmyla" gender="F" lastname="Khiresh" nation="UKR" athleteid="1660">
              <RESULTS>
                <RESULT eventid="1119" points="291" swimtime="00:00:40.81" resultid="1661" heatid="6984" lane="5" entrytime="00:00:41.75" />
                <RESULT eventid="1453" points="262" swimtime="00:00:37.05" resultid="1662" heatid="7117" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-11-30" firstname="Tetiana" gender="F" lastname="Kozakova" nation="UKR" athleteid="1663">
              <RESULTS>
                <RESULT eventid="1119" points="138" swimtime="00:00:52.26" resultid="1664" heatid="6983" lane="8" entrytime="00:00:51.20" />
                <RESULT eventid="1453" points="118" swimtime="00:00:48.36" resultid="1665" heatid="7115" lane="1" entrytime="00:00:50.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-11" firstname="Lyudmyla" gender="F" lastname="Maksymiv" nation="UKR" athleteid="1666">
              <RESULTS>
                <RESULT eventid="1271" points="209" swimtime="00:00:50.17" resultid="1667" heatid="7049" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1528" points="223" swimtime="00:01:46.28" resultid="1668" heatid="7152" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="1669">
              <RESULTS>
                <RESULT eventid="1119" points="336" swimtime="00:00:38.92" resultid="1670" heatid="6986" lane="9" entrytime="00:00:38.20" />
                <RESULT eventid="1240" points="343" swimtime="00:00:35.81" resultid="1671" heatid="7033" lane="4" entrytime="00:00:35.20" />
                <RESULT eventid="1301" points="275" swimtime="00:01:29.32" resultid="1672" heatid="7065" lane="0" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="284" swimtime="00:01:37.98" resultid="1673" heatid="7153" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-06" firstname="Mariia" gender="F" lastname="Vasylko" nation="UKR" athleteid="1674">
              <RESULTS>
                <RESULT eventid="1240" points="174" swimtime="00:00:44.90" resultid="1675" heatid="7031" lane="5" entrytime="00:00:45.50" />
                <RESULT eventid="1361" points="137" swimtime="00:03:38.76" resultid="1676" heatid="7078" lane="6" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.75" />
                    <SPLIT distance="100" swimtime="00:01:43.77" />
                    <SPLIT distance="150" swimtime="00:02:43.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="127" swimtime="00:07:55.15" resultid="7626" heatid="7166" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                    <SPLIT distance="100" swimtime="00:01:49.24" />
                    <SPLIT distance="150" swimtime="00:02:50.76" />
                    <SPLIT distance="200" swimtime="00:03:53.02" />
                    <SPLIT distance="250" swimtime="00:04:54.09" />
                    <SPLIT distance="300" swimtime="00:05:57.13" />
                    <SPLIT distance="350" swimtime="00:06:59.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-06" firstname="Yuriy" gender="M" lastname="Chyrkov" nation="UKR" athleteid="1678">
              <RESULTS>
                <RESULT eventid="1256" points="256" swimtime="00:00:35.31" resultid="1679" heatid="7040" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1406" points="190" swimtime="00:03:18.20" resultid="1680" heatid="7097" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                    <SPLIT distance="150" swimtime="00:02:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="287" swimtime="00:00:31.70" resultid="1681" heatid="7126" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-10-14" firstname="Stepan" gender="M" lastname="Delyatynskyy" nation="UKR" athleteid="1682">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="1683" heatid="7018" lane="0" entrytime="00:01:04.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1684" heatid="7057" lane="5" entrytime="00:00:37.50" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="1685" heatid="7131" lane="8" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-08" firstname="Andriy" gender="M" lastname="Hertsyk" nation="UKR" athleteid="1686">
              <RESULTS>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1687" heatid="7056" lane="2" entrytime="00:00:39.85" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="1688" heatid="7159" lane="9" entrytime="00:01:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="1689">
              <RESULTS>
                <RESULT eventid="1134" points="258" swimtime="00:00:37.76" resultid="1690" heatid="6995" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1286" points="311" swimtime="00:00:39.34" resultid="1691" heatid="7058" lane="4" entrytime="00:00:36.42" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="1692" heatid="7100" lane="5" entrytime="00:02:45.39" />
                <RESULT eventid="1543" points="294" swimtime="00:01:28.03" resultid="1693" heatid="7159" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-08" firstname="Dmytro" gender="M" lastname="Konovalov" nation="UKR" athleteid="1694">
              <RESULTS>
                <RESULT eventid="1286" points="583" swimtime="00:00:31.91" resultid="1695" heatid="7061" lane="5" entrytime="00:00:30.75" />
                <RESULT eventid="1543" points="500" swimtime="00:01:13.78" resultid="1696" heatid="7163" lane="3" entrytime="00:01:08.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-31" firstname="Roman" gender="M" lastname="Koretskyy" nation="UKR" athleteid="1697">
              <RESULTS>
                <RESULT eventid="1134" points="133" swimtime="00:00:47.07" resultid="1698" heatid="6990" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1468" points="156" swimtime="00:00:38.79" resultid="1699" heatid="7124" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-05-31" firstname="Zenoviy" gender="M" lastname="Kushnir" nation="UKR" athleteid="1700">
              <RESULTS>
                <RESULT eventid="1134" points="78" swimtime="00:00:56.26" resultid="1701" heatid="6989" lane="8" entrytime="00:00:51.00" />
                <RESULT eventid="1286" points="95" swimtime="00:00:58.32" resultid="1702" heatid="7053" lane="1" entrytime="00:00:55.50" />
                <RESULT eventid="1468" points="85" swimtime="00:00:47.52" resultid="5583" heatid="7122" lane="0" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-27" firstname="Iurii" gender="M" lastname="Martyniuk" nation="UKR" athleteid="1703">
              <RESULTS>
                <RESULT eventid="1194" points="279" swimtime="00:01:11.75" resultid="1704" heatid="7016" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="298" swimtime="00:00:31.30" resultid="1705" heatid="7130" lane="2" entrytime="00:00:28.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="1706">
              <RESULTS>
                <RESULT eventid="1286" points="443" swimtime="00:00:34.97" resultid="1707" heatid="7060" lane="3" entrytime="00:00:33.50" />
                <RESULT eventid="1543" points="371" swimtime="00:01:21.46" resultid="1708" heatid="7162" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-13" firstname="Bogdan" gender="M" lastname="Osidach" nation="UKR" athleteid="1709">
              <RESULTS>
                <RESULT eventid="1468" points="298" swimtime="00:00:31.28" resultid="1710" heatid="7129" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1194" points="305" swimtime="00:01:09.66" resultid="5584" heatid="7016" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-08" firstname="Igor" gender="M" lastname="Rudnyk" nation="UKR" athleteid="1711">
              <RESULTS>
                <RESULT eventid="1376" points="234" swimtime="00:02:45.39" resultid="1712" heatid="7085" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                    <SPLIT distance="150" swimtime="00:01:59.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="1713" heatid="7098" lane="6" entrytime="00:03:00.00" />
                <RESULT eventid="1468" points="282" swimtime="00:00:31.87" resultid="1714" heatid="7126" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1134" points="231" swimtime="00:00:39.17" resultid="5585" heatid="6992" lane="2" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-23" firstname="Oleksandr" gender="M" lastname="Shavrov" nation="UKR" athleteid="1715">
              <RESULTS>
                <RESULT eventid="1286" points="386" swimtime="00:00:36.60" resultid="1716" heatid="7059" lane="3" entrytime="00:00:35.16" />
                <RESULT eventid="1543" points="305" swimtime="00:01:26.99" resultid="1717" heatid="7161" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-13" firstname="Igor" gender="M" lastname="Yaskevych" nation="UKR" athleteid="1718">
              <RESULTS>
                <RESULT eventid="1286" points="299" swimtime="00:00:39.86" resultid="1719" heatid="7057" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1543" points="253" swimtime="00:01:32.52" resultid="1720" heatid="7159" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-11-07" firstname="Bohdan" gender="M" lastname="Yatsura" nation="UKR" athleteid="1721">
              <RESULTS>
                <RESULT eventid="1194" points="213" swimtime="00:01:18.54" resultid="1722" heatid="7012" lane="4" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="161" swimtime="00:00:41.23" resultid="1723" heatid="7037" lane="7" entrytime="00:00:40.45" />
                <RESULT eventid="1468" points="225" swimtime="00:00:34.37" resultid="1724" heatid="7125" lane="3" entrytime="00:00:33.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-02" firstname="Serhiy" gender="M" lastname="Zhykh" nation="UKR" athleteid="1725">
              <RESULTS>
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="1726" heatid="6995" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="1727" heatid="7131" lane="9" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-10" firstname="Serhiy" gender="M" lastname="Fedorov" nation="UKR" athleteid="1728">
              <RESULTS>
                <RESULT eventid="1256" points="286" swimtime="00:00:34.02" resultid="1729" heatid="7041" lane="0" entrytime="00:00:33.30" />
                <RESULT eventid="1468" points="328" swimtime="00:00:30.29" resultid="1730" heatid="7129" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-05" firstname="Oleksiy" gender="M" lastname="Shalayev" nation="UKR" athleteid="5586">
              <RESULTS>
                <RESULT eventid="1406" points="339" swimtime="00:02:43.34" resultid="5587" heatid="7101" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="377" swimtime="00:01:08.93" resultid="5588" heatid="7110" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1164" points="379" swimtime="00:02:09.10" resultid="7221" heatid="7001" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:38.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1689" number="1" />
                    <RELAYPOSITION athleteid="1694" number="2" />
                    <RELAYPOSITION athleteid="1706" number="3" />
                    <RELAYPOSITION athleteid="1728" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1346" points="362" swimtime="00:01:59.00" resultid="7607" heatid="7074" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:01.22" />
                    <SPLIT distance="150" swimtime="00:01:27.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1694" number="1" />
                    <RELAYPOSITION athleteid="1711" number="2" />
                    <RELAYPOSITION athleteid="1678" number="3" />
                    <RELAYPOSITION athleteid="1728" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1149" points="240" swimtime="00:02:50.76" resultid="7220" heatid="6998" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                    <SPLIT distance="100" swimtime="00:01:39.88" />
                    <SPLIT distance="150" swimtime="00:02:15.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1663" number="1" />
                    <RELAYPOSITION athleteid="1666" number="2" />
                    <RELAYPOSITION athleteid="1674" number="3" />
                    <RELAYPOSITION athleteid="1669" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1331" points="265" swimtime="00:02:30.48" resultid="7610" heatid="7608" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:01:52.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1658" number="1" />
                    <RELAYPOSITION athleteid="1674" number="2" />
                    <RELAYPOSITION athleteid="1669" number="3" />
                    <RELAYPOSITION athleteid="1660" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1513" points="233" swimtime="00:02:31.63" resultid="7622" heatid="7147" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1663" number="1" />
                    <RELAYPOSITION athleteid="1694" number="2" />
                    <RELAYPOSITION athleteid="1669" number="3" />
                    <RELAYPOSITION athleteid="1703" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1513" points="226" swimtime="00:02:33.31" resultid="7623" heatid="7147" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:01:25.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1660" number="1" />
                    <RELAYPOSITION athleteid="1689" number="2" />
                    <RELAYPOSITION athleteid="1674" number="3" />
                    <RELAYPOSITION athleteid="1678" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01910" name="KS Delfin Gdynia" nation="POL" region="POM">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" license="S01910200065" athleteid="1732">
              <RESULTS>
                <RESULT eventid="1224" points="293" swimtime="00:02:47.84" resultid="1733" heatid="7028" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:04.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="425" swimtime="00:00:29.81" resultid="1734" heatid="7044" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1438" points="387" swimtime="00:01:08.34" resultid="1735" heatid="7111" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="413" swimtime="00:00:28.07" resultid="1736" heatid="7131" lane="4" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-24" firstname="Aleksandra" gender="F" lastname="Sypniewska" nation="POL" license="S01910100045" athleteid="1737">
              <RESULTS>
                <RESULT eventid="1361" points="337" swimtime="00:02:42.33" resultid="1738" heatid="7081" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:58.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="354" swimtime="00:05:38.03" resultid="1739" heatid="7167" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="150" swimtime="00:02:01.41" />
                    <SPLIT distance="200" swimtime="00:02:44.29" />
                    <SPLIT distance="250" swimtime="00:03:27.73" />
                    <SPLIT distance="300" swimtime="00:04:11.64" />
                    <SPLIT distance="350" swimtime="00:04:55.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEGLI" name="KS Delfin Gliwice" nation="POL" region="SLA">
          <CONTACT city="Gliwice" email="ksdelfin@op.pl" name="Cupiał" phone="605065587" state="ŚLASK" street="Stwosza" street2="8/3" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="1741">
              <RESULTS>
                <RESULT eventid="1104" points="58" swimtime="00:05:28.75" resultid="1742" heatid="6974" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.98" />
                    <SPLIT distance="100" swimtime="00:02:35.69" />
                    <SPLIT distance="150" swimtime="00:04:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="43" swimtime="00:01:08.51" resultid="1743" heatid="6987" lane="7" />
                <RESULT eventid="1286" points="87" swimtime="00:01:00.02" resultid="1744" heatid="7052" lane="4" entrytime="00:00:58.86" entrycourse="LCM" />
                <RESULT eventid="1316" points="24" swimtime="00:02:58.63" resultid="1745" heatid="7066" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="47" swimtime="00:00:57.63" resultid="1746" heatid="7121" lane="6" entrytime="00:00:56.48" entrycourse="LCM" />
                <RESULT eventid="1543" points="67" swimtime="00:02:24.01" resultid="1747" heatid="7155" lane="3" entrytime="00:02:17.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01202" name="KP Delfin Inowrocław" nation="POL" region="KUJ">
          <CONTACT city="Inowrocław" email="jarek.molenda@gmail.com" name="Molenda Jarosław" phone="660 899 358" state="KUJ" street="Wierzbińskiego 11" zip="88-100" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-28" firstname="Krzysztof" gender="M" lastname="Derkowski" nation="POL" license="M01202200043" athleteid="1749">
              <RESULTS>
                <RESULT eventid="1134" points="137" swimtime="00:00:46.53" resultid="1750" heatid="6990" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1194" points="206" swimtime="00:01:19.37" resultid="1751" heatid="7012" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="222" swimtime="00:00:36.99" resultid="1752" heatid="7038" lane="4" entrytime="00:00:37.20" />
                <RESULT eventid="1286" points="241" swimtime="00:00:42.85" resultid="1753" heatid="7056" lane="9" entrytime="00:00:41.65" />
                <RESULT eventid="1468" points="236" swimtime="00:00:33.80" resultid="1754" heatid="7126" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1543" points="206" swimtime="00:01:39.11" resultid="1755" heatid="7157" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZKRA" name="AZS UJ Kraków" nation="POL" region="MAL">
          <CONTACT city="Kraków" name="Michał Syryca" state="MAL" street="ul. Piastowska 26d" zip="30-067" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-01" firstname="Karolina" gender="F" lastname="Zadrożna" nation="POL" athleteid="1757">
              <RESULTS>
                <RESULT eventid="1119" points="327" swimtime="00:00:39.27" resultid="1758" heatid="6986" lane="2" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1179" points="415" swimtime="00:01:09.76" resultid="1759" heatid="7008" lane="7" entrytime="00:01:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="292" swimtime="00:01:27.57" resultid="1760" heatid="7065" lane="3" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="381" swimtime="00:02:35.73" resultid="1761" heatid="7081" lane="6" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                    <SPLIT distance="150" swimtime="00:01:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="393" swimtime="00:00:32.37" resultid="1762" heatid="7119" lane="4" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1558" points="411" swimtime="00:05:21.62" resultid="1763" heatid="7167" lane="5" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:56.87" />
                    <SPLIT distance="200" swimtime="00:02:37.93" />
                    <SPLIT distance="250" swimtime="00:03:19.50" />
                    <SPLIT distance="300" swimtime="00:04:00.69" />
                    <SPLIT distance="350" swimtime="00:04:42.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KUAZ" name="KU AZS Uniwersytet Rolniczy im H  Kołłątaja" nation="POL" region="MAZ">
          <CONTACT city="Kraków" email="manuela.nawrocka@gmail.com" name="Nawrocka Manuela" phone="606704926" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="1765">
              <RESULTS>
                <RESULT eventid="1058" points="352" swimtime="00:03:18.37" resultid="1766" heatid="6973" lane="3" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:33.34" />
                    <SPLIT distance="150" swimtime="00:02:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="398" swimtime="00:00:36.77" resultid="1767" heatid="6986" lane="6" entrytime="00:00:35.70" />
                <RESULT eventid="1271" points="365" swimtime="00:00:41.68" resultid="1768" heatid="7051" lane="9" entrytime="00:00:39.50" />
                <RESULT eventid="1391" points="393" swimtime="00:02:52.13" resultid="1769" heatid="7094" lane="6" entrytime="00:02:44.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="433" swimtime="00:00:31.36" resultid="1770" heatid="7120" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="1771" heatid="7154" lane="2" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-16" firstname="Michalina" gender="F" lastname="Bąk" nation="POL" athleteid="1772">
              <RESULTS>
                <RESULT eventid="1179" points="548" swimtime="00:01:03.60" resultid="1773" heatid="7008" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="489" swimtime="00:00:31.80" resultid="1774" heatid="7034" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1361" points="433" swimtime="00:02:29.27" resultid="1775" heatid="7081" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:49.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ODOPO" name="Odrzańskie Ratownictwo Specjalistyczne Opole" nation="POL" region="OPO">
          <CONTACT name="Waldemar Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="1785">
              <RESULTS>
                <RESULT eventid="1194" points="277" swimtime="00:01:11.91" resultid="1786" heatid="7015" lane="8" entrytime="00:01:10.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="271" swimtime="00:02:37.57" resultid="1787" heatid="7086" lane="6" entrytime="00:02:35.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:56.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="139" swimtime="00:03:35.72" resultid="1788" heatid="7142" lane="7" entrytime="00:03:40.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:48.01" />
                    <SPLIT distance="150" swimtime="00:02:43.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="271" swimtime="00:05:39.81" resultid="1789" heatid="7171" lane="9" entrytime="00:05:35.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:05.07" />
                    <SPLIT distance="200" swimtime="00:02:48.51" />
                    <SPLIT distance="250" swimtime="00:03:31.81" />
                    <SPLIT distance="300" swimtime="00:04:15.26" />
                    <SPLIT distance="350" swimtime="00:04:59.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="1790">
              <RESULTS>
                <RESULT eventid="1179" points="272" swimtime="00:01:20.29" resultid="1791" heatid="7005" lane="5" entrytime="00:01:22.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="277" swimtime="00:01:29.12" resultid="1792" heatid="7064" lane="7" entrytime="00:01:30.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="276" swimtime="00:03:13.65" resultid="1793" heatid="7093" lane="6" entrytime="00:03:15.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:02:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="265" swimtime="00:03:14.15" resultid="1794" heatid="7139" lane="0" entrytime="00:03:09.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:02:25.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01805" name="Z-Ł Wopr Ozorków" nation="POL" region="LOD">
          <CONTACT city="OZORKÓW" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁODZK" street="LOTNICZA 1" zip="95-035" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-09" firstname="WŁODZIMIERZ" gender="M" lastname="PRZYTULSKI" nation="POL" license="M0180520005" athleteid="1796">
              <RESULTS>
                <RESULT eventid="1134" points="289" swimtime="00:00:36.34" resultid="1797" heatid="6993" lane="3" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="319" swimtime="00:00:32.81" resultid="1798" heatid="7041" lane="4" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="1799" heatid="7087" lane="0" entrytime="00:02:32.00" entrycourse="LCM" />
                <RESULT eventid="1438" points="239" swimtime="00:01:20.19" resultid="1800" heatid="7109" lane="2" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-20" firstname="BOGDAN" gender="M" lastname="WĄSIK" nation="POL" license="M0180520002" athleteid="1801">
              <RESULTS>
                <RESULT eventid="1104" points="280" swimtime="00:03:14.56" resultid="1802" heatid="6977" lane="2" entrytime="00:03:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:34.85" />
                    <SPLIT distance="150" swimtime="00:02:24.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="1803" heatid="7026" lane="1" entrytime="00:03:40.00" entrycourse="LCM" />
                <RESULT eventid="1286" points="288" swimtime="00:00:40.38" resultid="1804" heatid="7056" lane="7" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="1805" heatid="7097" lane="7" entrytime="00:03:20.00" entrycourse="LCM" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="1806" heatid="7107" lane="5" entrytime="00:01:36.00" entrycourse="LCM" />
                <RESULT eventid="1543" points="287" swimtime="00:01:28.74" resultid="1807" heatid="7158" lane="4" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="ZBIGNIEW" gender="M" lastname="MACIEJCZYK" nation="POL" license="M01805" athleteid="1808">
              <RESULTS>
                <RESULT eventid="1194" points="250" swimtime="00:01:14.39" resultid="1809" heatid="7014" lane="8" entrytime="00:01:14.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="207" swimtime="00:00:37.91" resultid="1810" heatid="7039" lane="8" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1438" points="116" swimtime="00:01:42.00" resultid="1811" heatid="7107" lane="3" entrytime="00:01:38.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="239" swimtime="00:00:33.65" resultid="1812" heatid="7125" lane="4" entrytime="00:00:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="ROMAN" gender="M" lastname="WICZEL" nation="POL" license="M0180520003" athleteid="1813">
              <RESULTS>
                <RESULT eventid="1104" points="229" swimtime="00:03:27.94" resultid="1814" heatid="6977" lane="7" entrytime="00:03:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                    <SPLIT distance="100" swimtime="00:01:36.72" />
                    <SPLIT distance="150" swimtime="00:02:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="254" swimtime="00:00:42.07" resultid="1815" heatid="7056" lane="3" entrytime="00:00:39.01" entrycourse="LCM" />
                <RESULT eventid="1543" points="249" swimtime="00:01:33.07" resultid="1816" heatid="7159" lane="0" entrytime="00:01:29.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="URSZULA" gender="F" lastname="MRÓZ" nation="POL" license="M0180510002" athleteid="1817">
              <RESULTS>
                <RESULT eventid="1119" points="319" swimtime="00:00:39.57" resultid="1818" heatid="6985" lane="1" entrytime="00:00:40.01" entrycourse="LCM" />
                <RESULT eventid="1179" points="279" swimtime="00:01:19.66" resultid="1819" heatid="7004" lane="8" entrytime="00:01:30.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="298" swimtime="00:00:37.52" resultid="1820" heatid="7033" lane="7" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1361" points="233" swimtime="00:03:03.45" resultid="1821" heatid="7080" lane="0" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="243" swimtime="00:01:29.76" resultid="1822" heatid="7105" lane="2" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="311" swimtime="00:00:34.99" resultid="1823" heatid="7118" lane="0" entrytime="00:00:35.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="EWA" gender="F" lastname="STĘPIEŃ" nation="POL" license="M0180510003" athleteid="1824">
              <RESULTS>
                <RESULT eventid="1119" points="312" swimtime="00:00:39.87" resultid="1825" heatid="6984" lane="6" entrytime="00:00:42.08" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters w kat. F /50-54/" eventid="1179" points="339" swimtime="00:01:14.62" resultid="1826" heatid="7006" lane="6" entrytime="00:01:16.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. F /50-54/" eventid="1271" points="388" swimtime="00:00:40.84" resultid="1827" heatid="7050" lane="7" entrytime="00:00:41.30" entrycourse="LCM" />
                <RESULT eventid="1361" points="276" swimtime="00:02:53.45" resultid="1828" heatid="7080" lane="8" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="150" swimtime="00:02:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat F /50-54/" eventid="1453" points="382" swimtime="00:00:32.69" resultid="1829" heatid="7119" lane="9" entrytime="00:00:33.15" entrycourse="LCM" />
                <RESULT eventid="1528" points="334" swimtime="00:01:32.81" resultid="1830" heatid="7153" lane="6" entrytime="00:01:31.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-13" firstname="MIROSŁAWA" gender="F" lastname="RAJTAR" nation="POL" license="M0180510004" athleteid="1831">
              <RESULTS>
                <RESULT eventid="1119" points="217" swimtime="00:00:44.97" resultid="1832" heatid="6984" lane="7" entrytime="00:00:44.60" entrycourse="LCM" />
                <RESULT eventid="1179" points="252" swimtime="00:01:22.38" resultid="1833" heatid="7005" lane="6" entrytime="00:01:22.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="185" swimtime="00:00:43.99" resultid="1834" heatid="7032" lane="9" entrytime="00:00:43.80" entrycourse="LCM" />
                <RESULT eventid="1391" points="203" swimtime="00:03:34.46" resultid="1835" heatid="7094" lane="4" entrytime="00:02:31.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:38.70" />
                    <SPLIT distance="150" swimtime="00:02:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="244" swimtime="00:00:37.97" resultid="1836" heatid="7117" lane="9" entrytime="00:00:37.60" entrycourse="LCM" />
                <RESULT eventid="1558" points="198" swimtime="00:06:49.98" resultid="1837" heatid="7165" lane="6" entrytime="00:06:47.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                    <SPLIT distance="200" swimtime="00:03:16.96" />
                    <SPLIT distance="250" swimtime="00:04:10.63" />
                    <SPLIT distance="300" swimtime="00:05:04.57" />
                    <SPLIT distance="350" swimtime="00:05:57.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="TADEUSZ" gender="M" lastname="OBIEDZIŃSKI" nation="POL" license="M01805" athleteid="2745">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="2746" heatid="6976" lane="8" entrytime="00:03:40.00" entrycourse="LCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="2747" heatid="7037" lane="5" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2748" heatid="7056" lane="1" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2749" heatid="7158" lane="0" entrytime="00:01:35.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="229" swimtime="00:02:32.65" resultid="1838" heatid="7000" lane="9" entrytime="00:02:27.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1796" number="1" />
                    <RELAYPOSITION athleteid="1813" number="2" />
                    <RELAYPOSITION athleteid="1801" number="3" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1346" points="232" swimtime="00:02:17.92" resultid="1839" heatid="7074" lane="4" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:45.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1796" number="1" />
                    <RELAYPOSITION athleteid="1801" number="2" />
                    <RELAYPOSITION athleteid="1813" number="3" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1513" points="248" swimtime="00:02:28.52" resultid="1840" heatid="7149" lane="8" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1817" number="1" />
                    <RELAYPOSITION athleteid="1796" number="2" />
                    <RELAYPOSITION athleteid="1824" number="3" />
                    <RELAYPOSITION athleteid="1808" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KUPOZ" name="Ku Azs Uam Poznań" nation="POL" region="WIE">
          <CONTACT city="Poznań" name="Ziemniarski Bartosz" phone="691679381" state="WLKP" street="ul. Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-22" firstname="Bartosz" gender="M" lastname="Ziemniarski" nation="POL" license="S03315100001" athleteid="1856">
              <RESULTS>
                <RESULT eventid="1194" points="653" swimtime="00:00:54.06" resultid="1857" heatid="7022" lane="6" entrytime="00:00:54.81" entrycourse="LCM" />
                <RESULT eventid="1256" points="589" swimtime="00:00:26.75" resultid="1858" heatid="7045" lane="6" entrytime="00:00:27.39" entrycourse="LCM" />
                <RESULT eventid="1468" points="638" swimtime="00:00:24.28" resultid="1859" heatid="7136" lane="6" entrytime="00:00:24.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" name="MKS &quot;Neptun&quot; Stargard Szcz." nation="POL" region="SZ">
          <CONTACT city="Stargard Szcz" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Międzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1982-10-19" firstname="Tomasz" gender="M" lastname="SULEJA" nation="POL" athleteid="1861">
              <RESULTS>
                <RESULT eventid="1194" points="552" swimtime="00:00:57.16" resultid="1862" heatid="7021" lane="5" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="404" swimtime="00:02:17.88" resultid="1863" heatid="7088" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="517" swimtime="00:00:26.05" resultid="1864" heatid="7135" lane="5" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04514" name="Uks 307" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" name="Ilczyszyn" state="MAZ" street="barcelońska 8" zip="02-762" />
          <ATHLETES>
            <ATHLETE birthdate="1983-07-13" firstname="Krzysztof" gender="M" lastname="Ilczyszyn" nation="POL" athleteid="1866">
              <RESULTS>
                <RESULT eventid="1194" points="394" swimtime="00:01:03.94" resultid="1867" heatid="7019" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="408" swimtime="00:00:30.23" resultid="1868" heatid="7042" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="1376" points="275" swimtime="00:02:36.78" resultid="1869" heatid="7087" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:01:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="274" swimtime="00:01:16.62" resultid="1870" heatid="7109" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="352" swimtime="00:00:29.60" resultid="1871" heatid="7132" lane="5" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="Ziółkowski" nation="POL" athleteid="1872">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="1873" heatid="7019" lane="9" entrytime="00:01:03.00" />
                <RESULT eventid="1256" points="360" swimtime="00:00:31.52" resultid="1874" heatid="7043" lane="9" entrytime="00:00:30.50" />
                <RESULT eventid="1376" points="329" swimtime="00:02:27.67" resultid="1875" heatid="7087" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="241" swimtime="00:01:19.99" resultid="1876" heatid="7109" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="387" swimtime="00:00:28.67" resultid="1877" heatid="7132" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2959" heatid="7100" lane="8" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEINO" name="Delfin Inowrocław" nation="POL" region="KUJ">
          <CONTACT city="INOWROCŁAW" name="LEWANDOWSKI ZYGMUNT" state="KUJ-P" street="WIERZBIŃSKIEGO" zip="88-100" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="ZYGMUNT" gender="M" lastname="LEWANDOWSKI" nation="POL" athleteid="1879">
              <RESULTS>
                <RESULT eventid="1134" points="115" swimtime="00:00:49.33" resultid="1880" heatid="6988" lane="6" entrytime="00:00:55.00" entrycourse="LCM" />
                <RESULT eventid="1194" points="132" swimtime="00:01:31.90" resultid="1881" heatid="7011" lane="8" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="90" swimtime="00:00:49.96" resultid="1882" heatid="7036" lane="6" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1376" points="121" swimtime="00:03:25.86" resultid="1883" heatid="7083" lane="1" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:39.99" />
                    <SPLIT distance="150" swimtime="00:02:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="65" swimtime="00:02:03.68" resultid="1884" heatid="7106" lane="5" entrytime="00:01:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="134" swimtime="00:07:09.95" resultid="1885" heatid="7168" lane="3" entrytime="00:07:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:42.73" />
                    <SPLIT distance="150" swimtime="00:02:38.22" />
                    <SPLIT distance="200" swimtime="00:03:33.85" />
                    <SPLIT distance="250" swimtime="00:04:29.31" />
                    <SPLIT distance="300" swimtime="00:05:25.61" />
                    <SPLIT distance="350" swimtime="00:06:19.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WEZAB" name="Weteran Zabrze" nation="POL" region="SLA">
          <CONTACT email="WETERANZABRZE@OP.PL" name="BOSOWSKI WŁODZIMIERZ" />
          <ATHLETES>
            <ATHLETE birthdate="1947-01-01" firstname="Henryk" gender="M" lastname="Wachnik" nation="POL" athleteid="1887">
              <RESULTS>
                <RESULT eventid="1134" points="22" swimtime="00:01:25.60" resultid="1888" heatid="6987" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1194" points="31" swimtime="00:02:28.10" resultid="1889" heatid="7010" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="1890" heatid="7066" lane="3" entrytime="00:02:35.00" />
                <RESULT eventid="1468" points="27" swimtime="00:01:09.47" resultid="1891" heatid="7121" lane="3" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="1892">
              <RESULTS>
                <RESULT eventid="1134" points="180" swimtime="00:00:42.55" resultid="1893" heatid="6992" lane="9" entrytime="00:00:40.50" />
                <RESULT eventid="1194" points="294" swimtime="00:01:10.52" resultid="1894" heatid="7016" lane="8" entrytime="00:01:09.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="220" swimtime="00:02:48.95" resultid="1895" heatid="7086" lane="0" entrytime="00:02:41.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:19.67" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="309" swimtime="00:00:30.90" resultid="1896" heatid="7128" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="1897" heatid="7170" lane="8" entrytime="00:05:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" athleteid="1898">
              <RESULTS>
                <RESULT eventid="1104" points="214" swimtime="00:03:32.64" resultid="1899" heatid="6976" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:45.66" />
                    <SPLIT distance="150" swimtime="00:02:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="193" swimtime="00:00:46.09" resultid="1900" heatid="7055" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1543" points="192" swimtime="00:01:41.45" resultid="1901" heatid="7158" lane="7" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" athleteid="1902">
              <RESULTS>
                <RESULT eventid="1058" points="206" swimtime="00:03:57.15" resultid="1903" heatid="6971" lane="5" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.27" />
                    <SPLIT distance="100" swimtime="00:01:56.27" />
                    <SPLIT distance="150" swimtime="00:02:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1209" points="126" swimtime="00:04:02.53" resultid="1904" heatid="7024" lane="1" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.52" />
                    <SPLIT distance="100" swimtime="00:01:59.66" />
                    <SPLIT distance="150" swimtime="00:03:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="176" swimtime="00:00:53.13" resultid="1905" heatid="7049" lane="9" entrytime="00:00:54.00" />
                <RESULT eventid="1422" points="131" swimtime="00:01:50.29" resultid="1906" heatid="7104" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="185" swimtime="00:01:52.95" resultid="1907" heatid="7152" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" athleteid="1908">
              <RESULTS>
                <RESULT eventid="1194" points="220" swimtime="00:01:17.64" resultid="1909" heatid="7015" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="238" swimtime="00:00:36.19" resultid="1910" heatid="7039" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1468" points="257" swimtime="00:00:32.86" resultid="1911" heatid="7128" lane="9" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" athleteid="1912">
              <RESULTS>
                <RESULT eventid="1058" points="400" swimtime="00:03:10.09" resultid="1913" heatid="6973" lane="6" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:20.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="403" swimtime="00:01:10.48" resultid="1914" heatid="7008" lane="9" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="378" swimtime="00:00:41.20" resultid="1915" heatid="7051" lane="1" entrytime="00:00:39.00" />
                <RESULT comment="Rekord Polski Masters w kat. D /40-45/" eventid="1391" points="402" swimtime="00:02:50.92" resultid="1916" heatid="7094" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="382" swimtime="00:01:28.76" resultid="1917" heatid="7154" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Tadeusz" gender="M" lastname="Stuchlik" nation="POL" athleteid="1918">
              <RESULTS>
                <RESULT eventid="1134" points="448" swimtime="00:00:31.41" resultid="1919" heatid="6996" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1256" points="456" swimtime="00:00:29.12" resultid="1920" heatid="7044" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1286" points="418" swimtime="00:00:35.66" resultid="1921" heatid="7060" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1543" points="363" swimtime="00:01:22.09" resultid="1922" heatid="7161" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Marek" gender="M" lastname="Roter" nation="POL" athleteid="1923">
              <RESULTS>
                <RESULT eventid="1134" points="433" swimtime="00:00:31.76" resultid="1924" heatid="6996" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1316" points="415" swimtime="00:01:09.61" resultid="1925" heatid="7072" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="381" swimtime="00:02:20.64" resultid="1926" heatid="7088" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="402" swimtime="00:02:31.64" resultid="1927" heatid="7146" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" athleteid="1928">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat.H /60-64/" eventid="1119" points="316" swimtime="00:00:39.70" resultid="1929" heatid="6985" lane="3" entrytime="00:00:40.00" />
                <RESULT comment="Rekord Polski Masters w kat. H /60-64/" eventid="1209" points="169" swimtime="00:03:40.22" resultid="1930" heatid="7024" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                    <SPLIT distance="100" swimtime="00:01:46.04" />
                    <SPLIT distance="150" swimtime="00:02:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. H /60-64/" eventid="1240" points="248" swimtime="00:00:39.85" resultid="1931" heatid="7032" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1301" points="281" swimtime="00:01:28.70" resultid="1932" heatid="7064" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat H /60-64/" eventid="1483" points="259" swimtime="00:03:15.60" resultid="1933" heatid="7138" lane="6" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:35.11" />
                    <SPLIT distance="150" swimtime="00:02:26.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Stanisław" gender="M" lastname="Kiszczak" nation="POL" athleteid="1934">
              <RESULTS>
                <RESULT eventid="1134" points="147" swimtime="00:00:45.48" resultid="1935" heatid="6990" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1468" points="237" swimtime="00:00:33.76" resultid="1936" heatid="7125" lane="2" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" athleteid="1937">
              <RESULTS>
                <RESULT eventid="1179" points="173" swimtime="00:01:33.28" resultid="1938" heatid="7003" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="134" swimtime="00:03:40.41" resultid="1939" heatid="7078" lane="8" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.19" />
                    <SPLIT distance="100" swimtime="00:01:43.32" />
                    <SPLIT distance="150" swimtime="00:02:42.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="184" swimtime="00:00:41.69" resultid="1940" heatid="7116" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" athleteid="1941">
              <RESULTS>
                <RESULT eventid="1134" points="173" swimtime="00:00:43.14" resultid="1942" heatid="6990" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1316" points="132" swimtime="00:01:41.95" resultid="1943" heatid="7068" lane="9" entrytime="00:01:37.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="111" swimtime="00:03:52.25" resultid="1944" heatid="7142" lane="1" entrytime="00:03:42.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                    <SPLIT distance="100" swimtime="00:01:50.08" />
                    <SPLIT distance="150" swimtime="00:02:52.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Maria" gender="F" lastname="Buczkowska" nation="POL" athleteid="1945">
              <RESULTS>
                <RESULT eventid="1058" points="192" swimtime="00:04:02.71" resultid="1946" heatid="6971" lane="7" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.49" />
                    <SPLIT distance="100" swimtime="00:01:58.76" />
                    <SPLIT distance="150" swimtime="00:03:01.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="1948" heatid="7031" lane="8" entrytime="00:00:51.00" />
                <RESULT eventid="1271" points="236" swimtime="00:00:48.21" resultid="1949" heatid="7049" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1528" points="206" swimtime="00:01:49.03" resultid="1950" heatid="7152" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="Władysław" gender="M" lastname="Buczkowski" nation="POL" athleteid="1951">
              <RESULTS>
                <RESULT eventid="1134" points="180" swimtime="00:00:42.50" resultid="1952" heatid="6991" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1194" points="211" swimtime="00:01:18.75" resultid="1953" heatid="7013" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="252" swimtime="00:00:42.20" resultid="1954" heatid="7056" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1316" points="130" swimtime="00:01:42.42" resultid="1955" heatid="7068" lane="6" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="217" swimtime="00:00:34.76" resultid="1956" heatid="7125" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1543" points="200" swimtime="00:01:40.01" resultid="1957" heatid="7158" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Renata" gender="F" lastname="Bastek" nation="POL" athleteid="1958">
              <RESULTS>
                <RESULT eventid="1119" points="247" swimtime="00:00:43.09" resultid="1959" heatid="6984" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1240" points="149" swimtime="00:00:47.23" resultid="1960" heatid="7031" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1453" points="290" swimtime="00:00:35.83" resultid="1961" heatid="7117" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Daniel" gender="M" lastname="Weselak" nation="POL" athleteid="1962">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. B /30-34/" eventid="1224" points="415" swimtime="00:02:29.46" resultid="1963" heatid="7029" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="389" swimtime="00:02:36.13" resultid="1964" heatid="7102" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:02:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="428" swimtime="00:01:06.06" resultid="1965" heatid="7111" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="326" swimtime="00:02:42.48" resultid="1966" heatid="7145" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="150" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Bartosz" gender="M" lastname="Kwestorowski" nation="POL" athleteid="1967">
              <RESULTS>
                <RESULT eventid="1224" points="433" swimtime="00:02:27.38" resultid="1968" heatid="7029" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="1969" heatid="7072" lane="7" entrytime="00:01:05.00" />
                <RESULT eventid="1406" points="514" swimtime="00:02:22.28" resultid="1970" heatid="7103" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="458" swimtime="00:02:25.11" resultid="1971" heatid="7146" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="529" swimtime="00:04:32.07" resultid="1972" heatid="7171" lane="2" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:01:02.52" />
                    <SPLIT distance="150" swimtime="00:01:37.17" />
                    <SPLIT distance="200" swimtime="00:02:12.25" />
                    <SPLIT distance="250" swimtime="00:02:47.32" />
                    <SPLIT distance="300" swimtime="00:03:22.88" />
                    <SPLIT distance="350" swimtime="00:03:57.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Aleksander" gender="M" lastname="Nawrat" nation="POL" athleteid="1973">
              <RESULTS>
                <RESULT eventid="1194" points="199" swimtime="00:01:20.27" resultid="1974" heatid="7012" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="167" swimtime="00:00:40.67" resultid="1975" heatid="7037" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="1976" heatid="7126" lane="1" entrytime="00:00:32.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" athleteid="1977">
              <RESULTS>
                <RESULT eventid="1119" points="140" swimtime="00:00:52.00" resultid="1978" heatid="6982" lane="4" entrytime="00:00:54.00" />
                <RESULT eventid="1271" points="193" swimtime="00:00:51.48" resultid="1979" heatid="7049" lane="1" entrytime="00:00:52.00" />
                <RESULT eventid="1453" points="158" swimtime="00:00:43.88" resultid="1980" heatid="7115" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" athleteid="1981">
              <RESULTS>
                <RESULT eventid="1134" points="79" swimtime="00:00:55.88" resultid="1982" heatid="6989" lane="3" entrytime="00:00:48.50" />
                <RESULT eventid="1256" points="127" swimtime="00:00:44.52" resultid="1983" heatid="7038" lane="0" entrytime="00:00:38.50" />
                <RESULT eventid="1468" points="155" swimtime="00:00:38.92" resultid="1984" heatid="7124" lane="2" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Daniel" gender="M" lastname="Hoszczewski" nation="POL" athleteid="1985">
              <RESULTS>
                <RESULT eventid="1194" points="430" swimtime="00:01:02.13" resultid="1986" heatid="7020" lane="2" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="340" swimtime="00:00:32.13" resultid="1987" heatid="7044" lane="0" entrytime="00:00:29.99" />
                <RESULT eventid="1468" points="427" swimtime="00:00:27.76" resultid="1988" heatid="7136" lane="8" entrytime="00:00:25.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1164" points="239" swimtime="00:02:30.55" resultid="1990" heatid="7000" lane="1" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:57.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1923" number="1" />
                    <RELAYPOSITION athleteid="1951" number="2" />
                    <RELAYPOSITION athleteid="1981" number="3" />
                    <RELAYPOSITION athleteid="1908" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1164" points="416" swimtime="00:02:05.15" resultid="1991" heatid="7001" lane="6" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="150" swimtime="00:01:38.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1967" number="1" />
                    <RELAYPOSITION athleteid="1918" number="2" />
                    <RELAYPOSITION athleteid="1962" number="3" />
                    <RELAYPOSITION athleteid="1985" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1346" points="460" swimtime="00:01:49.89" resultid="1993" heatid="7076" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.97" />
                    <SPLIT distance="100" swimtime="00:00:55.13" />
                    <SPLIT distance="150" swimtime="00:01:23.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1967" number="1" />
                    <RELAYPOSITION athleteid="1962" number="2" />
                    <RELAYPOSITION athleteid="1918" number="3" />
                    <RELAYPOSITION athleteid="1985" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="6">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. E /240-279/" eventid="1346" points="242" swimtime="00:02:16.12" resultid="1994" heatid="7075" lane="0" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1951" number="1" />
                    <RELAYPOSITION athleteid="1908" number="2" />
                    <RELAYPOSITION athleteid="1934" number="3" />
                    <RELAYPOSITION athleteid="1892" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. E /240-279/" eventid="1149" points="232" swimtime="00:02:52.50" resultid="1989" heatid="6998" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:31.40" />
                    <SPLIT distance="150" swimtime="00:02:12.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1958" number="1" />
                    <RELAYPOSITION athleteid="1945" number="2" />
                    <RELAYPOSITION athleteid="1928" number="3" />
                    <RELAYPOSITION athleteid="1937" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1331" points="229" swimtime="00:02:38.03" resultid="1992" heatid="7073" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1937" number="1" />
                    <RELAYPOSITION athleteid="1977" number="2" />
                    <RELAYPOSITION athleteid="1928" number="3" />
                    <RELAYPOSITION athleteid="1958" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1513" status="DNF" swimtime="00:00:00.00" resultid="1995" heatid="7148" lane="7" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1941" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1977" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="1981" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="1937" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1513" points="153" swimtime="00:02:54.45" resultid="1996" heatid="7148" lane="2" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:29.02" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1958" number="1" />
                    <RELAYPOSITION athleteid="1898" number="2" />
                    <RELAYPOSITION athleteid="1902" number="3" />
                    <RELAYPOSITION athleteid="1951" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3283" heatid="7148" lane="6" entrytime="00:02:49.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1958" number="1" />
                    <RELAYPOSITION athleteid="1898" number="2" />
                    <RELAYPOSITION athleteid="1902" number="3" />
                    <RELAYPOSITION athleteid="1951" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MABOL" name="Klub Pływacki Masters Bolesławiec" nation="POL" region="DOL">
          <CONTACT email="sekretarz-masters@o2.pl" name="Marta Satoła" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="2036">
              <RESULTS>
                <RESULT eventid="1134" points="120" swimtime="00:00:48.72" resultid="2037" heatid="6989" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1224" points="60" swimtime="00:04:43.98" resultid="2038" heatid="7025" lane="4" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.72" />
                    <SPLIT distance="100" swimtime="00:02:08.99" />
                    <SPLIT distance="150" swimtime="00:03:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="109" swimtime="00:01:48.59" resultid="2039" heatid="7067" lane="5" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="96" swimtime="00:04:08.69" resultid="2040" heatid="7096" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.85" />
                    <SPLIT distance="100" swimtime="00:02:00.35" />
                    <SPLIT distance="150" swimtime="00:03:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="58" swimtime="00:02:08.63" resultid="2041" heatid="7106" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="104" swimtime="00:03:57.69" resultid="2042" heatid="7142" lane="9" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.67" />
                    <SPLIT distance="100" swimtime="00:01:59.82" />
                    <SPLIT distance="150" swimtime="00:03:00.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-25" firstname="Fryderyk" gender="M" lastname="Popieliński" nation="POL" athleteid="2043">
              <RESULTS>
                <RESULT eventid="1104" points="279" swimtime="00:03:14.67" resultid="2044" heatid="6977" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:33.25" />
                    <SPLIT distance="150" swimtime="00:02:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="134" swimtime="00:03:37.43" resultid="2045" heatid="7026" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:41.42" />
                    <SPLIT distance="150" swimtime="00:02:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="268" swimtime="00:02:38.17" resultid="2046" heatid="7087" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="241" swimtime="00:03:03.14" resultid="2047" heatid="7097" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:21.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G-9 - Ukończenie wyścigu nie w położeniu na plecach" eventid="1498" status="DSQ" swimtime="00:03:14.71" resultid="2048" heatid="7143" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:33.72" />
                    <SPLIT distance="150" swimtime="00:02:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="235" swimtime="00:05:56.42" resultid="2049" heatid="7170" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:03.48" />
                    <SPLIT distance="200" swimtime="00:02:50.12" />
                    <SPLIT distance="250" swimtime="00:03:36.76" />
                    <SPLIT distance="300" swimtime="00:04:24.40" />
                    <SPLIT distance="350" swimtime="00:05:11.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-11" firstname="Henryk" gender="M" lastname="Kopaniecki" nation="POL" athleteid="2050">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="2051" heatid="6977" lane="0" entrytime="00:03:20.00" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2052" heatid="7026" lane="2" entrytime="00:03:30.00" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="2053" heatid="7086" lane="5" entrytime="00:02:35.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2055" heatid="7143" lane="3" entrytime="00:03:10.00" />
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="2056" heatid="7170" lane="3" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASBYD" name="Astoria Bydgoszcz" nation="POL" region="KUJ">
          <CONTACT email="sikoreczka7@o2.pl" name="Sikorska Małgorzata" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Kawecki" nation="POL" athleteid="2058">
              <RESULTS>
                <RESULT eventid="1104" points="258" swimtime="00:03:19.75" resultid="2059" heatid="6978" lane="9" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:34.59" />
                    <SPLIT distance="150" swimtime="00:02:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="151" swimtime="00:03:29.24" resultid="2060" heatid="7027" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                    <SPLIT distance="100" swimtime="00:01:37.65" />
                    <SPLIT distance="150" swimtime="00:02:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="224" swimtime="00:00:43.85" resultid="2061" heatid="7057" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2062" heatid="7099" lane="6" entrytime="00:02:52.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2063" heatid="7144" lane="6" entrytime="00:02:55.00" />
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="2064" heatid="7170" lane="7" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIGLI" name="Sikret Gliwice" nation="POL" region="SLA">
          <CONTACT city="GLIWICE" email="J.ZAGALA@ECOTRADE.PL" name="ZAGAŁA JOANNA" phone="601427257" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-24" firstname="JOANNA" gender="F" lastname="ZAGAŁA" nation="POL" athleteid="2264">
              <RESULTS>
                <RESULT eventid="1058" points="175" swimtime="00:04:10.11" resultid="2265" heatid="6971" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.42" />
                    <SPLIT distance="100" swimtime="00:02:01.33" />
                    <SPLIT distance="150" swimtime="00:03:05.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="155" swimtime="00:00:50.28" resultid="2266" heatid="6982" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1271" points="196" swimtime="00:00:51.29" resultid="2267" heatid="7048" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="1391" points="144" swimtime="00:04:00.65" resultid="2268" heatid="7092" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                    <SPLIT distance="100" swimtime="00:01:59.46" />
                    <SPLIT distance="150" swimtime="00:03:05.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="216" swimtime="00:00:39.49" resultid="2269" heatid="7115" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2270" heatid="7151" lane="4" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="ZOFIA" gender="F" lastname="DĄBROWSKA" nation="POL" athleteid="2271">
              <RESULTS>
                <RESULT eventid="1179" points="162" swimtime="00:01:35.51" resultid="2272" heatid="7003" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="127" swimtime="00:00:49.80" resultid="2273" heatid="7031" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="1391" points="117" swimtime="00:04:17.59" resultid="2274" heatid="7092" lane="8" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                    <SPLIT distance="100" swimtime="00:02:11.04" />
                    <SPLIT distance="150" swimtime="00:03:17.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="190" swimtime="00:00:41.24" resultid="2275" heatid="7116" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1558" points="134" swimtime="00:07:46.76" resultid="2276" heatid="7164" lane="2" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                    <SPLIT distance="100" swimtime="00:01:51.80" />
                    <SPLIT distance="150" swimtime="00:02:53.31" />
                    <SPLIT distance="200" swimtime="00:03:52.81" />
                    <SPLIT distance="250" swimtime="00:04:53.86" />
                    <SPLIT distance="300" swimtime="00:05:53.52" />
                    <SPLIT distance="350" swimtime="00:06:53.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-14" firstname="DANUTA" gender="F" lastname="ZIARKO" nation="POL" athleteid="2277">
              <RESULTS>
                <RESULT eventid="1119" points="185" swimtime="00:00:47.47" resultid="2278" heatid="6984" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1209" points="145" swimtime="00:03:51.58" resultid="2279" heatid="7024" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="100" swimtime="00:01:47.46" />
                    <SPLIT distance="150" swimtime="00:02:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="283" swimtime="00:00:38.15" resultid="2280" heatid="7033" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1361" points="267" swimtime="00:02:55.30" resultid="2281" heatid="7079" lane="4" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="198" swimtime="00:01:36.18" resultid="2282" heatid="7104" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="237" swimtime="00:06:26.09" resultid="2283" heatid="7166" lane="8" entrytime="00:06:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                    <SPLIT distance="100" swimtime="00:01:31.19" />
                    <SPLIT distance="150" swimtime="00:02:20.38" />
                    <SPLIT distance="200" swimtime="00:03:10.08" />
                    <SPLIT distance="250" swimtime="00:04:00.45" />
                    <SPLIT distance="300" swimtime="00:04:50.85" />
                    <SPLIT distance="350" swimtime="00:05:41.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03001" name="MUKP Just Swim Jelenia Góra" nation="POL" region="DOL">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz" phone="509071929" zip="58-506" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-07" firstname="Wojciech" gender="M" lastname="Woźny" nation="POL" license="M031-0120003" athleteid="2291">
              <RESULTS>
                <RESULT eventid="1134" points="280" swimtime="00:00:36.73" resultid="2292" heatid="6994" lane="1" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1194" points="351" swimtime="00:01:06.47" resultid="2293" heatid="7017" lane="9" entrytime="00:01:06.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2294" heatid="7055" lane="5" entrytime="00:00:42.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="Waszkewicz" nation="POL" license="M0300120009" athleteid="2295">
              <RESULTS>
                <RESULT eventid="1256" points="586" swimtime="00:00:26.80" resultid="2296" heatid="7046" lane="3" entrytime="00:00:25.91" />
                <RESULT eventid="1468" points="603" swimtime="00:00:24.75" resultid="2297" heatid="7136" lane="3" entrytime="00:00:24.27" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VIJOZ" name="UKS Victoria Józefów" nation="POL" region="MAZ">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1980-11-08" firstname="Alicja" gender="F" lastname="Kowalczyk-kędzierska" nation="POL" athleteid="2299">
              <RESULTS>
                <RESULT eventid="1119" points="342" swimtime="00:00:38.66" resultid="2300" heatid="6985" lane="5" entrytime="00:00:38.65" />
                <RESULT eventid="1179" points="299" swimtime="00:01:17.80" resultid="2301" heatid="7006" lane="3" entrytime="00:01:16.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="352" swimtime="00:00:35.50" resultid="2302" heatid="7033" lane="3" entrytime="00:00:36.54" />
                <RESULT eventid="1301" points="309" swimtime="00:01:25.90" resultid="2303" heatid="7064" lane="4" entrytime="00:01:25.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="258" swimtime="00:01:27.98" resultid="2304" heatid="7105" lane="1" entrytime="00:01:30.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="285" swimtime="00:03:09.56" resultid="2305" heatid="7139" lane="9" entrytime="00:03:10.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:23.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="2306">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="2307" heatid="6978" lane="4" entrytime="00:03:08.05" />
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="2308" heatid="7017" lane="1" entrytime="00:01:06.02" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="2309" heatid="7056" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2310" heatid="7099" lane="3" entrytime="00:02:50.09" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="2311" heatid="7159" lane="8" entrytime="00:01:28.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZKAT" name="AZS AWF Katowice" nation="POL" region="SLA">
          <CONTACT city="Gliwice" email="tomasz-czermak@wp.pl" name="Tomasz Czermak" phone="515 585 011" street="Żeromskiego 84/7" zip="44-119" />
          <ATHLETES>
            <ATHLETE birthdate="1991-09-13" firstname="Tomasz" gender="M" lastname="Czermak" nation="POL" license="S00611200197" athleteid="2320">
              <RESULTS>
                <RESULT eventid="1104" points="582" swimtime="00:02:32.46" resultid="2321" heatid="6980" lane="5" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="410" swimtime="00:02:30.09" resultid="2322" heatid="7029" lane="9" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="596" swimtime="00:00:31.68" resultid="2323" heatid="7061" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1406" points="518" swimtime="00:02:21.94" resultid="2324" heatid="7103" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="575" swimtime="00:01:10.43" resultid="2325" heatid="7163" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="505" swimtime="00:04:36.25" resultid="2326" heatid="7174" lane="7" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:40.74" />
                    <SPLIT distance="200" swimtime="00:02:15.87" />
                    <SPLIT distance="250" swimtime="00:02:51.66" />
                    <SPLIT distance="300" swimtime="00:03:27.32" />
                    <SPLIT distance="350" swimtime="00:04:02.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KOKRA" name="Masters Korona Kraków" nation="POL" region="MAL">
          <CONTACT email="masterskorona@wp.pl" internet="www.masterskorona.pl" name="mariola Kuliś" phone="500677133" state="KR" />
          <ATHLETES>
            <ATHLETE birthdate="1933-04-07" firstname="Tadeusz" gender="M" lastname="Banach" nation="POL" athleteid="2328">
              <RESULTS>
                <RESULT eventid="1134" points="30" swimtime="00:01:16.82" resultid="2329" heatid="6987" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1468" points="25" swimtime="00:01:10.74" resultid="2330" heatid="7121" lane="7" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="2331">
              <RESULTS>
                <RESULT eventid="1194" points="455" swimtime="00:01:00.99" resultid="2332" heatid="7020" lane="6" entrytime="00:00:59.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="361" swimtime="00:00:37.45" resultid="2333" heatid="7059" lane="5" entrytime="00:00:35.12" />
                <RESULT eventid="1376" points="342" swimtime="00:02:25.78" resultid="2334" heatid="7088" lane="9" entrytime="00:02:21.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:08.94" />
                    <SPLIT distance="150" swimtime="00:01:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="461" swimtime="00:00:27.05" resultid="2335" heatid="7135" lane="2" entrytime="00:00:26.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-04-24" firstname="Krzysztof" gender="M" lastname="Chołda" nation="POL" athleteid="2337">
              <RESULTS>
                <RESULT eventid="1134" points="184" swimtime="00:00:42.24" resultid="2338" heatid="6991" lane="6" entrytime="00:00:41.05" />
                <RESULT eventid="1194" points="265" swimtime="00:01:13.00" resultid="2339" heatid="7015" lane="7" entrytime="00:01:10.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="264" swimtime="00:00:41.55" resultid="2340" heatid="7054" lane="5" entrytime="00:00:44.90" />
                <RESULT eventid="1406" points="217" swimtime="00:03:09.70" resultid="2341" heatid="7098" lane="8" entrytime="00:03:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:33.72" />
                    <SPLIT distance="150" swimtime="00:02:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="252" swimtime="00:00:33.08" resultid="2342" heatid="7127" lane="7" entrytime="00:00:31.14" />
                <RESULT eventid="1573" points="211" swimtime="00:06:09.28" resultid="2343" heatid="7170" lane="0" entrytime="00:05:55.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:02:08.81" />
                    <SPLIT distance="200" swimtime="00:02:55.93" />
                    <SPLIT distance="250" swimtime="00:03:44.35" />
                    <SPLIT distance="300" swimtime="00:04:33.19" />
                    <SPLIT distance="350" swimtime="00:05:22.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="Data" nation="POL" athleteid="2344">
              <RESULTS>
                <RESULT eventid="1104" points="185" swimtime="00:03:43.35" resultid="2345" heatid="6977" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:43.51" />
                    <SPLIT distance="150" swimtime="00:02:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="198" swimtime="00:01:20.46" resultid="2346" heatid="7014" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="196" swimtime="00:00:45.87" resultid="2347" heatid="7055" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1406" points="154" swimtime="00:03:32.23" resultid="2348" heatid="7098" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                    <SPLIT distance="100" swimtime="00:01:42.84" />
                    <SPLIT distance="150" swimtime="00:02:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="197" swimtime="00:01:40.53" resultid="2349" heatid="7158" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="179" swimtime="00:06:30.18" resultid="2350" heatid="7169" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                    <SPLIT distance="150" swimtime="00:02:16.67" />
                    <SPLIT distance="200" swimtime="00:03:07.61" />
                    <SPLIT distance="250" swimtime="00:03:59.30" />
                    <SPLIT distance="300" swimtime="00:04:51.02" />
                    <SPLIT distance="350" swimtime="00:05:42.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-07" firstname="Robert" gender="M" lastname="Grela" nation="POL" athleteid="2351">
              <RESULTS>
                <RESULT eventid="1224" points="338" swimtime="00:02:39.93" resultid="2352" heatid="7029" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="415" swimtime="00:00:30.05" resultid="2353" heatid="7045" lane="0" entrytime="00:00:28.00" />
                <RESULT comment="O-4 - Przedwczwsny start" eventid="1438" status="DSQ" swimtime="00:01:08.18" resultid="2354" heatid="7111" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Mariusz" gender="M" lastname="Kaliszyk" nation="POL" athleteid="2355">
              <RESULTS>
                <RESULT eventid="1134" points="413" swimtime="00:00:32.28" resultid="2356" heatid="6996" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1194" points="428" swimtime="00:01:02.21" resultid="2357" heatid="7018" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="354" swimtime="00:01:13.38" resultid="2358" heatid="7070" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2359" heatid="7101" lane="8" entrytime="00:02:45.00" />
                <RESULT eventid="1468" points="396" swimtime="00:00:28.46" resultid="2360" heatid="7134" lane="0" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-11" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="2361">
              <RESULTS>
                <RESULT eventid="1134" points="34" swimtime="00:01:13.65" resultid="2362" heatid="6987" lane="6" entrytime="00:01:11.00" />
                <RESULT eventid="1194" points="82" swimtime="00:01:47.84" resultid="2363" heatid="7010" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="32" swimtime="00:02:43.09" resultid="2364" heatid="7066" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="104" swimtime="00:00:44.33" resultid="2365" heatid="7122" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2366" heatid="7141" lane="0" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="2367">
              <RESULTS>
                <RESULT eventid="1104" points="321" swimtime="00:03:05.75" resultid="2368" heatid="6979" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:15.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="410" swimtime="00:00:30.18" resultid="2369" heatid="7044" lane="8" entrytime="00:00:29.70" />
                <RESULT eventid="1286" points="397" swimtime="00:00:36.28" resultid="2370" heatid="7059" lane="6" entrytime="00:00:35.80" />
                <RESULT eventid="1543" points="360" swimtime="00:01:22.33" resultid="2371" heatid="7162" lane="9" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="2372">
              <RESULTS>
                <RESULT eventid="1194" points="234" swimtime="00:01:16.06" resultid="2373" heatid="7013" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="70" swimtime="00:04:29.90" resultid="2374" heatid="7026" lane="9" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.62" />
                    <SPLIT distance="100" swimtime="00:02:07.70" />
                    <SPLIT distance="150" swimtime="00:03:18.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="187" swimtime="00:02:58.20" resultid="2375" heatid="7084" lane="4" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="135" swimtime="00:03:41.74" resultid="2376" heatid="7096" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:53.60" />
                    <SPLIT distance="150" swimtime="00:02:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="105" swimtime="00:01:45.37" resultid="2377" heatid="7107" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="159" swimtime="00:06:45.74" resultid="2378" heatid="7169" lane="8" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                    <SPLIT distance="100" swimtime="00:01:38.09" />
                    <SPLIT distance="150" swimtime="00:02:30.97" />
                    <SPLIT distance="200" swimtime="00:03:25.78" />
                    <SPLIT distance="250" swimtime="00:04:18.35" />
                    <SPLIT distance="300" swimtime="00:05:12.82" />
                    <SPLIT distance="350" swimtime="00:06:04.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="2379">
              <RESULTS>
                <RESULT eventid="1134" points="294" swimtime="00:00:36.13" resultid="2380" heatid="6994" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1256" points="392" swimtime="00:00:30.63" resultid="2381" heatid="7040" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1316" points="276" swimtime="00:01:19.69" resultid="2382" heatid="7070" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="2383" heatid="7109" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1498" points="244" swimtime="00:02:59.05" resultid="2384" heatid="7144" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:26.76" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="2385">
              <RESULTS>
                <RESULT eventid="1224" points="329" swimtime="00:02:41.49" resultid="2386" heatid="7028" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="363" swimtime="00:00:31.44" resultid="2387" heatid="7042" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1438" points="373" swimtime="00:01:09.17" resultid="2388" heatid="7111" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="346" swimtime="00:05:13.37" resultid="2389" heatid="7173" lane="8" entrytime="00:04:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:52.76" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:13.78" />
                    <SPLIT distance="300" swimtime="00:03:54.46" />
                    <SPLIT distance="350" swimtime="00:04:34.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Robert" gender="M" lastname="Trzos" nation="POL" athleteid="2390">
              <RESULTS>
                <RESULT eventid="1104" points="314" swimtime="00:03:07.24" resultid="2391" heatid="6979" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:29.12" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="189" swimtime="00:01:30.47" resultid="2392" heatid="7070" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="271" swimtime="00:01:30.50" resultid="2393" heatid="7161" lane="0" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="2394">
              <RESULTS>
                <RESULT eventid="1119" points="235" swimtime="00:00:43.83" resultid="2395" heatid="6983" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1301" points="208" swimtime="00:01:38.05" resultid="2396" heatid="7063" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="183" swimtime="00:03:18.90" resultid="2397" heatid="7078" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:35.73" />
                    <SPLIT distance="150" swimtime="00:02:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="211" swimtime="00:03:31.80" resultid="2398" heatid="7092" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:42.28" />
                    <SPLIT distance="150" swimtime="00:02:43.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="210" swimtime="00:03:29.87" resultid="2399" heatid="7137" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                    <SPLIT distance="100" swimtime="00:01:44.38" />
                    <SPLIT distance="150" swimtime="00:02:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="186" swimtime="00:06:58.75" resultid="2400" heatid="7165" lane="8" entrytime="00:07:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:37.07" />
                    <SPLIT distance="150" swimtime="00:02:30.20" />
                    <SPLIT distance="200" swimtime="00:03:25.05" />
                    <SPLIT distance="250" swimtime="00:04:19.22" />
                    <SPLIT distance="300" swimtime="00:05:13.25" />
                    <SPLIT distance="350" swimtime="00:06:07.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Koźmin" nation="POL" athleteid="2401">
              <RESULTS>
                <RESULT eventid="1058" points="141" swimtime="00:04:28.93" resultid="2402" heatid="6971" lane="0" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.89" />
                    <SPLIT distance="100" swimtime="00:02:07.27" />
                    <SPLIT distance="150" swimtime="00:03:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="174" swimtime="00:00:53.36" resultid="2403" heatid="7049" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1391" points="111" swimtime="00:04:22.25" resultid="2404" heatid="7091" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.79" />
                    <SPLIT distance="100" swimtime="00:02:08.66" />
                    <SPLIT distance="150" swimtime="00:03:21.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="143" swimtime="00:02:02.97" resultid="2405" heatid="7152" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="2406">
              <RESULTS>
                <RESULT eventid="1119" points="380" swimtime="00:00:37.33" resultid="2407" heatid="6983" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1179" points="383" swimtime="00:01:11.67" resultid="2408" heatid="7007" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. E /45-49/" eventid="1271" points="403" swimtime="00:00:40.33" resultid="2410" heatid="7051" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1453" points="401" swimtime="00:00:32.16" resultid="2411" heatid="7119" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="2412" heatid="7154" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1301" points="342" swimtime="00:01:23.10" resultid="5651" heatid="7065" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="2413">
              <RESULTS>
                <RESULT eventid="1058" points="318" swimtime="00:03:25.13" resultid="2414" heatid="6973" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:37.05" />
                    <SPLIT distance="150" swimtime="00:02:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="318" swimtime="00:00:43.65" resultid="2415" heatid="7050" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1528" points="295" swimtime="00:01:36.77" resultid="2416" heatid="7154" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="2417">
              <RESULTS>
                <RESULT eventid="1119" points="236" swimtime="00:00:43.75" resultid="2418" heatid="6981" lane="6" />
                <RESULT comment="Rekord Polski Masters w kat. G /55-59/" eventid="1209" points="140" swimtime="00:03:54.40" resultid="2419" heatid="7024" lane="3" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.44" />
                    <SPLIT distance="100" swimtime="00:01:51.70" />
                    <SPLIT distance="150" swimtime="00:02:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="214" swimtime="00:00:41.85" resultid="2420" heatid="7030" lane="1" />
                <RESULT eventid="1391" points="209" swimtime="00:03:32.31" resultid="2421" heatid="7093" lane="9" entrytime="00:03:40.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                    <SPLIT distance="100" swimtime="00:01:44.47" />
                    <SPLIT distance="150" swimtime="00:02:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat G /55-59/" eventid="1422" points="169" swimtime="00:01:41.39" resultid="2422" heatid="7104" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="156" swimtime="00:03:51.52" resultid="2423" heatid="7138" lane="0" entrytime="00:03:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.69" />
                    <SPLIT distance="100" swimtime="00:01:54.65" />
                    <SPLIT distance="150" swimtime="00:02:56.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="2424">
              <RESULTS>
                <RESULT eventid="1058" points="92" swimtime="00:05:09.57" resultid="2425" heatid="6970" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.18" />
                    <SPLIT distance="100" swimtime="00:02:29.57" />
                    <SPLIT distance="150" swimtime="00:03:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="69" swimtime="00:02:06.83" resultid="2426" heatid="7002" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="34" swimtime="00:01:16.74" resultid="2427" heatid="7030" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1391" points="51" swimtime="00:05:38.48" resultid="2428" heatid="7091" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.40" />
                    <SPLIT distance="100" swimtime="00:02:36.57" />
                    <SPLIT distance="150" swimtime="00:04:02.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="64" swimtime="00:00:59.29" resultid="2429" heatid="7114" lane="6" entrytime="00:01:06.00" />
                <RESULT eventid="1528" points="97" swimtime="00:02:20.24" resultid="2430" heatid="7151" lane="7" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="2431">
              <RESULTS>
                <RESULT eventid="1119" points="412" swimtime="00:00:36.34" resultid="2432" heatid="6986" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1271" points="354" swimtime="00:00:42.11" resultid="2433" heatid="7050" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1301" points="401" swimtime="00:01:18.76" resultid="2434" heatid="7065" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="366" swimtime="00:02:54.47" resultid="2435" heatid="7139" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="2436">
              <RESULTS>
                <RESULT eventid="1179" points="135" swimtime="00:01:41.47" resultid="2437" heatid="7003" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="78" swimtime="00:00:58.43" resultid="2438" heatid="7031" lane="9" entrytime="00:00:58.00" />
                <RESULT eventid="1361" points="114" swimtime="00:03:52.83" resultid="2439" heatid="7077" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:52.78" />
                    <SPLIT distance="150" swimtime="00:02:55.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="68" swimtime="00:02:16.98" resultid="2440" heatid="7104" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="2441">
              <RESULTS>
                <RESULT eventid="1179" points="312" swimtime="00:01:16.70" resultid="2442" heatid="7007" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="356" swimtime="00:00:35.37" resultid="2443" heatid="7034" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1391" points="327" swimtime="00:03:03.06" resultid="2444" heatid="7093" lane="5" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="336" swimtime="00:01:20.56" resultid="2445" heatid="7105" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="309" swimtime="00:05:53.46" resultid="2446" heatid="7167" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="150" swimtime="00:02:07.41" />
                    <SPLIT distance="200" swimtime="00:02:51.70" />
                    <SPLIT distance="250" swimtime="00:03:36.60" />
                    <SPLIT distance="300" swimtime="00:04:22.45" />
                    <SPLIT distance="350" swimtime="00:05:08.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="2447">
              <RESULTS>
                <RESULT eventid="1058" points="347" swimtime="00:03:19.29" resultid="2448" heatid="6973" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:33.32" />
                    <SPLIT distance="150" swimtime="00:02:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="272" swimtime="00:01:20.29" resultid="2449" heatid="7006" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="349" swimtime="00:00:42.29" resultid="2450" heatid="7050" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1453" points="274" swimtime="00:00:36.52" resultid="2451" heatid="7118" lane="1" entrytime="00:00:35.00" />
                <RESULT comment="Rekord Polski Masters w kat F /50-54/" eventid="1528" points="356" swimtime="00:01:30.91" resultid="2452" heatid="7153" lane="5" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-18" firstname="Jadwiga" gender="F" lastname="Gorecka" nation="POL" athleteid="2453">
              <RESULTS>
                <RESULT eventid="1119" points="201" swimtime="00:00:46.13" resultid="2454" heatid="6984" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1179" points="220" swimtime="00:01:26.13" resultid="2455" heatid="7006" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="208" swimtime="00:00:42.28" resultid="2456" heatid="7032" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1453" points="285" swimtime="00:00:36.02" resultid="2457" heatid="7118" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-16" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="2458">
              <RESULTS>
                <RESULT eventid="1058" points="129" swimtime="00:04:36.88" resultid="2459" heatid="6970" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.42" />
                    <SPLIT distance="100" swimtime="00:02:17.95" />
                    <SPLIT distance="150" swimtime="00:03:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="110" swimtime="00:00:56.33" resultid="2460" heatid="6983" lane="9" entrytime="00:00:53.58" />
                <RESULT eventid="1271" points="130" swimtime="00:00:58.69" resultid="2461" heatid="7048" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1301" points="85" swimtime="00:02:11.83" resultid="2462" heatid="7063" lane="2" entrytime="00:02:05.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="85" swimtime="00:04:43.82" resultid="2463" heatid="7137" lane="7" entrytime="00:04:58.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.32" />
                    <SPLIT distance="100" swimtime="00:02:21.74" />
                    <SPLIT distance="150" swimtime="00:03:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="115" swimtime="00:02:12.35" resultid="2464" heatid="7151" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kr C" number="3">
              <RESULTS>
                <RESULT eventid="1346" points="396" swimtime="00:01:55.52" resultid="2466" heatid="7075" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="100" swimtime="00:00:57.72" />
                    <SPLIT distance="150" swimtime="00:01:27.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2355" number="1" />
                    <RELAYPOSITION athleteid="2351" number="2" />
                    <RELAYPOSITION athleteid="2385" number="3" />
                    <RELAYPOSITION athleteid="2367" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1164" points="385" swimtime="00:02:08.39" resultid="2467" heatid="7000" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:38.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2355" number="1" />
                    <RELAYPOSITION athleteid="2367" number="2" />
                    <RELAYPOSITION athleteid="2351" number="3" />
                    <RELAYPOSITION athleteid="2385" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kr D" number="4">
              <RESULTS>
                <RESULT eventid="1164" points="252" swimtime="00:02:27.78" resultid="2472" heatid="7000" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2379" number="1" />
                    <RELAYPOSITION athleteid="2390" number="2" />
                    <RELAYPOSITION athleteid="2337" number="3" />
                    <RELAYPOSITION athleteid="2372" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kr E" number="9">
              <RESULTS>
                <RESULT eventid="1346" points="125" swimtime="00:02:49.66" resultid="2476" heatid="7074" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.69" />
                    <SPLIT distance="100" swimtime="00:01:45.04" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2328" number="1" />
                    <RELAYPOSITION athleteid="2337" number="2" />
                    <RELAYPOSITION athleteid="2372" number="3" />
                    <RELAYPOSITION athleteid="2379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kr D" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. D /200-239/" eventid="1331" points="353" swimtime="00:02:16.84" resultid="2468" heatid="7073" lane="5" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:42.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2406" number="1" />
                    <RELAYPOSITION athleteid="2441" number="2" />
                    <RELAYPOSITION athleteid="2417" number="3" />
                    <RELAYPOSITION athleteid="2447" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kat. D /200-239/" eventid="1149" points="347" swimtime="00:02:30.98" resultid="2469" heatid="6998" lane="5" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                    <SPLIT distance="150" swimtime="00:01:54.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2406" number="1" />
                    <RELAYPOSITION athleteid="2447" number="2" />
                    <RELAYPOSITION athleteid="2441" number="3" />
                    <RELAYPOSITION athleteid="2417" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kr B" number="2">
              <RESULTS>
                <RESULT eventid="1149" points="287" swimtime="00:02:40.80" resultid="2470" heatid="6998" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2431" number="1" />
                    <RELAYPOSITION athleteid="2413" number="2" />
                    <RELAYPOSITION athleteid="2453" number="3" />
                    <RELAYPOSITION athleteid="2394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1331" points="294" swimtime="00:02:25.44" resultid="2471" heatid="7073" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:52.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2394" number="1" />
                    <RELAYPOSITION athleteid="2413" number="2" />
                    <RELAYPOSITION athleteid="2453" number="3" />
                    <RELAYPOSITION athleteid="2431" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kr C" number="6">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat C /160-199/" eventid="1513" points="328" swimtime="00:02:15.40" resultid="2473" heatid="7149" lane="7" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:43.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2355" number="1" />
                    <RELAYPOSITION athleteid="2367" number="2" />
                    <RELAYPOSITION athleteid="2441" number="3" />
                    <RELAYPOSITION athleteid="2406" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kr D" number="7">
              <RESULTS>
                <RESULT eventid="1513" points="272" swimtime="00:02:24.06" resultid="2474" heatid="7149" lane="0" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:18.90" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2379" number="1" />
                    <RELAYPOSITION athleteid="2447" number="2" />
                    <RELAYPOSITION athleteid="2351" number="3" />
                    <RELAYPOSITION athleteid="2453" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kr E" number="8">
              <RESULTS>
                <RESULT eventid="1513" points="122" swimtime="00:03:07.95" resultid="2465" heatid="7148" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:40.89" />
                    <SPLIT distance="150" swimtime="00:02:23.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2417" number="1" />
                    <RELAYPOSITION athleteid="2401" number="2" />
                    <RELAYPOSITION athleteid="2372" number="3" />
                    <RELAYPOSITION athleteid="2361" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kr B" number="9">
              <RESULTS>
                <RESULT eventid="1513" points="276" swimtime="00:02:23.35" resultid="2475" heatid="7149" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:01:48.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2431" number="1" />
                    <RELAYPOSITION athleteid="2390" number="2" />
                    <RELAYPOSITION athleteid="2385" number="3" />
                    <RELAYPOSITION athleteid="2394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" name="Straz Miejska miasta kraków" nation="POL" region="KR">
          <CONTACT name="Jawień Krzysztof" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-12" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="2505">
              <RESULTS>
                <RESULT eventid="1104" points="391" swimtime="00:02:54.10" resultid="2506" heatid="6980" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:21.37" />
                    <SPLIT distance="150" swimtime="00:02:07.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="244" swimtime="00:02:58.31" resultid="2507" heatid="7028" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:17.01" />
                    <SPLIT distance="150" swimtime="00:02:06.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="401" swimtime="00:00:36.16" resultid="2508" heatid="7060" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1376" points="291" swimtime="00:02:33.88" resultid="2509" heatid="7087" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:55.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2510" heatid="7141" lane="5" entrytime="00:04:00.00" />
                <RESULT eventid="1543" points="388" swimtime="00:01:20.30" resultid="2511" heatid="7162" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" name="Masters Kraśnik" nation="POL" region="LBL">
          <CONTACT city="Kraśnik" email="jurek@krasnik. info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601 69 89 77" state="LUB." street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="2513">
              <RESULTS>
                <RESULT eventid="1104" points="159" swimtime="00:03:54.61" resultid="2514" heatid="6975" lane="1" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:52.77" />
                    <SPLIT distance="150" swimtime="00:02:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="111" swimtime="00:00:46.54" resultid="2515" heatid="7036" lane="4" entrytime="00:00:47.30" />
                <RESULT eventid="1286" points="175" swimtime="00:00:47.65" resultid="2516" heatid="7053" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1438" points="76" swimtime="00:01:57.15" resultid="2517" heatid="7107" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="2518">
              <RESULTS>
                <RESULT eventid="1104" points="296" swimtime="00:03:11.01" resultid="2519" heatid="6977" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:32.34" />
                    <SPLIT distance="150" swimtime="00:02:22.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="319" swimtime="00:00:39.00" resultid="2520" heatid="7057" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1543" points="293" swimtime="00:01:28.12" resultid="2521" heatid="7160" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="2522">
              <RESULTS>
                <RESULT eventid="1134" points="224" swimtime="00:00:39.55" resultid="2523" heatid="6992" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="2524" heatid="7014" lane="1" entrytime="00:01:14.00" />
                <RESULT eventid="1316" points="206" swimtime="00:01:27.86" resultid="2526" heatid="7068" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="2527" heatid="7127" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1498" points="170" swimtime="00:03:21.89" resultid="2528" heatid="7143" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                    <SPLIT distance="150" swimtime="00:02:35.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-30" firstname="Bartłomiej" gender="M" lastname="Sieczyński" nation="POL" athleteid="5652">
              <RESULTS>
                <RESULT eventid="1194" points="298" swimtime="00:01:10.23" resultid="5653" heatid="7016" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="229" swimtime="00:00:36.66" resultid="5654" heatid="7039" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1376" points="284" swimtime="00:02:35.00" resultid="5655" heatid="7088" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="309" swimtime="00:00:30.91" resultid="5656" heatid="7128" lane="7" entrytime="00:00:30.70" />
                <RESULT eventid="1573" points="282" swimtime="00:05:35.30" resultid="5657" heatid="7171" lane="3" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:56.36" />
                    <SPLIT distance="200" swimtime="00:02:39.29" />
                    <SPLIT distance="250" swimtime="00:03:23.32" />
                    <SPLIT distance="300" swimtime="00:04:07.97" />
                    <SPLIT distance="350" swimtime="00:04:52.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRLOD" name="MKS &quot;Trójka&quot; Łódź" nation="POL" region="LO">
          <CONTACT city="Łódź" name="Międzyszkolny Klub Sportowy" state="LOD" street="Sienkiewicza 46" zip="90-012" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-08" firstname="Marcin" gender="M" lastname="Babuchowski" nation="POL" athleteid="2545">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat A /25-29/" eventid="1194" points="735" swimtime="00:00:51.96" resultid="2546" heatid="7022" lane="4" entrytime="00:00:52.40" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters w kat. A /25-29/" eventid="1256" points="732" swimtime="00:00:24.88" resultid="2547" heatid="7046" lane="4" entrytime="00:00:24.58" entrycourse="LCM" />
                <RESULT eventid="1316" points="648" swimtime="00:01:00.00" resultid="2548" heatid="7072" lane="5" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat A /25-29/" eventid="1438" points="754" swimtime="00:00:54.73" resultid="2549" heatid="7112" lane="4" entrytime="00:00:53.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="645" swimtime="00:00:24.20" resultid="2550" heatid="7136" lane="2" entrytime="00:00:25.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MABIA" name="Masters Białystok" nation="POL" region="PDL">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko Wojciech" phone="797309140" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="2552">
              <RESULTS>
                <RESULT eventid="1119" points="310" swimtime="00:00:39.95" resultid="2553" heatid="6985" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1179" points="348" swimtime="00:01:13.99" resultid="2554" heatid="7007" lane="1" entrytime="00:01:13.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="301" swimtime="00:01:26.69" resultid="2555" heatid="7064" lane="2" entrytime="00:01:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="315" swimtime="00:02:45.93" resultid="2556" heatid="7080" lane="5" entrytime="00:02:44.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="371" swimtime="00:00:33.00" resultid="2557" heatid="7119" lane="0" entrytime="00:00:33.10" />
                <RESULT eventid="1483" points="283" swimtime="00:03:10.02" resultid="2558" heatid="7139" lane="8" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:02:21.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Bartek" gender="M" lastname="Bogdanowicz" nation="POL" athleteid="2559">
              <RESULTS>
                <RESULT eventid="1134" points="414" swimtime="00:00:32.23" resultid="2560" heatid="6995" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1316" points="396" swimtime="00:01:10.69" resultid="2561" heatid="7071" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="330" swimtime="00:02:41.90" resultid="2562" heatid="7145" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:02.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Hubert" gender="M" lastname="Milewski" nation="POL" athleteid="2563">
              <RESULTS>
                <RESULT eventid="1194" points="324" swimtime="00:01:08.27" resultid="2564" heatid="7015" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="346" swimtime="00:00:37.98" resultid="2565" heatid="7059" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1406" points="260" swimtime="00:02:58.55" resultid="2566" heatid="7100" lane="7" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:26.02" />
                    <SPLIT distance="150" swimtime="00:02:16.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="335" swimtime="00:00:30.08" resultid="2567" heatid="7127" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1543" status="DNF" swimtime="00:00:00.00" resultid="2568" heatid="7160" lane="1" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="2569">
              <RESULTS>
                <RESULT eventid="1179" points="409" swimtime="00:01:10.10" resultid="2570" heatid="7007" lane="4" entrytime="00:01:09.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="404" swimtime="00:02:32.73" resultid="2571" heatid="7081" lane="0" entrytime="00:02:32.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="412" swimtime="00:05:21.17" resultid="2572" heatid="7167" lane="3" entrytime="00:05:17.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:01:55.46" />
                    <SPLIT distance="200" swimtime="00:02:36.33" />
                    <SPLIT distance="250" swimtime="00:03:17.67" />
                    <SPLIT distance="300" swimtime="00:03:59.19" />
                    <SPLIT distance="350" swimtime="00:04:41.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="2573">
              <RESULTS>
                <RESULT eventid="1134" points="276" swimtime="00:00:36.90" resultid="2574" heatid="6992" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1194" points="210" swimtime="00:01:18.87" resultid="2575" heatid="7013" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="230" swimtime="00:01:24.66" resultid="2576" heatid="7069" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="180" swimtime="00:03:00.33" resultid="2577" heatid="7084" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="235" swimtime="00:00:33.87" resultid="2578" heatid="7126" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1498" points="199" swimtime="00:03:11.45" resultid="2579" heatid="7143" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:30.81" />
                    <SPLIT distance="150" swimtime="00:02:21.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="2580">
              <RESULTS>
                <RESULT eventid="1179" points="197" swimtime="00:01:29.39" resultid="2581" heatid="7005" lane="0" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="191" swimtime="00:03:15.95" resultid="2582" heatid="7079" lane="0" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:02:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="2583" heatid="7117" lane="2" entrytime="00:00:36.50" />
                <RESULT eventid="1558" points="168" swimtime="00:07:13.00" resultid="2584" heatid="7165" lane="1" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:36.00" />
                    <SPLIT distance="150" swimtime="00:02:31.11" />
                    <SPLIT distance="200" swimtime="00:03:27.15" />
                    <SPLIT distance="250" swimtime="00:04:24.35" />
                    <SPLIT distance="300" swimtime="00:05:22.16" />
                    <SPLIT distance="350" swimtime="00:06:19.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="2585">
              <RESULTS>
                <RESULT eventid="1104" points="259" swimtime="00:03:19.66" resultid="2586" heatid="6977" lane="4" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                    <SPLIT distance="150" swimtime="00:02:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="291" swimtime="00:00:33.83" resultid="2587" heatid="7035" lane="5" />
                <RESULT eventid="1286" points="379" swimtime="00:00:36.85" resultid="2588" heatid="7058" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1468" points="239" swimtime="00:00:33.69" resultid="2589" heatid="7127" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1543" points="336" swimtime="00:01:24.24" resultid="2590" heatid="7160" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="2591">
              <RESULTS>
                <RESULT eventid="1194" points="438" swimtime="00:01:01.73" resultid="2592" heatid="7019" lane="7" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="391" swimtime="00:00:30.67" resultid="2593" heatid="7042" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="1406" points="364" swimtime="00:02:39.57" resultid="2594" heatid="7101" lane="5" entrytime="00:02:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:02:02.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="368" swimtime="00:01:09.49" resultid="2595" heatid="7111" lane="8" entrytime="00:01:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="388" swimtime="00:00:28.65" resultid="2596" heatid="7130" lane="6" entrytime="00:00:28.75" />
                <RESULT eventid="1498" points="301" swimtime="00:02:46.90" resultid="2597" heatid="7145" lane="2" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:02:05.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEPL" name="K.S. niezrzeszeni.pl" nation="POL" region="MAZ">
          <CONTACT email="niezrzeszenipl@gmail.com" internet="niezrzeszeni.pl" name="Wawer Matylda Katarzyna" phone="501701359" />
          <ATHLETES>
            <ATHLETE birthdate="1960-07-16" firstname="Matylda Katarzyna" gender="F" lastname="Wawer" nation="POL" athleteid="2602">
              <RESULTS>
                <RESULT eventid="1179" points="233" swimtime="00:01:24.52" resultid="2603" heatid="7005" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="150" swimtime="00:00:47.16" resultid="2604" heatid="7032" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1361" points="150" swimtime="00:03:32.26" resultid="2605" heatid="7079" lane="9" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:43.05" />
                    <SPLIT distance="150" swimtime="00:02:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="284" swimtime="00:00:36.10" resultid="2606" heatid="7117" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1558" points="133" swimtime="00:07:48.02" resultid="2607" heatid="7165" lane="9" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:46.60" />
                    <SPLIT distance="150" swimtime="00:02:46.08" />
                    <SPLIT distance="200" swimtime="00:03:45.82" />
                    <SPLIT distance="250" swimtime="00:04:47.33" />
                    <SPLIT distance="300" swimtime="00:05:48.82" />
                    <SPLIT distance="350" swimtime="00:06:49.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="2608">
              <RESULTS>
                <RESULT eventid="1104" points="189" swimtime="00:03:41.74" resultid="2609" heatid="6976" lane="3" entrytime="00:03:29.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="100" swimtime="00:01:45.09" />
                    <SPLIT distance="150" swimtime="00:02:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="169" swimtime="00:01:24.76" resultid="2610" heatid="7012" lane="7" entrytime="00:01:20.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="203" swimtime="00:00:45.35" resultid="2611" heatid="7055" lane="1" entrytime="00:00:43.84" />
                <RESULT eventid="1376" points="164" swimtime="00:03:06.30" resultid="2612" heatid="7084" lane="6" entrytime="00:02:59.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:30.63" />
                    <SPLIT distance="150" swimtime="00:02:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="178" swimtime="00:00:37.16" resultid="2613" heatid="7124" lane="7" entrytime="00:00:35.53" />
                <RESULT eventid="1573" points="177" swimtime="00:06:31.82" resultid="2614" heatid="7169" lane="3" entrytime="00:06:17.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="150" swimtime="00:02:21.40" />
                    <SPLIT distance="200" swimtime="00:03:11.66" />
                    <SPLIT distance="250" swimtime="00:04:02.89" />
                    <SPLIT distance="300" swimtime="00:04:54.38" />
                    <SPLIT distance="350" swimtime="00:05:45.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="2615">
              <RESULTS>
                <RESULT eventid="1134" points="180" swimtime="00:00:42.52" resultid="2616" heatid="6992" lane="0" entrytime="00:00:40.26" />
                <RESULT eventid="1256" points="120" swimtime="00:00:45.40" resultid="2617" heatid="7037" lane="0" entrytime="00:00:44.96" />
                <RESULT eventid="1316" points="167" swimtime="00:01:34.29" resultid="2618" heatid="7069" lane="0" entrytime="00:01:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="172" swimtime="00:03:21.02" resultid="2619" heatid="7143" lane="1" entrytime="00:03:17.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="150" swimtime="00:02:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="167" swimtime="00:01:46.27" resultid="2620" heatid="7157" lane="0" entrytime="00:01:41.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-31" firstname="Zofia" gender="F" lastname="Kalinowska" nation="POL" athleteid="2621">
              <RESULTS>
                <RESULT eventid="1209" points="157" swimtime="00:03:45.72" resultid="2622" heatid="7023" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                    <SPLIT distance="100" swimtime="00:01:45.98" />
                    <SPLIT distance="150" swimtime="00:02:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="223" swimtime="00:01:32.31" resultid="2623" heatid="7105" lane="8" entrytime="00:01:31.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-09-16" firstname="Lina" gender="F" lastname="Varela-Machado" nation="POL" athleteid="2624">
              <RESULTS>
                <RESULT eventid="1058" points="224" swimtime="00:03:50.40" resultid="2625" heatid="6972" lane="9" entrytime="00:03:40.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.73" />
                    <SPLIT distance="100" swimtime="00:01:48.20" />
                    <SPLIT distance="150" swimtime="00:02:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="237" swimtime="00:01:24.07" resultid="2626" heatid="7005" lane="1" entrytime="00:01:23.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="175" swimtime="00:00:44.81" resultid="2627" heatid="7032" lane="6" entrytime="00:00:41.68" />
                <RESULT eventid="1361" points="209" swimtime="00:03:10.08" resultid="2628" heatid="7079" lane="2" entrytime="00:03:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:26.94" />
                    <SPLIT distance="150" swimtime="00:02:18.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="280" swimtime="00:00:36.27" resultid="2629" heatid="7118" lane="9" entrytime="00:00:35.59" />
                <RESULT eventid="1558" points="190" swimtime="00:06:55.54" resultid="2630" heatid="7165" lane="5" entrytime="00:06:43.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="150" swimtime="00:02:26.58" />
                    <SPLIT distance="200" swimtime="00:03:20.43" />
                    <SPLIT distance="250" swimtime="00:04:14.97" />
                    <SPLIT distance="300" swimtime="00:05:09.88" />
                    <SPLIT distance="350" swimtime="00:06:06.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-08" firstname="Paweł" gender="M" lastname="Salamończyk" nation="POL" athleteid="2631">
              <RESULTS>
                <RESULT eventid="1134" points="316" swimtime="00:00:35.29" resultid="2632" heatid="6994" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1194" points="401" swimtime="00:01:03.58" resultid="2633" heatid="7017" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="363" swimtime="00:00:31.43" resultid="2634" heatid="7042" lane="2" entrytime="00:00:30.92" />
                <RESULT eventid="1316" points="297" swimtime="00:01:17.81" resultid="2635" heatid="7070" lane="5" entrytime="00:01:14.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="402" swimtime="00:00:28.31" resultid="2636" heatid="7132" lane="8" entrytime="00:00:27.94" />
                <RESULT eventid="1498" points="279" swimtime="00:02:51.17" resultid="2637" heatid="7144" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:06.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Agnieszka" gender="F" lastname="Misiewicz" nation="POL" athleteid="7593" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1331" points="233" swimtime="00:02:37.13" resultid="7592" heatid="7073" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:02:01.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2621" number="1" />
                    <RELAYPOSITION athleteid="2624" number="2" />
                    <RELAYPOSITION athleteid="7593" number="3" />
                    <RELAYPOSITION athleteid="2602" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1513" points="190" swimtime="00:02:42.40" resultid="2638" heatid="7149" lane="9" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2631" number="1" />
                    <RELAYPOSITION athleteid="2608" number="2" />
                    <RELAYPOSITION athleteid="2621" number="3" />
                    <RELAYPOSITION athleteid="2624" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAOPO" name="Tp Masters Opole" nation="POL" region="OPO">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="TADEUSZ" gender="M" lastname="WITKOWSKI" nation="POL" athleteid="2653">
              <RESULTS>
                <RESULT eventid="1134" points="116" swimtime="00:00:49.26" resultid="2654" heatid="6988" lane="2" entrytime="00:00:55.50" />
                <RESULT eventid="1194" points="156" swimtime="00:01:27.07" resultid="2655" heatid="7011" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="143" swimtime="00:00:50.94" resultid="2656" heatid="7052" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1316" points="93" swimtime="00:01:54.57" resultid="2657" heatid="7067" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="204" swimtime="00:00:35.49" resultid="2658" heatid="7123" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1498" points="91" swimtime="00:04:08.33" resultid="2659" heatid="7141" lane="4" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.29" />
                    <SPLIT distance="100" swimtime="00:02:03.20" />
                    <SPLIT distance="150" swimtime="00:03:08.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="OLGIERD" gender="M" lastname="MIKOSZA" nation="POL" athleteid="2660">
              <RESULTS>
                <RESULT eventid="1134" points="235" swimtime="00:00:38.93" resultid="2661" heatid="6993" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1194" points="273" swimtime="00:01:12.27" resultid="2662" heatid="7015" lane="2" entrytime="00:01:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="222" swimtime="00:01:25.66" resultid="2663" heatid="7069" lane="2" entrytime="00:01:24.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="197" swimtime="00:02:55.20" resultid="2664" heatid="7085" lane="7" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                    <SPLIT distance="150" swimtime="00:02:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="321" swimtime="00:00:30.53" resultid="2665" heatid="7129" lane="6" entrytime="00:00:29.80" />
                <RESULT eventid="1498" points="178" swimtime="00:03:18.62" resultid="2666" heatid="7143" lane="7" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:36.89" />
                    <SPLIT distance="150" swimtime="00:02:30.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="JANUSZ" gender="M" lastname="SZPALA" nation="POL" athleteid="2667">
              <RESULTS>
                <RESULT eventid="1134" points="94" swimtime="00:00:52.81" resultid="2668" heatid="6990" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1256" points="99" swimtime="00:00:48.47" resultid="2669" heatid="7037" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1406" points="95" swimtime="00:04:09.33" resultid="2670" heatid="7096" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                    <SPLIT distance="100" swimtime="00:02:00.15" />
                    <SPLIT distance="150" swimtime="00:03:13.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="75" swimtime="00:01:58.03" resultid="2671" heatid="7107" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="JERZY" gender="M" lastname="MINKIEWICZ" nation="POL" athleteid="2672">
              <RESULTS>
                <RESULT eventid="1134" points="190" swimtime="00:00:41.81" resultid="2673" heatid="6991" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1194" points="290" swimtime="00:01:10.83" resultid="2674" heatid="7015" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="235" swimtime="00:00:36.34" resultid="2675" heatid="7040" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1316" points="172" swimtime="00:01:33.23" resultid="2676" heatid="7069" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="301" swimtime="00:00:31.18" resultid="2677" heatid="7127" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-01-01" firstname="JÓZEF" gender="M" lastname="KASPEREK" nation="POL" athleteid="2678">
              <RESULTS>
                <RESULT eventid="1316" points="21" swimtime="00:03:07.44" resultid="2679" heatid="7066" lane="7" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="19" swimtime="00:06:20.67" resultid="2680" heatid="7082" lane="6" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.17" />
                    <SPLIT distance="100" swimtime="00:02:59.16" />
                    <SPLIT distance="150" swimtime="00:04:44.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-01-01" firstname="BRONISŁAW" gender="M" lastname="PICHURSKI" nation="POL" athleteid="2681">
              <RESULTS>
                <RESULT eventid="1104" points="15" swimtime="00:08:33.95" resultid="2682" heatid="6974" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.84" />
                    <SPLIT distance="100" swimtime="00:03:59.42" />
                    <SPLIT distance="150" swimtime="00:06:21.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="16" swimtime="00:01:44.20" resultid="2683" heatid="7052" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1543" points="15" swimtime="00:03:56.89" resultid="2684" heatid="7155" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1164" points="159" swimtime="00:02:52.36" resultid="7176" heatid="6999" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:02:12.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2660" number="1" />
                    <RELAYPOSITION athleteid="2672" number="2" />
                    <RELAYPOSITION athleteid="2667" number="3" />
                    <RELAYPOSITION athleteid="2653" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="231" swimtime="00:02:18.25" resultid="7177" heatid="7074" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:40.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2653" number="1" />
                    <RELAYPOSITION athleteid="2672" number="2" />
                    <RELAYPOSITION athleteid="2667" number="3" />
                    <RELAYPOSITION athleteid="2660" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" name="MOSiR Ostrowiec Świętokrzyski" nation="POL" region="SWI">
          <CONTACT city="Ostrowiec Św." email="basen@mosir.ostrowiec.pl" name="Różalski" street="Józef" zip="27-400" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="M01012200001" athleteid="2686">
              <RESULTS>
                <RESULT eventid="1104" points="169" swimtime="00:03:50.07" resultid="2687" heatid="6975" lane="6" entrytime="00:03:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.57" />
                    <SPLIT distance="100" swimtime="00:01:50.35" />
                    <SPLIT distance="150" swimtime="00:02:50.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="235" swimtime="00:01:15.97" resultid="2688" heatid="7014" lane="9" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="241" swimtime="00:00:36.01" resultid="2689" heatid="7040" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1406" points="145" swimtime="00:03:36.50" resultid="2690" heatid="7096" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                    <SPLIT distance="100" swimtime="00:01:49.10" />
                    <SPLIT distance="150" swimtime="00:02:51.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="117" swimtime="00:01:41.58" resultid="2691" heatid="7107" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="258" swimtime="00:00:32.82" resultid="2692" heatid="7126" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOPIE" name="MOSiR Piekary Śląskie" nation="POL" region="SLA">
          <CONTACT email="bartolomeo863@wp.pl" name="Sz" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Bartosz" gender="M" lastname="Szymik" nation="POL" athleteid="2751">
              <RESULTS>
                <RESULT eventid="1104" points="321" swimtime="00:03:05.75" resultid="2752" heatid="6978" lane="7" entrytime="00:03:10.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                    <SPLIT distance="150" swimtime="00:02:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2753" heatid="7027" lane="5" entrytime="00:03:08.48" />
                <RESULT eventid="1286" points="395" swimtime="00:00:36.34" resultid="2754" heatid="7059" lane="2" entrytime="00:00:35.86" />
                <RESULT eventid="1406" points="293" swimtime="00:02:51.51" resultid="2755" heatid="7100" lane="1" entrytime="00:02:49.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:09.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2756" heatid="7144" lane="9" entrytime="00:03:02.67" />
                <RESULT eventid="1543" points="336" swimtime="00:01:24.21" resultid="2757" heatid="7160" lane="4" entrytime="00:01:23.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" name="KS Masters Polkowice" nation="POL" region="DOL">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-05-30" firstname="Grażyna" gender="F" lastname="Grzegorzewska" nation="POL" athleteid="2772">
              <RESULTS>
                <RESULT eventid="1119" points="106" swimtime="00:00:57.12" resultid="2773" heatid="6982" lane="5" entrytime="00:00:54.50" entrycourse="SCM" />
                <RESULT eventid="1179" points="165" swimtime="00:01:34.86" resultid="2774" heatid="7004" lane="9" entrytime="00:01:34.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="88" swimtime="00:00:56.28" resultid="2775" heatid="7031" lane="0" entrytime="00:00:52.30" entrycourse="SCM" />
                <RESULT eventid="1361" points="136" swimtime="00:03:39.48" resultid="2776" heatid="7078" lane="2" entrytime="00:03:33.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:44.72" />
                    <SPLIT distance="150" swimtime="00:02:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="193" swimtime="00:00:41.05" resultid="2777" heatid="7116" lane="0" entrytime="00:00:40.20" entrycourse="SCM" />
                <RESULT eventid="1558" points="138" swimtime="00:07:42.44" resultid="2778" heatid="7164" lane="5" entrytime="00:07:30.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:47.01" />
                    <SPLIT distance="150" swimtime="00:02:46.43" />
                    <SPLIT distance="200" swimtime="00:03:46.72" />
                    <SPLIT distance="250" swimtime="00:04:46.75" />
                    <SPLIT distance="300" swimtime="00:05:46.91" />
                    <SPLIT distance="350" swimtime="00:06:46.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="2779">
              <RESULTS>
                <RESULT eventid="1134" points="295" swimtime="00:00:36.11" resultid="2780" heatid="6994" lane="5" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1316" points="276" swimtime="00:01:19.72" resultid="2781" heatid="7070" lane="4" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="262" swimtime="00:02:54.87" resultid="2782" heatid="7145" lane="5" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                    <SPLIT distance="150" swimtime="00:02:08.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="2783">
              <RESULTS>
                <RESULT eventid="1104" points="96" swimtime="00:04:37.13" resultid="2784" heatid="6974" lane="2" entrytime="00:04:44.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.08" />
                    <SPLIT distance="100" swimtime="00:02:15.73" />
                    <SPLIT distance="150" swimtime="00:03:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="98" swimtime="00:01:41.63" resultid="2785" heatid="7010" lane="6" entrytime="00:01:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="119" swimtime="00:00:54.09" resultid="2786" heatid="7053" lane="7" entrytime="00:00:53.10" entrycourse="LCM" />
                <RESULT eventid="1406" points="75" swimtime="00:04:30.27" resultid="2787" heatid="7095" lane="5" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.63" />
                    <SPLIT distance="100" swimtime="00:02:16.15" />
                    <SPLIT distance="150" swimtime="00:03:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="57" swimtime="00:04:49.99" resultid="2788" heatid="7141" lane="7" entrytime="00:04:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.28" />
                    <SPLIT distance="100" swimtime="00:02:21.12" />
                    <SPLIT distance="150" swimtime="00:03:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="102" swimtime="00:02:05.03" resultid="2789" heatid="7156" lane="9" entrytime="00:02:06.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WAPOZ" name="Ks Warta Poznań" nation="POL" region="WIE">
          <CONTACT city="POZNAŃ" email="j.thiem@glos.com" name="THIEM JACEK" phone="502 499 565" state="WIE" street="OS. DĘBINA 19 M 34" zip="61450" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="JACEK" gender="M" lastname="THIEM" nation="POL" athleteid="2794">
              <RESULTS>
                <RESULT eventid="1224" points="193" swimtime="00:03:12.93" resultid="2795" heatid="7027" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:32.64" />
                    <SPLIT distance="150" swimtime="00:02:22.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="212" swimtime="00:00:37.58" resultid="2796" heatid="7038" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="2797" heatid="7085" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="1438" points="184" swimtime="00:01:27.58" resultid="2798" heatid="7108" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="138" swimtime="00:03:36.25" resultid="2799" heatid="7142" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.48" />
                    <SPLIT distance="100" swimtime="00:01:50.94" />
                    <SPLIT distance="150" swimtime="00:02:45.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="ANNA" gender="F" lastname="KOTECKA" nation="POL" athleteid="2801">
              <RESULTS>
                <RESULT eventid="1119" points="190" swimtime="00:00:47.02" resultid="2802" heatid="6983" lane="4" entrytime="00:00:46.90" />
                <RESULT eventid="1179" points="261" swimtime="00:01:21.42" resultid="2803" heatid="7005" lane="2" entrytime="00:01:22.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="213" swimtime="00:01:37.23" resultid="2804" heatid="7064" lane="0" entrytime="00:01:38.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" status="DNS" swimtime="00:00:00.00" resultid="2805" heatid="7079" lane="6" entrytime="00:03:04.50" />
                <RESULT eventid="1483" status="DNS" swimtime="00:00:00.00" resultid="2806" heatid="7138" lane="7" entrytime="00:03:28.10" />
                <RESULT eventid="1558" points="244" swimtime="00:06:22.42" resultid="2807" heatid="7164" lane="3" entrytime="00:06:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                    <SPLIT distance="150" swimtime="00:02:18.46" />
                    <SPLIT distance="200" swimtime="00:03:07.18" />
                    <SPLIT distance="250" swimtime="00:03:56.61" />
                    <SPLIT distance="300" swimtime="00:04:45.63" />
                    <SPLIT distance="350" swimtime="00:05:35.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="PAWEŁ" gender="M" lastname="OLSZEWSKI" nation="POL" athleteid="2808">
              <RESULTS>
                <RESULT eventid="1194" points="451" swimtime="00:01:01.14" resultid="2809" heatid="7019" lane="4" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="384" swimtime="00:02:20.33" resultid="2810" heatid="7089" lane="9" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="415" swimtime="00:00:28.02" resultid="2811" heatid="7130" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1573" points="369" swimtime="00:05:06.58" resultid="2812" heatid="7173" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:45.74" />
                    <SPLIT distance="200" swimtime="00:02:23.57" />
                    <SPLIT distance="250" swimtime="00:03:02.82" />
                    <SPLIT distance="300" swimtime="00:03:42.87" />
                    <SPLIT distance="350" swimtime="00:04:25.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-07-08" firstname="TOMASZ" gender="M" lastname="RYBAK" nation="POL" athleteid="2813">
              <RESULTS>
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="2814" heatid="6994" lane="8" entrytime="00:00:35.50" />
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="2815" heatid="7016" lane="7" entrytime="00:01:08.00" />
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="2816" heatid="7070" lane="7" entrytime="00:01:17.90" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="2817" heatid="7098" lane="5" entrytime="00:02:57.90" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="2818" heatid="7144" lane="2" entrytime="00:02:56.30" />
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="2819" heatid="7170" lane="1" entrytime="00:05:45.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="DARIUSZ" gender="M" lastname="JANYGA" nation="POL" athleteid="2820">
              <RESULTS>
                <RESULT eventid="1134" points="309" swimtime="00:00:35.54" resultid="2821" heatid="6994" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1194" points="346" swimtime="00:01:06.80" resultid="2822" heatid="7016" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="278" swimtime="00:01:19.49" resultid="2823" heatid="7069" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="346" swimtime="00:00:29.77" resultid="2824" heatid="7128" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="1498" points="231" swimtime="00:03:02.39" resultid="2825" heatid="7142" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:13.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-30" firstname="ALEKSANDRA" gender="F" lastname="GÓRNIAK" nation="POL" athleteid="2826">
              <RESULTS>
                <RESULT eventid="1119" points="361" swimtime="00:00:38.00" resultid="2827" heatid="6986" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1301" points="334" swimtime="00:01:23.69" resultid="2828" heatid="7065" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="330" swimtime="00:03:00.55" resultid="2829" heatid="7139" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="150" swimtime="00:02:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="PRZEMYSŁAW" gender="M" lastname="WARACZEWSKI" nation="POL" athleteid="2830">
              <RESULTS>
                <RESULT eventid="1104" points="283" swimtime="00:03:13.70" resultid="2831" heatid="6977" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:31.90" />
                    <SPLIT distance="150" swimtime="00:02:22.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="241" swimtime="00:00:38.58" resultid="2832" heatid="6990" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1286" points="326" swimtime="00:00:38.74" resultid="2833" heatid="7054" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1316" points="211" swimtime="00:01:27.18" resultid="2834" heatid="7068" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="288" swimtime="00:01:28.63" resultid="2835" heatid="7158" lane="1" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="2837" heatid="7000" lane="3" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2820" number="1" />
                    <RELAYPOSITION athleteid="2808" number="2" />
                    <RELAYPOSITION athleteid="2813" number="3" />
                    <RELAYPOSITION athleteid="2830" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="2836" heatid="7075" lane="6" entrytime="00:01:59.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2808" number="1" />
                    <RELAYPOSITION athleteid="2830" number="2" />
                    <RELAYPOSITION athleteid="2813" number="3" />
                    <RELAYPOSITION athleteid="2820" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1513" points="201" swimtime="00:02:39.46" resultid="2838" heatid="7148" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                    <SPLIT distance="150" swimtime="00:02:05.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2801" number="1" />
                    <RELAYPOSITION athleteid="2830" number="2" />
                    <RELAYPOSITION athleteid="2794" number="3" />
                    <RELAYPOSITION athleteid="2826" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MKSZC" name="MKP Szczecin" nation="POL" region="ZAC">
          <CONTACT city="Szczecin" email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" state="ZACHO" street="Kaliny 45/9" zip="71-118" />
          <ATHLETES>
            <ATHLETE birthdate="1942-07-12" firstname="Jerzy" gender="M" lastname="Rabiej" nation="POL" license="S001166200549" athleteid="2846">
              <RESULTS>
                <RESULT eventid="1134" points="106" swimtime="00:00:50.78" resultid="2847" heatid="6992" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1316" points="72" swimtime="00:02:04.72" resultid="2848" heatid="7068" lane="0" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="61" swimtime="00:04:43.53" resultid="2849" heatid="7142" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.21" />
                    <SPLIT distance="100" swimtime="00:02:19.38" />
                    <SPLIT distance="150" swimtime="00:03:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="78" swimtime="00:08:34.48" resultid="2850" heatid="7168" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.14" />
                    <SPLIT distance="100" swimtime="00:02:05.47" />
                    <SPLIT distance="150" swimtime="00:03:13.48" />
                    <SPLIT distance="200" swimtime="00:04:19.63" />
                    <SPLIT distance="250" swimtime="00:05:26.46" />
                    <SPLIT distance="300" swimtime="00:06:32.68" />
                    <SPLIT distance="350" swimtime="00:07:37.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="2863">
              <RESULTS>
                <RESULT eventid="1194" points="463" swimtime="00:01:00.61" resultid="2864" heatid="7019" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="396" swimtime="00:02:18.89" resultid="2865" heatid="7088" lane="3" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="384" swimtime="00:05:02.65" resultid="2866" heatid="7173" lane="9" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                    <SPLIT distance="200" swimtime="00:02:29.19" />
                    <SPLIT distance="250" swimtime="00:03:08.03" />
                    <SPLIT distance="300" swimtime="00:03:47.88" />
                    <SPLIT distance="350" swimtime="00:04:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-08" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="2867">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. E /45-49/" eventid="1179" points="444" swimtime="00:01:08.25" resultid="2868" heatid="7008" lane="8" entrytime="00:01:08.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. E /45-49/" eventid="1361" points="486" swimtime="00:02:23.65" resultid="2869" heatid="7081" lane="3" entrytime="00:02:22.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="451" swimtime="00:05:11.76" resultid="2870" heatid="7167" lane="4" entrytime="00:04:59.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:53.59" />
                    <SPLIT distance="200" swimtime="00:02:33.28" />
                    <SPLIT distance="250" swimtime="00:03:13.15" />
                    <SPLIT distance="300" swimtime="00:03:53.19" />
                    <SPLIT distance="350" swimtime="00:04:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="2871">
              <RESULTS>
                <RESULT eventid="1134" points="154" swimtime="00:00:44.82" resultid="2872" heatid="6990" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1194" status="DNF" swimtime="00:00:00.00" resultid="2873" heatid="7011" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1376" points="175" swimtime="00:03:02.34" resultid="2874" heatid="7083" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:27.46" />
                    <SPLIT distance="150" swimtime="00:02:15.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="195" swimtime="00:00:36.00" resultid="2875" heatid="7123" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOSIE" name="Wodnik Siemianowice Śląskie" nation="POL" region="SLA">
          <CONTACT email="bartolomeo863@wp.pl" name="Szymik Bartosz" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="2852">
              <RESULTS>
                <RESULT eventid="1104" points="208" swimtime="00:03:34.75" resultid="2853" heatid="6977" lane="9" entrytime="00:03:20.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.65" />
                    <SPLIT distance="100" swimtime="00:01:43.52" />
                    <SPLIT distance="150" swimtime="00:02:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="186" swimtime="00:03:15.15" resultid="2854" heatid="7027" lane="1" entrytime="00:03:16.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="241" swimtime="00:00:36.04" resultid="2855" heatid="7039" lane="6" entrytime="00:00:35.35" />
                <RESULT eventid="1406" points="268" swimtime="00:02:56.68" resultid="2856" heatid="7098" lane="3" entrytime="00:02:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:25.20" />
                    <SPLIT distance="150" swimtime="00:02:17.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="209" swimtime="00:01:23.88" resultid="2857" heatid="7109" lane="9" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="277" swimtime="00:05:37.55" resultid="2858" heatid="7171" lane="8" entrytime="00:05:32.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:05.07" />
                    <SPLIT distance="200" swimtime="00:02:48.10" />
                    <SPLIT distance="250" swimtime="00:03:31.27" />
                    <SPLIT distance="300" swimtime="00:04:14.05" />
                    <SPLIT distance="350" swimtime="00:04:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TAKAS" name="Takas" nation="LTU">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Romaldas Bickauskas" phone="+37068687934" street="Lentvario g. 19-1" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas" gender="M" lastname="JUODESKA" nation="LTU" athleteid="2877">
              <RESULTS>
                <RESULT comment="K-3 - Brak wynurzenia głowy w drugim cyklu po nawrocie" eventid="1104" status="DSQ" swimtime="00:03:12.07" resultid="2878" heatid="6977" lane="5" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:32.31" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="363" swimtime="00:00:37.36" resultid="2879" heatid="7058" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1406" points="272" swimtime="00:02:55.82" resultid="2880" heatid="7099" lane="7" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="340" swimtime="00:00:29.94" resultid="2881" heatid="7130" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1543" points="318" swimtime="00:01:25.81" resultid="2882" heatid="7160" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-08" firstname="Pavelas" gender="M" lastname="bezzubovas" nation="LTU" athleteid="2883">
              <RESULTS>
                <RESULT eventid="1256" points="140" swimtime="00:00:43.12" resultid="2884" heatid="7038" lane="8" entrytime="00:00:38.50" />
                <RESULT eventid="1286" points="145" swimtime="00:00:50.76" resultid="2885" heatid="7055" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1468" points="190" swimtime="00:00:36.36" resultid="2886" heatid="7124" lane="6" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-25" firstname="Arturas" gender="M" lastname="tuomas" nation="LTU" athleteid="2887">
              <RESULTS>
                <RESULT eventid="1224" points="221" swimtime="00:03:04.32" resultid="2888" heatid="7028" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:35.21" />
                    <SPLIT distance="150" swimtime="00:02:25.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="286" swimtime="00:02:52.85" resultid="2889" heatid="7100" lane="3" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:12.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="268" swimtime="00:01:17.21" resultid="2890" heatid="7111" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-22" firstname="Arvydas" gender="M" lastname="burinskas" nation="LTU" athleteid="2891">
              <RESULTS>
                <RESULT eventid="1224" points="260" swimtime="00:02:54.52" resultid="2892" heatid="7028" lane="6" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="366" swimtime="00:00:31.35" resultid="2893" heatid="7043" lane="0" entrytime="00:00:30.50" />
                <RESULT eventid="1438" points="321" swimtime="00:01:12.75" resultid="2894" heatid="7111" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1927-04-21" firstname="Vladas" gender="M" lastname="vimbaras" nation="LTU" athleteid="2895">
              <RESULTS>
                <RESULT eventid="1134" points="39" swimtime="00:01:10.46" resultid="2896" heatid="6988" lane="9" entrytime="00:01:05.00" />
                <RESULT eventid="1194" points="34" swimtime="00:02:24.77" resultid="2897" heatid="7009" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="22" swimtime="00:03:04.28" resultid="2898" heatid="7066" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="72" swimtime="00:00:50.12" resultid="2899" heatid="7122" lane="8" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-09-25" firstname="Vytautas" gender="M" lastname="svetikas" nation="LTU" athleteid="2900">
              <RESULTS>
                <RESULT eventid="1194" points="126" swimtime="00:01:33.54" resultid="2901" heatid="7011" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="2902" heatid="7085" lane="8" entrytime="00:02:50.00" />
                <RESULT eventid="1468" points="158" swimtime="00:00:38.62" resultid="2903" heatid="7124" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-14" firstname="Romaldas" gender="M" lastname="bickauskas" nation="LTU" athleteid="2904">
              <RESULTS>
                <RESULT eventid="1256" points="155" swimtime="00:00:41.73" resultid="2905" heatid="7039" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="1438" points="85" swimtime="00:01:52.98" resultid="6417" heatid="7107" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-25" firstname="Dalicija" gender="F" lastname="fedoraviciene" nation="LTU" athleteid="2907">
              <RESULTS>
                <RESULT eventid="1179" points="70" swimtime="00:02:06.03" resultid="2908" heatid="7003" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="67" swimtime="00:04:36.82" resultid="2909" heatid="7077" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.15" />
                    <SPLIT distance="100" swimtime="00:02:18.67" />
                    <SPLIT distance="150" swimtime="00:03:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="92" swimtime="00:00:52.43" resultid="2910" heatid="7115" lane="9" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-02" firstname="Elena" gender="F" lastname="baumanaite" nation="LTU" athleteid="2911">
              <RESULTS>
                <RESULT eventid="1119" points="16" swimtime="00:01:46.33" resultid="2912" heatid="6982" lane="8" entrytime="00:01:15.00" />
                <RESULT eventid="1453" points="26" swimtime="00:01:19.82" resultid="2913" heatid="7114" lane="1" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="ivanauskaite" nation="LTU" athleteid="2914">
              <RESULTS>
                <RESULT eventid="1119" points="277" swimtime="00:00:41.51" resultid="2915" heatid="6985" lane="0" entrytime="00:00:40.70" />
                <RESULT eventid="1301" points="300" swimtime="00:01:26.74" resultid="2916" heatid="7064" lane="6" entrytime="00:01:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="306" swimtime="00:02:47.63" resultid="2917" heatid="7080" lane="1" entrytime="00:02:50.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:01:20.53" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="306" swimtime="00:03:05.17" resultid="2918" heatid="7139" lane="7" entrytime="00:03:07.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="308" swimtime="00:05:54.11" resultid="2919" heatid="7166" lane="5" entrytime="00:05:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:22.21" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                    <SPLIT distance="200" swimtime="00:02:51.33" />
                    <SPLIT distance="250" swimtime="00:03:37.21" />
                    <SPLIT distance="300" swimtime="00:04:23.98" />
                    <SPLIT distance="350" swimtime="00:05:10.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="kersevicius" nation="LTU" athleteid="2920">
              <RESULTS>
                <RESULT eventid="1134" points="401" swimtime="00:00:32.59" resultid="2921" heatid="6996" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1316" points="406" swimtime="00:01:10.14" resultid="2922" heatid="7071" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="386" swimtime="00:02:33.61" resultid="2923" heatid="7146" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:54.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-15" firstname="Daiva" gender="F" lastname="Diedoniene" nation="LTU" athleteid="2924">
              <RESULTS>
                <RESULT eventid="1240" points="278" swimtime="00:00:38.39" resultid="2925" heatid="7033" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1453" points="276" swimtime="00:00:36.41" resultid="2926" heatid="7118" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-26" firstname="Ausra" gender="F" lastname="patasiene" nation="LTU" athleteid="2927">
              <RESULTS>
                <RESULT eventid="1240" points="175" swimtime="00:00:44.78" resultid="2928" heatid="7032" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1453" points="237" swimtime="00:00:38.33" resultid="2929" heatid="7116" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-08-11" firstname="Audrius" gender="M" lastname="kiauke" nation="LTU" athleteid="2930">
              <RESULTS>
                <RESULT eventid="1194" points="255" swimtime="00:01:13.94" resultid="2931" heatid="7014" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="217" swimtime="00:02:49.73" resultid="2932" heatid="7086" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="252" swimtime="00:00:33.10" resultid="2933" heatid="7126" lane="7" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="yliene" nation="LTU" athleteid="2934">
              <RESULTS>
                <RESULT eventid="1119" points="157" swimtime="00:00:50.14" resultid="2935" heatid="6983" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1301" points="118" swimtime="00:01:58.22" resultid="2936" heatid="7063" lane="3" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="102" swimtime="00:04:27.04" resultid="2937" heatid="7137" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.56" />
                    <SPLIT distance="100" swimtime="00:02:12.49" />
                    <SPLIT distance="150" swimtime="00:03:23.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-19" firstname="Pavel" gender="M" lastname="Protasciuk" nation="LTU" athleteid="2938">
              <RESULTS>
                <RESULT eventid="1134" points="411" swimtime="00:00:32.33" resultid="2939" heatid="6996" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1256" points="496" swimtime="00:00:28.33" resultid="2940" heatid="7044" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1406" points="457" swimtime="00:02:27.91" resultid="2941" heatid="7103" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="479" swimtime="00:00:26.72" resultid="2942" heatid="7134" lane="4" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-28" firstname="Giedrius" gender="M" lastname="Zalionis" nation="LTU" athleteid="2943">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="2944" heatid="7044" lane="7" entrytime="00:00:28.90" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="2945" heatid="7134" lane="6" entrytime="00:00:26.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-04-10" firstname="Loreta" gender="F" lastname="kabasinskiene" nation="LTU" athleteid="2946">
              <RESULTS>
                <RESULT eventid="1179" points="210" swimtime="00:01:27.55" resultid="2947" heatid="7004" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="209" swimtime="00:03:32.52" resultid="2948" heatid="7093" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                    <SPLIT distance="100" swimtime="00:01:45.49" />
                    <SPLIT distance="150" swimtime="00:02:45.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="159" swimtime="00:01:43.28" resultid="2949" heatid="7104" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-08" firstname="Viktoras" gender="M" lastname="SNIESKA" nation="LTU" athleteid="2950">
              <RESULTS>
                <RESULT eventid="1134" points="213" swimtime="00:00:40.23" resultid="2951" heatid="6990" lane="5" entrytime="00:00:42.10" />
                <RESULT eventid="1194" points="267" swimtime="00:01:12.76" resultid="2952" heatid="7013" lane="5" entrytime="00:01:14.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="175" swimtime="00:01:32.72" resultid="2953" heatid="7068" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="187" swimtime="00:02:58.25" resultid="2954" heatid="7084" lane="5" entrytime="00:02:52.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:02:14.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="255" swimtime="00:00:32.97" resultid="2955" heatid="7125" lane="1" entrytime="00:00:33.58" />
                <RESULT eventid="1498" points="161" swimtime="00:03:25.68" resultid="2956" heatid="7142" lane="4" entrytime="00:03:25.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:32.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-01" firstname="Nerimantas" gender="M" lastname="steponavicius" nation="LTU" athleteid="2957">
              <RESULTS>
                <RESULT eventid="1286" points="433" swimtime="00:00:35.23" resultid="2958" heatid="7060" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1164" points="106" swimtime="00:03:16.99" resultid="7223" heatid="6999" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.05" />
                    <SPLIT distance="100" swimtime="00:01:40.00" />
                    <SPLIT distance="150" swimtime="00:02:24.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2904" number="1" />
                    <RELAYPOSITION athleteid="2950" number="2" />
                    <RELAYPOSITION athleteid="2900" number="3" />
                    <RELAYPOSITION athleteid="2895" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="136" swimtime="00:02:44.87" resultid="7606" heatid="7074" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                    <SPLIT distance="150" swimtime="00:02:09.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2895" number="1" />
                    <RELAYPOSITION athleteid="2883" number="2" />
                    <RELAYPOSITION athleteid="2900" number="3" />
                    <RELAYPOSITION athleteid="2950" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1164" points="361" swimtime="00:02:11.15" resultid="7224" heatid="6999" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:44.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2877" number="1" />
                    <RELAYPOSITION athleteid="2920" number="2" />
                    <RELAYPOSITION athleteid="2938" number="3" />
                    <RELAYPOSITION athleteid="2887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1331" points="176" swimtime="00:02:52.41" resultid="7605" heatid="7073" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.37" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:01:32.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2907" number="1" />
                    <RELAYPOSITION athleteid="2914" number="2" />
                    <RELAYPOSITION athleteid="2946" number="3" />
                    <RELAYPOSITION athleteid="2934" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1513" status="DSQ" swimtime="00:03:08.36" resultid="7616" heatid="7148" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:32.88" />
                    <SPLIT distance="150" swimtime="00:01:23.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2950" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2883" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2946" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2907" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1513" points="246" swimtime="00:02:28.92" resultid="7617" heatid="7148" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:13.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2877" number="1" />
                    <RELAYPOSITION athleteid="2891" number="2" />
                    <RELAYPOSITION athleteid="2924" number="3" />
                    <RELAYPOSITION athleteid="2927" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1513" points="184" swimtime="00:02:44.26" resultid="7621" heatid="7148" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                    <SPLIT distance="100" swimtime="00:01:37.06" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2934" number="1" />
                    <RELAYPOSITION athleteid="2914" number="2" />
                    <RELAYPOSITION athleteid="2887" number="3" />
                    <RELAYPOSITION athleteid="2930" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WMT" name="Warsaw Masters Team" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="jstobnic@gmail.com" internet="masters.waw.pl" name="Justyna Marta Stobnicka" state="MAZ" />
          <ATHLETES>
            <ATHLETE birthdate="1978-02-01" firstname="Dariusz" gender="M" lastname="Dębski" nation="POL" athleteid="2972">
              <RESULTS>
                <RESULT eventid="1194" points="369" swimtime="00:01:05.36" resultid="2973" heatid="7017" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="282" swimtime="00:00:34.17" resultid="2974" heatid="7040" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1468" points="378" swimtime="00:00:28.91" resultid="2975" heatid="7130" lane="8" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-01" firstname="Paweł" gender="M" lastname="Kowalewski" nation="POL" athleteid="2976">
              <RESULTS>
                <RESULT eventid="1406" points="371" swimtime="00:02:38.52" resultid="2977" heatid="7102" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:02:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="308" swimtime="00:01:13.74" resultid="2978" heatid="7110" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="407" swimtime="00:04:56.76" resultid="2979" heatid="7173" lane="1" entrytime="00:04:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                    <SPLIT distance="200" swimtime="00:02:28.37" />
                    <SPLIT distance="250" swimtime="00:03:06.09" />
                    <SPLIT distance="300" swimtime="00:03:43.47" />
                    <SPLIT distance="350" swimtime="00:04:20.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="2980">
              <RESULTS>
                <RESULT eventid="1104" points="98" swimtime="00:04:35.21" resultid="2981" heatid="6974" lane="3" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.42" />
                    <SPLIT distance="100" swimtime="00:02:15.44" />
                    <SPLIT distance="150" swimtime="00:03:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. K /75-79/" eventid="1224" points="41" swimtime="00:05:23.13" resultid="2982" heatid="7025" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.13" />
                    <SPLIT distance="100" swimtime="00:02:37.19" />
                    <SPLIT distance="150" swimtime="00:04:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="61" swimtime="00:02:11.39" resultid="2983" heatid="7066" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="77" swimtime="00:04:27.59" resultid="2984" heatid="7095" lane="3" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                    <SPLIT distance="100" swimtime="00:02:11.22" />
                    <SPLIT distance="150" swimtime="00:03:22.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="69" swimtime="00:04:32.40" resultid="2985" heatid="7141" lane="8" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.53" />
                    <SPLIT distance="100" swimtime="00:02:14.81" />
                    <SPLIT distance="150" swimtime="00:03:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="106" swimtime="00:02:03.77" resultid="2986" heatid="7155" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-10" firstname="Maciej" gender="M" lastname="Burny" nation="POL" athleteid="2987">
              <RESULTS>
                <RESULT eventid="1468" points="491" swimtime="00:00:26.49" resultid="2988" heatid="7133" lane="4" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-06-24" firstname="Krzysztof" gender="M" lastname="Tomaszewski" nation="POL" athleteid="2989">
              <RESULTS>
                <RESULT eventid="1134" points="98" swimtime="00:00:52.01" resultid="2990" heatid="6989" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1286" points="113" swimtime="00:00:55.05" resultid="2991" heatid="7053" lane="2" entrytime="00:00:53.00" />
                <RESULT eventid="1468" points="119" swimtime="00:00:42.46" resultid="2992" heatid="7122" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1543" points="76" swimtime="00:02:17.85" resultid="2993" heatid="7155" lane="4" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-15" firstname="Jerzy" gender="M" lastname="Leszczyński" nation="POL" athleteid="2994">
              <RESULTS>
                <RESULT eventid="1104" points="318" swimtime="00:03:06.44" resultid="2995" heatid="6979" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                    <SPLIT distance="150" swimtime="00:02:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="330" swimtime="00:01:07.85" resultid="2996" heatid="7016" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="349" swimtime="00:00:37.87" resultid="2997" heatid="7057" lane="3" entrytime="00:00:37.70" />
                <RESULT eventid="1406" points="269" swimtime="00:02:56.52" resultid="2998" heatid="7099" lane="2" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:26.83" />
                    <SPLIT distance="150" swimtime="00:02:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="339" swimtime="00:00:29.97" resultid="2999" heatid="7130" lane="3" entrytime="00:00:28.70" />
                <RESULT eventid="1543" points="326" swimtime="00:01:25.05" resultid="3000" heatid="7161" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-01" firstname="Andrzej" gender="M" lastname="Ciesliński" nation="POL" athleteid="3001">
              <RESULTS>
                <RESULT eventid="1104" points="212" swimtime="00:03:33.27" resultid="3002" heatid="6976" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:41.91" />
                    <SPLIT distance="150" swimtime="00:02:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="195" swimtime="00:00:38.65" resultid="3003" heatid="7038" lane="5" entrytime="00:00:37.70" />
                <RESULT eventid="1468" points="248" swimtime="00:00:33.25" resultid="3004" heatid="7125" lane="6" entrytime="00:00:33.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-11-05" firstname="Mirosława" gender="F" lastname="Przyłuska" nation="POL" athleteid="3005">
              <RESULTS>
                <RESULT eventid="1271" points="149" swimtime="00:00:56.09" resultid="3006" heatid="7048" lane="5" entrytime="00:00:56.00" />
                <RESULT eventid="1361" points="67" swimtime="00:04:37.62" resultid="3007" heatid="7077" lane="5" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.35" />
                    <SPLIT distance="100" swimtime="00:02:15.77" />
                    <SPLIT distance="150" swimtime="00:03:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="129" swimtime="00:02:07.41" resultid="3008" heatid="7151" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="124" swimtime="00:04:40.50" resultid="5682" heatid="6971" lane="8" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.21" />
                    <SPLIT distance="100" swimtime="00:02:14.14" />
                    <SPLIT distance="150" swimtime="00:03:27.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="Dobczyńska" nation="POL" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1179" points="208" swimtime="00:01:27.75" resultid="3010" heatid="7004" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="222" swimtime="00:01:35.89" resultid="3011" heatid="7063" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="208" swimtime="00:03:10.45" resultid="3012" heatid="7079" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:30.92" />
                    <SPLIT distance="150" swimtime="00:02:21.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="211" swimtime="00:03:29.36" resultid="3013" heatid="7138" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.06" />
                    <SPLIT distance="100" swimtime="00:01:43.03" />
                    <SPLIT distance="150" swimtime="00:02:38.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-18" firstname="Robert" gender="M" lastname="Nowicki" nation="POL" athleteid="3014">
              <RESULTS>
                <RESULT eventid="1194" points="120" swimtime="00:01:35.06" resultid="3015" heatid="7010" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="123" swimtime="00:03:24.81" resultid="3016" heatid="7083" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="128" swimtime="00:00:41.42" resultid="3017" heatid="7122" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1573" points="137" swimtime="00:07:06.48" resultid="3018" heatid="7168" lane="4" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:33.17" />
                    <SPLIT distance="200" swimtime="00:03:29.00" />
                    <SPLIT distance="250" swimtime="00:04:24.44" />
                    <SPLIT distance="300" swimtime="00:05:19.98" />
                    <SPLIT distance="350" swimtime="00:06:16.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="3019">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. C /35-39/" eventid="1134" points="616" swimtime="00:00:28.25" resultid="3020" heatid="6997" lane="5" entrytime="00:00:27.99" />
                <RESULT comment="Rekord Polski Masters w kat. C /35-39/" eventid="1256" points="607" swimtime="00:00:26.49" resultid="3021" heatid="7046" lane="2" entrytime="00:00:26.26" />
                <RESULT comment="Rekord Polski Masters w kat. C /35-39/" eventid="1316" points="598" swimtime="00:01:01.64" resultid="3022" heatid="7072" lane="3" entrytime="00:01:02.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat C /35-39/" eventid="1438" points="569" swimtime="00:01:00.11" resultid="3023" heatid="7112" lane="2" entrytime="00:01:00.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-02" firstname="Andrzej" gender="M" lastname="Wiszniewski" nation="POL" athleteid="3024">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="3025" heatid="6976" lane="5" entrytime="00:03:27.20" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3026" heatid="7026" lane="8" entrytime="00:03:49.11" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3027" heatid="7036" lane="5" entrytime="00:00:48.10" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3028" heatid="7054" lane="9" entrytime="00:00:46.80" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="3029" heatid="7107" lane="0" entrytime="00:01:51.10" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="3030" heatid="7157" lane="2" entrytime="00:01:38.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-12-31" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="3031">
              <RESULTS>
                <RESULT eventid="1134" points="265" swimtime="00:00:37.40" resultid="3032" heatid="6993" lane="6" entrytime="00:00:36.55" />
                <RESULT eventid="1194" points="393" swimtime="00:01:04.02" resultid="3033" heatid="7017" lane="2" entrytime="00:01:05.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="304" swimtime="00:01:17.18" resultid="3034" heatid="7070" lane="2" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="327" swimtime="00:02:45.43" resultid="3035" heatid="7101" lane="3" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:09.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="295" swimtime="00:02:47.97" resultid="3036" heatid="7145" lane="7" entrytime="00:02:43.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:05.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-11-09" firstname="Tadeusz" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="3037">
              <RESULTS>
                <RESULT eventid="1468" points="150" swimtime="00:00:39.35" resultid="3038" heatid="7123" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Arkadiusz" gender="M" lastname="Dobrzyński" nation="POL" athleteid="3039">
              <RESULTS>
                <RESULT eventid="1134" points="396" swimtime="00:00:32.73" resultid="3040" heatid="6996" lane="8" entrytime="00:00:31.80" />
                <RESULT eventid="1316" points="355" swimtime="00:01:13.33" resultid="3041" heatid="7071" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="404" swimtime="00:00:28.27" resultid="3042" heatid="7134" lane="5" entrytime="00:00:26.70" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3043" heatid="7144" lane="5" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="3044">
              <RESULTS>
                <RESULT eventid="1134" points="391" swimtime="00:00:32.87" resultid="3045" heatid="6996" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1316" points="399" swimtime="00:01:10.51" resultid="3046" heatid="7071" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="406" swimtime="00:02:17.72" resultid="3047" heatid="7089" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:08.05" />
                    <SPLIT distance="150" swimtime="00:01:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3048" heatid="7146" lane="9" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="3049">
              <RESULTS>
                <RESULT eventid="1104" points="199" swimtime="00:03:37.93" resultid="3050" heatid="6976" lane="1" entrytime="00:03:35.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.32" />
                    <SPLIT distance="100" swimtime="00:01:42.25" />
                    <SPLIT distance="150" swimtime="00:02:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="87" swimtime="00:00:54.22" resultid="3051" heatid="6988" lane="5" entrytime="00:00:53.74" />
                <RESULT eventid="1194" points="146" swimtime="00:01:29.01" resultid="3052" heatid="7010" lane="5" entrytime="00:01:32.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="176" swimtime="00:00:47.51" resultid="3053" heatid="7054" lane="4" entrytime="00:00:44.26" />
                <RESULT eventid="1468" points="159" swimtime="00:00:38.52" resultid="3054" heatid="7122" lane="3" entrytime="00:00:40.46" />
                <RESULT eventid="1543" points="179" swimtime="00:01:43.77" resultid="3055" heatid="7157" lane="1" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="3056">
              <RESULTS>
                <RESULT eventid="1134" points="135" swimtime="00:00:46.86" resultid="3057" heatid="6989" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1194" points="183" swimtime="00:01:22.61" resultid="3058" heatid="7012" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="106" swimtime="00:01:49.53" resultid="3059" heatid="7067" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="131" swimtime="00:03:20.68" resultid="3060" heatid="7083" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:36.01" />
                    <SPLIT distance="150" swimtime="00:02:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="181" swimtime="00:00:36.92" resultid="3061" heatid="7123" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1573" points="125" swimtime="00:07:20.06" resultid="3062" heatid="7168" lane="5" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="100" swimtime="00:01:38.62" />
                    <SPLIT distance="150" swimtime="00:02:34.79" />
                    <SPLIT distance="200" swimtime="00:03:31.57" />
                    <SPLIT distance="250" swimtime="00:04:30.05" />
                    <SPLIT distance="300" swimtime="00:05:28.29" />
                    <SPLIT distance="350" swimtime="00:06:26.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="3063">
              <RESULTS>
                <RESULT eventid="1134" points="353" swimtime="00:00:33.99" resultid="3064" heatid="6995" lane="9" entrytime="00:00:34.11" />
                <RESULT comment="Rekord Polski Masters w kat. F /50-54/" eventid="1194" points="515" swimtime="00:00:58.52" resultid="3065" heatid="7020" lane="4" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="428" swimtime="00:00:29.75" resultid="3066" heatid="7043" lane="7" entrytime="00:00:30.09" />
                <RESULT comment="Rekord Polski Masters w kat. F /50-54/" eventid="1376" points="438" swimtime="00:02:14.31" resultid="3067" heatid="7089" lane="0" entrytime="00:02:16.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="445" swimtime="00:00:27.37" resultid="3068" heatid="7133" lane="2" entrytime="00:00:27.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-19" firstname="Dominik" gender="M" lastname="Bekierski" nation="POL" athleteid="3069">
              <RESULTS>
                <RESULT eventid="1134" points="506" swimtime="00:00:30.15" resultid="3070" heatid="6997" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1194" points="487" swimtime="00:00:59.61" resultid="3071" heatid="7021" lane="6" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="492" swimtime="00:01:05.79" resultid="3072" heatid="7072" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="418" swimtime="00:02:32.41" resultid="3073" heatid="7103" lane="2" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="440" swimtime="00:02:27.12" resultid="3074" heatid="7146" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="150" swimtime="00:01:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="421" swimtime="00:04:53.49" resultid="3075" heatid="7174" lane="0" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                    <SPLIT distance="150" swimtime="00:01:40.59" />
                    <SPLIT distance="200" swimtime="00:02:18.17" />
                    <SPLIT distance="250" swimtime="00:02:56.85" />
                    <SPLIT distance="300" swimtime="00:03:36.14" />
                    <SPLIT distance="350" swimtime="00:04:15.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="3076">
              <RESULTS>
                <RESULT eventid="1104" points="495" swimtime="00:02:40.93" resultid="3077" heatid="6980" lane="8" entrytime="00:02:48.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:15.99" />
                    <SPLIT distance="150" swimtime="00:01:59.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="622" swimtime="00:00:31.23" resultid="3078" heatid="7061" lane="6" entrytime="00:00:31.43" />
                <RESULT eventid="1406" points="351" swimtime="00:02:41.53" resultid="3079" heatid="7102" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="569" swimtime="00:01:10.67" resultid="3081" heatid="7163" lane="1" entrytime="00:01:12.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="3082">
              <RESULTS>
                <RESULT eventid="1134" points="75" swimtime="00:00:56.79" resultid="3083" heatid="6989" lane="9" entrytime="00:00:52.00" />
                <RESULT eventid="1194" points="146" swimtime="00:01:29.04" resultid="3084" heatid="7011" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="173" swimtime="00:00:40.18" resultid="3085" heatid="7038" lane="3" entrytime="00:00:38.00" />
                <RESULT comment="K-11 - Praca nóg w płaszczyźnie pionowej w dół" eventid="1286" status="DSQ" swimtime="00:01:10.42" resultid="3086" heatid="7053" lane="0" entrytime="00:00:56.00" />
                <RESULT eventid="1468" points="199" swimtime="00:00:35.79" resultid="5499" heatid="7125" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-28" firstname="Monika" gender="F" lastname="Figura" nation="POL" athleteid="3087">
              <RESULTS>
                <RESULT eventid="1453" points="359" swimtime="00:00:33.37" resultid="3088" heatid="7119" lane="6" entrytime="00:00:32.27" />
                <RESULT eventid="1483" points="288" swimtime="00:03:08.97" resultid="3089" heatid="7138" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                    <SPLIT distance="150" swimtime="00:02:21.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="3090">
              <RESULTS>
                <RESULT eventid="1179" points="219" swimtime="00:01:26.30" resultid="3091" heatid="7005" lane="8" entrytime="00:01:23.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="172" swimtime="00:00:45.04" resultid="3092" heatid="7032" lane="0" entrytime="00:00:43.25" />
                <RESULT eventid="1391" points="225" swimtime="00:03:27.24" resultid="3093" heatid="7093" lane="0" entrytime="00:03:21.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                    <SPLIT distance="100" swimtime="00:01:39.06" />
                    <SPLIT distance="150" swimtime="00:02:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="245" swimtime="00:00:37.88" resultid="3094" heatid="7117" lane="8" entrytime="00:00:37.18" />
                <RESULT eventid="1558" points="207" swimtime="00:06:44.15" resultid="3095" heatid="7166" lane="7" entrytime="00:06:15.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:27.14" />
                    <SPLIT distance="200" swimtime="00:03:19.19" />
                    <SPLIT distance="250" swimtime="00:04:10.98" />
                    <SPLIT distance="300" swimtime="00:05:02.67" />
                    <SPLIT distance="350" swimtime="00:05:54.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-31" firstname="Marianna" gender="F" lastname="Michalczyk" nation="POL" athleteid="3096">
              <RESULTS>
                <RESULT eventid="1058" points="311" swimtime="00:03:26.74" resultid="3236" heatid="6972" lane="6" entrytime="00:03:28.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:37.58" />
                    <SPLIT distance="150" swimtime="00:02:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="342" swimtime="00:00:35.83" resultid="3237" heatid="7033" lane="5" entrytime="00:00:35.57" />
                <RESULT eventid="1391" points="323" swimtime="00:03:03.69" resultid="3238" heatid="7094" lane="8" entrytime="00:03:01.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="306" swimtime="00:01:35.59" resultid="3239" heatid="7153" lane="3" entrytime="00:01:31.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-10" firstname="Alicja" gender="F" lastname="Stępniewska" nation="POL" athleteid="3101">
              <RESULTS>
                <RESULT eventid="1209" points="241" swimtime="00:03:15.68" resultid="3102" heatid="7024" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="150" swimtime="00:02:15.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="358" swimtime="00:00:35.29" resultid="3103" heatid="7034" lane="7" entrytime="00:00:33.90" />
                <RESULT eventid="1391" points="304" swimtime="00:03:07.44" resultid="3104" heatid="7094" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="328" swimtime="00:01:21.23" resultid="3105" heatid="7105" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-25" firstname="Barbara" gender="F" lastname="Ropa" nation="POL" athleteid="3106">
              <RESULTS>
                <RESULT eventid="1058" points="283" swimtime="00:03:33.23" resultid="3107" heatid="6972" lane="8" entrytime="00:03:34.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:41.33" />
                    <SPLIT distance="150" swimtime="00:02:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="278" swimtime="00:01:19.73" resultid="3108" heatid="7006" lane="0" entrytime="00:01:21.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="301" swimtime="00:00:44.44" resultid="3109" heatid="7049" lane="5" entrytime="00:00:45.06" />
                <RESULT eventid="1361" points="270" swimtime="00:02:54.77" resultid="3110" heatid="7079" lane="3" entrytime="00:03:02.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:24.39" />
                    <SPLIT distance="150" swimtime="00:02:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="275" swimtime="00:00:36.48" resultid="3111" heatid="7117" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1528" points="275" swimtime="00:01:39.03" resultid="3112" heatid="7152" lane="3" entrytime="00:01:42.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-15" firstname="Piotr" gender="M" lastname="Kober" nation="POL" athleteid="3113">
              <RESULTS>
                <RESULT eventid="1104" points="129" swimtime="00:04:11.75" resultid="3114" heatid="6975" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                    <SPLIT distance="100" swimtime="00:01:59.58" />
                    <SPLIT distance="150" swimtime="00:03:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="112" swimtime="00:00:49.80" resultid="3115" heatid="6991" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1194" points="159" swimtime="00:01:26.51" resultid="3116" heatid="7011" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="110" swimtime="00:01:48.38" resultid="3117" heatid="7068" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="127" swimtime="00:03:22.62" resultid="3118" heatid="7084" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:38.06" />
                    <SPLIT distance="150" swimtime="00:02:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="106" swimtime="00:04:00.32" resultid="3119" heatid="7097" lane="0" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.11" />
                    <SPLIT distance="100" swimtime="00:01:58.51" />
                    <SPLIT distance="150" swimtime="00:03:07.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-12-31" firstname="Dominik" gender="M" lastname="Matuzewicz" nation="POL" athleteid="3120">
              <RESULTS>
                <RESULT eventid="1468" points="497" swimtime="00:00:26.39" resultid="3121" heatid="7135" lane="7" entrytime="00:00:26.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-31" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="3122">
              <RESULTS>
                <RESULT eventid="1134" points="462" swimtime="00:00:31.09" resultid="3123" heatid="6997" lane="6" entrytime="00:00:30.30" />
                <RESULT comment="Rekord Polski Masters w kat. D /40-44/" eventid="1224" points="470" swimtime="00:02:23.33" resultid="3124" heatid="7029" lane="2" entrytime="00:02:25.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="514" swimtime="00:00:28.00" resultid="3125" heatid="7045" lane="7" entrytime="00:00:27.49" />
                <RESULT eventid="1376" points="460" swimtime="00:02:12.04" resultid="3126" heatid="7090" lane="1" entrytime="00:02:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="462" swimtime="00:01:04.42" resultid="3127" heatid="7112" lane="9" entrytime="00:01:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="381" swimtime="00:02:34.27" resultid="3128" heatid="7146" lane="6" entrytime="00:02:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:54.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-31" firstname="Monika" gender="F" lastname="Jarecka" nation="POL" athleteid="3129">
              <RESULTS>
                <RESULT eventid="1058" points="380" swimtime="00:03:13.37" resultid="3130" heatid="6973" lane="8" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:31.00" />
                    <SPLIT distance="150" swimtime="00:02:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="448" swimtime="00:00:38.93" resultid="3131" heatid="7051" lane="7" entrytime="00:00:38.50" />
                <RESULT eventid="1453" points="424" swimtime="00:00:31.58" resultid="3132" heatid="7119" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1528" points="404" swimtime="00:01:27.17" resultid="3133" heatid="7154" lane="3" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="3134">
              <RESULTS>
                <RESULT eventid="1104" points="354" swimtime="00:02:59.87" resultid="3135" heatid="6979" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:28.85" />
                    <SPLIT distance="150" swimtime="00:02:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="464" swimtime="00:01:00.56" resultid="3136" heatid="7018" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="444" swimtime="00:00:29.40" resultid="3137" heatid="7043" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1376" points="314" swimtime="00:02:30.05" resultid="3138" heatid="7086" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="446" swimtime="00:00:27.35" resultid="3139" heatid="7132" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1543" points="425" swimtime="00:01:17.88" resultid="3140" heatid="7162" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-02" firstname="Wojciech" gender="M" lastname="Czupryn" nation="POL" athleteid="3141">
              <RESULTS>
                <RESULT eventid="1104" points="158" swimtime="00:03:55.03" resultid="3142" heatid="6975" lane="2" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                    <SPLIT distance="100" swimtime="00:01:55.24" />
                    <SPLIT distance="150" swimtime="00:02:56.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="186" swimtime="00:01:22.15" resultid="3143" heatid="7012" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="130" swimtime="00:00:44.19" resultid="3144" heatid="7037" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1376" points="150" swimtime="00:03:11.90" resultid="3145" heatid="7084" lane="1" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:01:32.72" />
                    <SPLIT distance="150" swimtime="00:02:24.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="199" swimtime="00:00:35.79" resultid="3146" heatid="7122" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1573" points="156" swimtime="00:06:48.53" resultid="3147" heatid="7169" lane="7" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:37.17" />
                    <SPLIT distance="150" swimtime="00:02:30.27" />
                    <SPLIT distance="200" swimtime="00:03:24.13" />
                    <SPLIT distance="250" swimtime="00:04:17.20" />
                    <SPLIT distance="300" swimtime="00:05:11.21" />
                    <SPLIT distance="350" swimtime="00:06:03.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-01" firstname="Stanisław" gender="M" lastname="Fluder" nation="POL" athleteid="3148">
              <RESULTS>
                <RESULT eventid="1194" points="540" swimtime="00:00:57.58" resultid="3149" heatid="7022" lane="8" entrytime="00:00:57.30" />
                <RESULT eventid="1256" points="497" swimtime="00:00:28.31" resultid="3150" heatid="7044" lane="4" entrytime="00:00:28.30" />
                <RESULT eventid="1376" points="479" swimtime="00:02:10.32" resultid="3151" heatid="7090" lane="7" entrytime="00:02:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="491" swimtime="00:00:26.49" resultid="3152" heatid="7135" lane="1" entrytime="00:00:26.20" />
                <RESULT eventid="1573" points="470" swimtime="00:04:42.95" resultid="3153" heatid="7173" lane="5" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:43.70" />
                    <SPLIT distance="200" swimtime="00:02:19.98" />
                    <SPLIT distance="250" swimtime="00:02:55.69" />
                    <SPLIT distance="300" swimtime="00:03:32.08" />
                    <SPLIT distance="350" swimtime="00:04:08.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="3154">
              <RESULTS>
                <RESULT eventid="1134" points="255" swimtime="00:00:37.89" resultid="3155" heatid="6992" lane="7" entrytime="00:00:39.90" />
                <RESULT eventid="1194" points="334" swimtime="00:01:07.57" resultid="3156" heatid="7015" lane="1" entrytime="00:01:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="233" swimtime="00:01:24.32" resultid="3157" heatid="7069" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="321" swimtime="00:00:30.51" resultid="3159" heatid="7128" lane="8" entrytime="00:00:30.90" />
                <RESULT eventid="1573" points="280" swimtime="00:05:36.36" resultid="3160" heatid="7170" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                    <SPLIT distance="200" swimtime="00:02:43.99" />
                    <SPLIT distance="250" swimtime="00:03:27.80" />
                    <SPLIT distance="300" swimtime="00:04:11.87" />
                    <SPLIT distance="350" swimtime="00:04:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="285" swimtime="00:02:34.98" resultid="5493" heatid="7086" lane="9" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                    <SPLIT distance="150" swimtime="00:01:54.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-12-31" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="3161">
              <RESULTS>
                <RESULT eventid="1104" points="290" swimtime="00:03:12.28" resultid="3162" heatid="6978" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:34.03" />
                    <SPLIT distance="150" swimtime="00:02:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="274" swimtime="00:00:34.52" resultid="3163" heatid="7041" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1406" points="266" swimtime="00:02:57.21" resultid="3164" heatid="7100" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="230" swimtime="00:01:21.29" resultid="3165" heatid="7109" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="247" swimtime="00:05:50.57" resultid="3166" heatid="7171" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:09.02" />
                    <SPLIT distance="200" swimtime="00:02:54.65" />
                    <SPLIT distance="250" swimtime="00:03:39.32" />
                    <SPLIT distance="300" swimtime="00:04:23.86" />
                    <SPLIT distance="350" swimtime="00:05:08.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-09" firstname="Michał" gender="M" lastname="Sędrowski" nation="POL" athleteid="3167">
              <RESULTS>
                <RESULT eventid="1134" points="455" swimtime="00:00:31.25" resultid="3168" heatid="6996" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1316" points="380" swimtime="00:01:11.67" resultid="3169" heatid="7071" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3170" heatid="7100" lane="9" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="3171">
              <RESULTS>
                <RESULT eventid="1134" points="420" swimtime="00:00:32.08" resultid="3172" heatid="6995" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1194" points="496" swimtime="00:00:59.24" resultid="3173" heatid="7021" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="367" swimtime="00:01:12.54" resultid="3174" heatid="7071" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="382" swimtime="00:02:20.53" resultid="3175" heatid="7089" lane="2" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="457" swimtime="00:00:27.13" resultid="3176" heatid="7135" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1498" points="313" swimtime="00:02:44.83" resultid="3177" heatid="7145" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:06.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-31" firstname="Ewa" gender="F" lastname="Kosmol" nation="POL" athleteid="3178">
              <RESULTS>
                <RESULT eventid="1119" points="166" swimtime="00:00:49.23" resultid="3179" heatid="6983" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1179" points="145" swimtime="00:01:39.08" resultid="3180" heatid="7003" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="133" swimtime="00:00:49.02" resultid="3181" heatid="7031" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1361" points="122" swimtime="00:03:47.66" resultid="3182" heatid="7078" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                    <SPLIT distance="100" swimtime="00:01:50.81" />
                    <SPLIT distance="150" swimtime="00:02:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="146" swimtime="00:00:45.00" resultid="3183" heatid="7115" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1483" points="120" swimtime="00:04:12.79" resultid="3184" heatid="7137" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.82" />
                    <SPLIT distance="100" swimtime="00:02:03.19" />
                    <SPLIT distance="150" swimtime="00:03:08.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-05" firstname="Tomasz" gender="M" lastname="Bielan" nation="POL" athleteid="3185">
              <RESULTS>
                <RESULT eventid="1194" points="235" swimtime="00:01:15.98" resultid="3186" heatid="7013" lane="3" entrytime="00:01:14.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="234" swimtime="00:00:36.38" resultid="3187" heatid="7038" lane="1" entrytime="00:00:38.38" />
                <RESULT eventid="1468" points="259" swimtime="00:00:32.80" resultid="3188" heatid="7126" lane="2" entrytime="00:00:32.48" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-24" firstname="Ewa" gender="F" lastname="Szlagor" nation="POL" athleteid="3189">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. D /40-44/" eventid="1240" points="529" swimtime="00:00:30.99" resultid="3190" heatid="7030" lane="4" entrytime="00:00:59.00" />
                <RESULT comment="Rekord Polski Masters w kat. D /40-44/" eventid="1271" points="556" swimtime="00:00:36.22" resultid="3191" heatid="7051" lane="2" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="3192">
              <RESULTS>
                <RESULT eventid="1058" points="380" swimtime="00:03:13.31" resultid="3193" heatid="6973" lane="7" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:35.07" />
                    <SPLIT distance="150" swimtime="00:02:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="371" swimtime="00:00:41.46" resultid="3194" heatid="7050" lane="4" entrytime="00:00:40.50" />
                <RESULT eventid="1361" points="309" swimtime="00:02:47.07" resultid="3195" heatid="7080" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="150" swimtime="00:02:05.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="382" swimtime="00:01:28.79" resultid="3196" heatid="7154" lane="8" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-13" firstname="Ewa" gender="F" lastname="Krzyżanowska" nation="POL" athleteid="3197">
              <RESULTS>
                <RESULT eventid="1361" points="266" swimtime="00:02:55.49" resultid="3198" heatid="7079" lane="5" entrytime="00:03:02.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                    <SPLIT distance="150" swimtime="00:02:08.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="359" swimtime="00:00:33.36" resultid="3199" heatid="7118" lane="4" entrytime="00:00:33.29" />
                <RESULT eventid="1558" points="252" swimtime="00:06:18.38" resultid="3200" heatid="7166" lane="1" entrytime="00:06:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                    <SPLIT distance="200" swimtime="00:03:00.66" />
                    <SPLIT distance="250" swimtime="00:03:50.68" />
                    <SPLIT distance="300" swimtime="00:04:40.94" />
                    <SPLIT distance="350" swimtime="00:05:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-09-05" firstname="Joanna" gender="F" lastname="Maciąg" nation="POL" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1271" status="DNS" swimtime="00:00:00.00" resultid="3202" heatid="7049" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1528" points="274" swimtime="00:01:39.21" resultid="3203" heatid="7153" lane="7" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-07" firstname="Marta" gender="F" lastname="Paruszewska" nation="POL" athleteid="3204">
              <RESULTS>
                <RESULT eventid="1240" points="193" swimtime="00:00:43.33" resultid="3205" heatid="7031" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1361" points="211" swimtime="00:03:09.72" resultid="3206" heatid="7078" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:20.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="248" swimtime="00:00:37.75" resultid="3207" heatid="7116" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1558" points="182" swimtime="00:07:01.32" resultid="3208" heatid="7166" lane="9" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                    <SPLIT distance="150" swimtime="00:02:32.80" />
                    <SPLIT distance="200" swimtime="00:03:27.83" />
                    <SPLIT distance="250" swimtime="00:04:22.98" />
                    <SPLIT distance="300" swimtime="00:05:17.58" />
                    <SPLIT distance="350" swimtime="00:06:11.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="3209">
              <RESULTS>
                <RESULT eventid="1134" points="238" swimtime="00:00:38.76" resultid="3210" heatid="6992" lane="5" entrytime="00:00:38.63" />
                <RESULT eventid="1194" points="251" swimtime="00:01:14.28" resultid="3211" heatid="7014" lane="0" entrytime="00:01:14.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3212" heatid="7039" lane="2" entrytime="00:00:35.65" />
                <RESULT eventid="1286" points="349" swimtime="00:00:37.88" resultid="3213" heatid="7058" lane="7" entrytime="00:00:36.99" />
                <RESULT comment="O-4 - Przedwczwsny start" eventid="1468" status="DSQ" swimtime="00:00:31.45" resultid="3214" heatid="7128" lane="1" entrytime="00:00:30.73" />
                <RESULT eventid="1543" points="298" swimtime="00:01:27.67" resultid="3215" heatid="7159" lane="5" entrytime="00:01:25.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="3216">
              <RESULTS>
                <RESULT eventid="1179" points="120" swimtime="00:01:45.55" resultid="3217" heatid="7003" lane="1" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="107" swimtime="00:03:57.79" resultid="3218" heatid="7078" lane="9" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                    <SPLIT distance="100" swimtime="00:01:52.44" />
                    <SPLIT distance="150" swimtime="00:02:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="117" swimtime="00:00:48.42" resultid="3219" heatid="7115" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1558" points="117" swimtime="00:08:07.88" resultid="3220" heatid="7164" lane="6" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:53.93" />
                    <SPLIT distance="150" swimtime="00:02:57.20" />
                    <SPLIT distance="200" swimtime="00:04:01.42" />
                    <SPLIT distance="250" swimtime="00:05:03.03" />
                    <SPLIT distance="300" swimtime="00:06:07.35" />
                    <SPLIT distance="350" swimtime="00:07:08.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Bernard" gender="M" lastname="Wierzbik" nation="POL" athleteid="4513">
              <RESULTS>
                <RESULT eventid="1256" points="280" swimtime="00:00:34.26" resultid="4514" heatid="7040" lane="4" entrytime="00:00:33.54" />
                <RESULT eventid="1438" points="222" swimtime="00:01:22.21" resultid="4515" heatid="7109" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-01-01" firstname="Elżbieta" gender="F" lastname="Janik" nation="POL" athleteid="5494">
              <RESULTS>
                <RESULT eventid="1301" points="59" swimtime="00:02:29.22" resultid="5495" heatid="7063" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="28" swimtime="00:01:18.00" resultid="5496" heatid="7114" lane="8" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Wiesław" gender="M" lastname="Kurczyn" nation="POL" athleteid="6423">
              <RESULTS>
                <RESULT eventid="1286" points="95" swimtime="00:00:58.32" resultid="6424" heatid="7053" lane="9" entrytime="00:00:58.20" />
                <RESULT eventid="1468" points="52" swimtime="00:00:55.89" resultid="6425" heatid="7121" lane="4" entrytime="00:00:53.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. C /160-1199/" eventid="1164" points="453" swimtime="00:02:01.63" resultid="7215" heatid="7001" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:31.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3044" number="1" />
                    <RELAYPOSITION athleteid="3076" number="2" />
                    <RELAYPOSITION athleteid="3122" number="3" />
                    <RELAYPOSITION athleteid="3031" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="364" swimtime="00:01:58.81" resultid="7601" heatid="7075" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:00:59.67" />
                    <SPLIT distance="150" swimtime="00:01:30.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3167" number="1" />
                    <RELAYPOSITION athleteid="2994" number="2" />
                    <RELAYPOSITION athleteid="3031" number="3" />
                    <RELAYPOSITION athleteid="3076" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1164" status="DNF" swimtime="00:03:17.77" resultid="7216" heatid="7000" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:36.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3069" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3161" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3148" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3039" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="412" swimtime="00:01:53.95" resultid="7599" heatid="7076" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:00:58.33" />
                    <SPLIT distance="150" swimtime="00:01:28.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3044" number="1" />
                    <RELAYPOSITION athleteid="2972" number="2" />
                    <RELAYPOSITION athleteid="3154" number="3" />
                    <RELAYPOSITION athleteid="3148" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="475" swimtime="00:01:48.69" resultid="7600" heatid="7076" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="150" swimtime="00:01:22.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3069" number="1" />
                    <RELAYPOSITION athleteid="3122" number="2" />
                    <RELAYPOSITION athleteid="3039" number="3" />
                    <RELAYPOSITION athleteid="3171" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT comment="S-4 - Przedwczwsny start" eventid="1164" status="DSQ" swimtime="00:02:36.20" resultid="7217" heatid="6999" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3154" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3141" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3082" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3056" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="180" swimtime="00:02:30.17" resultid="7602" heatid="7074" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:54.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3001" number="1" />
                    <RELAYPOSITION athleteid="3113" number="2" />
                    <RELAYPOSITION athleteid="3141" number="3" />
                    <RELAYPOSITION athleteid="3082" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="372" swimtime="00:02:09.83" resultid="7212" heatid="7001" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:41.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3167" number="1" />
                    <RELAYPOSITION athleteid="2994" number="2" />
                    <RELAYPOSITION athleteid="2976" number="3" />
                    <RELAYPOSITION athleteid="2972" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1149" points="283" swimtime="00:02:41.63" resultid="7218" heatid="6998" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:04.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3009" number="1" />
                    <RELAYPOSITION athleteid="3106" number="2" />
                    <RELAYPOSITION athleteid="3096" number="3" />
                    <RELAYPOSITION athleteid="3090" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1331" points="449" swimtime="00:02:06.29" resultid="7603" heatid="7073" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:00.52" />
                    <SPLIT distance="150" swimtime="00:01:34.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3189" number="1" />
                    <RELAYPOSITION athleteid="3129" number="2" />
                    <RELAYPOSITION athleteid="3096" number="3" />
                    <RELAYPOSITION athleteid="3101" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1331" points="275" swimtime="00:02:28.67" resultid="7604" heatid="7073" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                    <SPLIT distance="150" swimtime="00:01:54.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3090" number="1" />
                    <RELAYPOSITION athleteid="3204" number="2" />
                    <RELAYPOSITION athleteid="3009" number="3" />
                    <RELAYPOSITION athleteid="3106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1513" points="379" swimtime="00:02:09.08" resultid="7612" heatid="7149" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:37.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3069" number="1" />
                    <RELAYPOSITION athleteid="3129" number="2" />
                    <RELAYPOSITION athleteid="3122" number="3" />
                    <RELAYPOSITION athleteid="3101" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" points="302" swimtime="00:02:19.19" resultid="7613" heatid="7149" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:01:45.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3087" number="1" />
                    <RELAYPOSITION athleteid="3161" number="2" />
                    <RELAYPOSITION athleteid="3148" number="3" />
                    <RELAYPOSITION athleteid="3096" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1513" points="219" swimtime="00:02:34.81" resultid="7614" heatid="7149" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:02.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3031" number="1" />
                    <RELAYPOSITION athleteid="3106" number="2" />
                    <RELAYPOSITION athleteid="3082" number="3" />
                    <RELAYPOSITION athleteid="3197" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1513" points="209" swimtime="00:02:37.28" resultid="7615" heatid="7149" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3154" number="1" />
                    <RELAYPOSITION athleteid="2994" number="2" />
                    <RELAYPOSITION athleteid="3090" number="3" />
                    <RELAYPOSITION athleteid="3204" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="DRZON" name="Drzonków" nation="POL" region="ZG">
          <CONTACT city="ŁĘŻYCA" email="PIOTRBARTA@O2.PL" name="BARTA PIOTR" phone="602347348" state="LUBUS" street="ODRZAŃSKA 21" zip="66016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="PIOTR" gender="M" lastname="BARTA" nation="POL" athleteid="3423">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. D /40-44/" eventid="1104" points="428" swimtime="00:02:48.83" resultid="3424" heatid="6979" lane="5" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:20.26" />
                    <SPLIT distance="150" swimtime="00:02:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="430" swimtime="00:00:35.33" resultid="3425" heatid="7059" lane="7" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1406" points="359" swimtime="00:02:40.30" resultid="3426" heatid="7101" lane="1" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="429" swimtime="00:01:17.67" resultid="3427" heatid="7162" lane="2" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="377" swimtime="00:05:04.51" resultid="3428" heatid="7171" lane="5" entrytime="00:05:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                    <SPLIT distance="200" swimtime="00:02:31.19" />
                    <SPLIT distance="250" swimtime="00:03:09.67" />
                    <SPLIT distance="300" swimtime="00:03:48.29" />
                    <SPLIT distance="350" swimtime="00:04:27.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSTA" name="MOTYL SENIOR MOSiR Stalowa Wola" nation="POL" region="PDK">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="15-8422562 wew.45" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="3430">
              <RESULTS>
                <RESULT eventid="1134" points="305" swimtime="00:00:35.69" resultid="3431" heatid="6995" lane="0" entrytime="00:00:34.10" />
                <RESULT eventid="1194" points="403" swimtime="00:01:03.46" resultid="3432" heatid="7018" lane="5" entrytime="00:01:03.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="343" swimtime="00:02:25.70" resultid="3433" heatid="7088" lane="5" entrytime="00:02:18.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="312" swimtime="00:02:48.03" resultid="3434" heatid="7101" lane="6" entrytime="00:02:43.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:17.09" />
                    <SPLIT distance="150" swimtime="00:02:08.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="404" swimtime="00:00:28.28" resultid="3435" heatid="7133" lane="1" entrytime="00:00:27.44" />
                <RESULT eventid="1573" points="329" swimtime="00:05:18.59" resultid="3436" heatid="7172" lane="3" entrytime="00:05:03.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:51.14" />
                    <SPLIT distance="200" swimtime="00:02:32.96" />
                    <SPLIT distance="250" swimtime="00:03:15.60" />
                    <SPLIT distance="300" swimtime="00:03:58.45" />
                    <SPLIT distance="350" swimtime="00:04:39.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="3437">
              <RESULTS>
                <RESULT eventid="1134" points="458" swimtime="00:00:31.18" resultid="3438" heatid="6996" lane="1" entrytime="00:00:31.67" />
                <RESULT eventid="1194" points="462" swimtime="00:01:00.66" resultid="3439" heatid="7020" lane="9" entrytime="00:01:01.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="344" swimtime="00:00:32.01" resultid="3440" heatid="7042" lane="1" entrytime="00:00:31.08" />
                <RESULT eventid="1316" points="405" swimtime="00:01:10.18" resultid="3441" heatid="7071" lane="3" entrytime="00:01:09.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="446" swimtime="00:00:27.36" resultid="3442" heatid="7132" lane="6" entrytime="00:00:27.61" />
                <RESULT eventid="1498" points="363" swimtime="00:02:36.83" resultid="3443" heatid="7145" lane="4" entrytime="00:02:37.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:01:58.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="3444">
              <RESULTS>
                <RESULT eventid="1224" points="466" swimtime="00:02:23.80" resultid="3445" heatid="7029" lane="3" entrytime="00:02:23.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:44.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="516" swimtime="00:00:27.96" resultid="3446" heatid="7045" lane="5" entrytime="00:00:27.30" />
                <RESULT eventid="1376" points="506" swimtime="00:02:07.92" resultid="3447" heatid="7090" lane="2" entrytime="00:02:08.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:02.34" />
                    <SPLIT distance="150" swimtime="00:01:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="532" swimtime="00:01:01.47" resultid="3448" heatid="7112" lane="7" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="500" swimtime="00:04:37.11" resultid="3449" heatid="7174" lane="6" entrytime="00:04:32.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                    <SPLIT distance="200" swimtime="00:02:17.31" />
                    <SPLIT distance="250" swimtime="00:02:53.21" />
                    <SPLIT distance="300" swimtime="00:03:29.22" />
                    <SPLIT distance="350" swimtime="00:04:04.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-07" firstname="Paweł" gender="M" lastname="Ciurko" nation="POL" athleteid="3450">
              <RESULTS>
                <RESULT eventid="1104" points="354" swimtime="00:02:59.96" resultid="3451" heatid="6980" lane="7" entrytime="00:02:45.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:02:13.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="170" swimtime="00:03:20.95" resultid="3452" heatid="7028" lane="1" entrytime="00:02:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:37.06" />
                    <SPLIT distance="150" swimtime="00:02:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="376" swimtime="00:00:36.93" resultid="3453" heatid="7059" lane="4" entrytime="00:00:35.11" />
                <RESULT eventid="1406" points="282" swimtime="00:02:53.82" resultid="3454" heatid="7100" lane="4" entrytime="00:02:45.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="150" swimtime="00:02:12.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="227" swimtime="00:01:21.64" resultid="3455" heatid="7110" lane="9" entrytime="00:01:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="369" swimtime="00:01:21.65" resultid="3456" heatid="7162" lane="5" entrytime="00:01:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="3457">
              <RESULTS>
                <RESULT eventid="1134" points="188" swimtime="00:00:41.96" resultid="3458" heatid="6989" lane="6" entrytime="00:00:48.94" />
                <RESULT eventid="1194" points="189" swimtime="00:01:21.72" resultid="3459" heatid="7012" lane="1" entrytime="00:01:21.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="172" swimtime="00:01:33.37" resultid="3460" heatid="7068" lane="8" entrytime="00:01:36.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="172" swimtime="00:03:24.91" resultid="3461" heatid="7096" lane="5" entrytime="00:03:38.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:42.32" />
                    <SPLIT distance="150" swimtime="00:02:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="264" swimtime="00:00:32.58" resultid="3462" heatid="7124" lane="4" entrytime="00:00:34.14" />
                <RESULT eventid="1498" points="152" swimtime="00:03:29.58" resultid="3463" heatid="7142" lane="6" entrytime="00:03:36.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                    <SPLIT distance="100" swimtime="00:01:45.39" />
                    <SPLIT distance="150" swimtime="00:02:39.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1194" points="299" swimtime="00:01:10.15" resultid="3465" heatid="7016" lane="0" entrytime="00:01:09.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="171" swimtime="00:03:20.56" resultid="3466" heatid="7027" lane="8" entrytime="00:03:18.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:31.81" />
                    <SPLIT distance="150" swimtime="00:02:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="3467" heatid="7086" lane="2" entrytime="00:02:38.11" />
                <RESULT eventid="1406" points="262" swimtime="00:02:58.13" resultid="3468" heatid="7099" lane="0" entrytime="00:02:56.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:18.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="3469" heatid="7108" lane="4" entrytime="00:01:22.41" />
                <RESULT eventid="1498" points="226" swimtime="00:03:03.60" resultid="3470" heatid="7144" lane="7" entrytime="00:02:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-04" firstname="Paweł" gender="M" lastname="Opaliński" nation="POL" athleteid="3471">
              <RESULTS>
                <RESULT eventid="1104" points="372" swimtime="00:02:57.01" resultid="3472" heatid="6979" lane="2" entrytime="00:03:00.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:08.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="408" swimtime="00:01:03.20" resultid="3473" heatid="7018" lane="4" entrytime="00:01:03.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="434" swimtime="00:00:35.21" resultid="3474" heatid="7058" lane="2" entrytime="00:00:36.59" />
                <RESULT eventid="1376" points="379" swimtime="00:02:20.86" resultid="3475" heatid="7088" lane="1" entrytime="00:02:20.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                    <SPLIT distance="150" swimtime="00:01:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="417" swimtime="00:01:18.36" resultid="3476" heatid="7162" lane="3" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="343" swimtime="00:05:14.09" resultid="3477" heatid="7172" lane="7" entrytime="00:05:15.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:51.10" />
                    <SPLIT distance="200" swimtime="00:02:31.34" />
                    <SPLIT distance="250" swimtime="00:03:12.53" />
                    <SPLIT distance="300" swimtime="00:03:54.04" />
                    <SPLIT distance="350" swimtime="00:04:36.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="3478">
              <RESULTS>
                <RESULT eventid="1104" points="290" swimtime="00:03:12.25" resultid="3479" heatid="6978" lane="1" entrytime="00:03:11.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:02:19.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3480" heatid="7027" lane="9" entrytime="00:03:22.10" />
                <RESULT eventid="1286" points="356" swimtime="00:00:37.60" resultid="3481" heatid="7058" lane="0" entrytime="00:00:37.15" />
                <RESULT eventid="1406" points="275" swimtime="00:02:55.20" resultid="3482" heatid="7098" lane="4" entrytime="00:02:57.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:14.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="234" swimtime="00:03:01.43" resultid="3483" heatid="7144" lane="0" entrytime="00:03:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="3484" heatid="7159" lane="3" entrytime="00:01:26.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="3485">
              <RESULTS>
                <RESULT eventid="1058" points="304" swimtime="00:03:28.18" resultid="3486" heatid="6972" lane="3" entrytime="00:03:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                    <SPLIT distance="100" swimtime="00:01:41.00" />
                    <SPLIT distance="150" swimtime="00:02:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="281" swimtime="00:01:19.42" resultid="3487" heatid="7006" lane="7" entrytime="00:01:18.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="310" swimtime="00:00:37.01" resultid="3488" heatid="7033" lane="1" entrytime="00:00:39.10" />
                <RESULT eventid="1391" points="296" swimtime="00:03:09.12" resultid="3489" heatid="7093" lane="2" entrytime="00:03:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:33.74" />
                    <SPLIT distance="150" swimtime="00:02:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="317" swimtime="00:00:34.80" resultid="3490" heatid="7117" lane="6" entrytime="00:00:36.10" />
                <RESULT eventid="1528" points="258" swimtime="00:01:41.20" resultid="3491" heatid="7153" lane="0" entrytime="00:01:36.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="3492">
              <RESULTS>
                <RESULT eventid="1134" points="264" swimtime="00:00:37.46" resultid="3493" heatid="6993" lane="0" entrytime="00:00:37.62" />
                <RESULT eventid="1224" points="152" swimtime="00:03:28.49" resultid="3494" heatid="7027" lane="0" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                    <SPLIT distance="150" swimtime="00:02:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="330" swimtime="00:00:32.44" resultid="3495" heatid="7041" lane="3" entrytime="00:00:32.75" />
                <RESULT eventid="1316" points="246" swimtime="00:01:22.80" resultid="3496" heatid="7069" lane="6" entrytime="00:01:24.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="241" swimtime="00:01:19.98" resultid="3497" heatid="7109" lane="1" entrytime="00:01:21.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="210" swimtime="00:03:08.17" resultid="3498" heatid="7144" lane="8" entrytime="00:03:00.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:01:31.34" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="3499">
              <RESULTS>
                <RESULT eventid="1104" points="421" swimtime="00:02:49.84" resultid="3500" heatid="6979" lane="4" entrytime="00:02:54.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:02:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="469" swimtime="00:00:34.31" resultid="3501" heatid="7060" lane="1" entrytime="00:00:34.80" />
                <RESULT eventid="1406" points="410" swimtime="00:02:33.39" resultid="3502" heatid="7101" lane="4" entrytime="00:02:40.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="319" swimtime="00:01:12.89" resultid="3503" heatid="7110" lane="2" entrytime="00:01:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="435" swimtime="00:01:17.29" resultid="3504" heatid="7162" lane="0" entrytime="00:01:19.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Paweł" gender="M" lastname="Cieśliński" nation="POL" athleteid="3505">
              <RESULTS>
                <RESULT eventid="1104" points="309" swimtime="00:03:08.22" resultid="3506" heatid="6978" lane="5" entrytime="00:03:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="150" swimtime="00:02:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="192" swimtime="00:03:13.12" resultid="3507" heatid="7028" lane="9" entrytime="00:03:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:35.06" />
                    <SPLIT distance="150" swimtime="00:02:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="310" swimtime="00:00:39.38" resultid="3508" heatid="7057" lane="1" entrytime="00:00:38.01" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3509" heatid="7098" lane="1" entrytime="00:03:05.10" />
                <RESULT eventid="1438" points="191" swimtime="00:01:26.36" resultid="3510" heatid="7109" lane="0" entrytime="00:01:22.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="301" swimtime="00:01:27.33" resultid="3511" heatid="7161" lane="2" entrytime="00:01:22.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="428" swimtime="00:02:03.92" resultid="3512" heatid="7000" lane="5" entrytime="00:02:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:35.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3437" number="1" />
                    <RELAYPOSITION athleteid="3499" number="2" />
                    <RELAYPOSITION athleteid="3444" number="3" />
                    <RELAYPOSITION athleteid="3471" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1164" points="285" swimtime="00:02:21.83" resultid="3513" heatid="7000" lane="7" entrytime="00:02:20.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:49.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3492" number="1" />
                    <RELAYPOSITION athleteid="3464" number="2" />
                    <RELAYPOSITION athleteid="3430" number="3" />
                    <RELAYPOSITION athleteid="3457" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1346" points="412" swimtime="00:01:53.97" resultid="3514" heatid="7076" lane="0" entrytime="00:01:52.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:00:56.30" />
                    <SPLIT distance="150" swimtime="00:01:26.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3437" number="1" />
                    <RELAYPOSITION athleteid="3499" number="2" />
                    <RELAYPOSITION athleteid="3478" number="3" />
                    <RELAYPOSITION athleteid="3471" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1346" points="337" swimtime="00:02:01.92" resultid="3515" heatid="7075" lane="7" entrytime="00:02:02.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:00.55" />
                    <SPLIT distance="150" swimtime="00:01:28.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3492" number="1" />
                    <RELAYPOSITION athleteid="3464" number="2" />
                    <RELAYPOSITION athleteid="3430" number="3" />
                    <RELAYPOSITION athleteid="3457" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="REWRO" name="Redeco Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="3532">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat B /30-34/" eventid="1058" points="581" swimtime="00:02:47.89" resultid="3533" heatid="6973" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. D /30-34/" eventid="1271" points="646" swimtime="00:00:34.46" resultid="3534" heatid="7051" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1528" points="591" swimtime="00:01:16.76" resultid="3535" heatid="7154" lane="5" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-28" firstname="Przemysław" gender="M" lastname="Matuszek" nation="POL" athleteid="3536">
              <RESULTS>
                <RESULT eventid="1194" points="366" swimtime="00:01:05.57" resultid="3537" heatid="7018" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="355" swimtime="00:00:31.65" resultid="3538" heatid="7043" lane="8" entrytime="00:00:30.50" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="3539" heatid="7085" lane="3" entrytime="00:02:45.00" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="3540" heatid="7110" lane="8" entrytime="00:01:15.00" />
                <RESULT eventid="1468" points="383" swimtime="00:00:28.77" resultid="3541" heatid="7131" lane="7" entrytime="00:00:28.28" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="3542" heatid="7160" lane="9" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Marta" gender="F" lastname="Frank" nation="POL" athleteid="3543">
              <RESULTS>
                <RESULT eventid="1119" points="373" swimtime="00:00:37.56" resultid="3544" heatid="6986" lane="0" entrytime="00:00:37.46" />
                <RESULT eventid="1179" points="297" swimtime="00:01:17.96" resultid="3545" heatid="7007" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="313" swimtime="00:01:25.55" resultid="3546" heatid="7065" lane="1" entrytime="00:01:20.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="298" swimtime="00:03:08.84" resultid="3547" heatid="7093" lane="4" entrytime="00:03:01.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:30.26" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="400" swimtime="00:00:32.19" resultid="3548" heatid="7120" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1483" points="279" swimtime="00:03:10.92" resultid="3549" heatid="7139" lane="1" entrytime="00:03:08.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:34.81" />
                    <SPLIT distance="150" swimtime="00:02:25.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Małgorzata" gender="F" lastname="Bogdan" nation="POL" athleteid="3550">
              <RESULTS>
                <RESULT eventid="1119" points="299" swimtime="00:00:40.46" resultid="3551" heatid="6985" lane="8" entrytime="00:00:40.09" />
                <RESULT eventid="1209" points="141" swimtime="00:03:53.56" resultid="3552" heatid="7024" lane="7" entrytime="00:03:54.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:52.66" />
                    <SPLIT distance="150" swimtime="00:02:52.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="262" swimtime="00:01:30.77" resultid="3553" heatid="7064" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="228" swimtime="00:03:26.43" resultid="3554" heatid="7093" lane="1" entrytime="00:03:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:37.98" />
                    <SPLIT distance="150" swimtime="00:02:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="143" swimtime="00:01:46.97" resultid="3555" heatid="7104" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="231" swimtime="00:03:23.26" resultid="3556" heatid="7138" lane="5" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                    <SPLIT distance="100" swimtime="00:01:37.81" />
                    <SPLIT distance="150" swimtime="00:02:30.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEOSI" name="Dęby Osielsko" nation="POL" region="MAZ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Adrian" gender="M" lastname="Teodorski" nation="POL" athleteid="3558">
              <RESULTS>
                <RESULT eventid="1194" points="512" swimtime="00:00:58.62" resultid="3559" heatid="7021" lane="7" entrytime="00:00:58.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="363" swimtime="00:02:36.23" resultid="3560" heatid="7029" lane="6" entrytime="00:02:23.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="505" swimtime="00:00:28.16" resultid="3561" heatid="7046" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1406" points="412" swimtime="00:02:33.19" resultid="3562" heatid="7103" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="463" swimtime="00:01:04.36" resultid="3563" heatid="7112" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POWAR" name="K.S Polonia Warszawa" nation="POL" region="MAZ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Lucjan" gender="M" lastname="Prządo" nation="POL" athleteid="3566">
              <RESULTS>
                <RESULT eventid="1104" points="113" swimtime="00:04:22.69" resultid="3567" heatid="6974" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.42" />
                    <SPLIT distance="100" swimtime="00:02:05.84" />
                    <SPLIT distance="150" swimtime="00:03:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="69" swimtime="00:00:58.39" resultid="3568" heatid="6987" lane="1" />
                <RESULT eventid="1286" points="120" swimtime="00:00:53.93" resultid="3569" heatid="7053" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1316" points="53" swimtime="00:02:17.57" resultid="3570" heatid="7066" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="56" swimtime="00:04:51.60" resultid="3571" heatid="7140" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.06" />
                    <SPLIT distance="100" swimtime="00:02:27.03" />
                    <SPLIT distance="150" swimtime="00:03:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="123" swimtime="00:01:57.61" resultid="3572" heatid="7156" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POSEI" name="Poseidonas" nation="LTU">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1977-01-28" firstname="Žalionis" gender="M" lastname="Giedrius" nation="LTU" athleteid="3630">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3631" heatid="7044" lane="6" entrytime="00:00:28.90" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="3632" heatid="7134" lane="2" entrytime="00:00:26.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Sergej" gender="M" lastname="Kolokolenkov" nation="LTU" athleteid="5477">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="5478" heatid="7014" lane="4" entrytime="00:01:12.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="5479" heatid="7041" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIWAR" name="Sinnet Club Warszawa" nation="POL" region="MAZ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1984-01-01" firstname="Joanna" gender="F" lastname="Janicka" nation="POL" athleteid="3634">
              <RESULTS>
                <RESULT eventid="1119" points="403" swimtime="00:00:36.63" resultid="3635" heatid="6986" lane="3" entrytime="00:00:34.89" />
                <RESULT eventid="1179" points="412" swimtime="00:01:09.96" resultid="3636" heatid="7008" lane="0" entrytime="00:01:08.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="343" swimtime="00:00:35.78" resultid="3637" heatid="7034" lane="2" entrytime="00:00:33.84" />
                <RESULT eventid="1361" points="349" swimtime="00:02:40.35" resultid="3638" heatid="7081" lane="7" entrytime="00:02:26.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="432" swimtime="00:00:31.38" resultid="3639" heatid="7120" lane="8" entrytime="00:00:30.59" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STPOZ" name="SSI Start Poznań" nation="POL" region="WLK">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="3641">
              <RESULTS>
                <RESULT eventid="1194" points="488" swimtime="00:00:59.57" resultid="3642" heatid="7020" lane="3" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="438" swimtime="00:02:14.25" resultid="3643" heatid="7089" lane="4" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="150" swimtime="00:01:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="388" swimtime="00:02:36.20" resultid="3644" heatid="7103" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:02:00.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="468" swimtime="00:00:26.93" resultid="3645" heatid="7134" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1573" points="429" swimtime="00:04:51.77" resultid="3646" heatid="7173" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                    <SPLIT distance="200" swimtime="00:02:24.59" />
                    <SPLIT distance="250" swimtime="00:03:02.81" />
                    <SPLIT distance="300" swimtime="00:03:39.81" />
                    <SPLIT distance="350" swimtime="00:04:16.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASZC" name="STP Masters Szczecinek" nation="POL" region="KUJ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1933-01-01" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="3648">
              <RESULTS>
                <RESULT eventid="1134" points="75" swimtime="00:00:56.86" resultid="3649" heatid="6988" lane="1" entrytime="00:00:57.00" />
                <RESULT eventid="1194" points="75" swimtime="00:01:50.97" resultid="3650" heatid="7010" lane="8" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="67" swimtime="00:02:07.62" resultid="3651" heatid="7067" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="71" swimtime="00:04:06.30" resultid="3652" heatid="7082" lane="4" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.48" />
                    <SPLIT distance="100" swimtime="00:01:59.04" />
                    <SPLIT distance="150" swimtime="00:03:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="61" swimtime="00:04:44.26" resultid="3653" heatid="7141" lane="2" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.02" />
                    <SPLIT distance="100" swimtime="00:02:20.90" />
                    <SPLIT distance="150" swimtime="00:03:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="71" swimtime="00:08:50.69" resultid="3654" heatid="7168" lane="2" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.42" />
                    <SPLIT distance="100" swimtime="00:02:02.47" />
                    <SPLIT distance="150" swimtime="00:03:09.22" />
                    <SPLIT distance="200" swimtime="00:04:17.67" />
                    <SPLIT distance="250" swimtime="00:05:26.29" />
                    <SPLIT distance="300" swimtime="00:06:35.32" />
                    <SPLIT distance="350" swimtime="00:07:44.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" name="Ts Masters Wisła Kraków" nation="POL" region="MAL">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="3656">
              <RESULTS>
                <RESULT eventid="1134" points="117" swimtime="00:00:49.06" resultid="3657" heatid="6988" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="1194" points="147" swimtime="00:01:28.70" resultid="3658" heatid="7010" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. L /80-84/" eventid="1256" points="79" swimtime="00:00:52.09" resultid="3659" heatid="7036" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1376" points="123" swimtime="00:03:24.75" resultid="3660" heatid="7083" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:34.33" />
                    <SPLIT distance="150" swimtime="00:02:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3661" heatid="7096" lane="8" entrytime="00:04:00.00" />
                <RESULT comment="Rekord Polski Masters w kat L /80-84/" eventid="1468" points="172" swimtime="00:00:37.55" resultid="3662" heatid="7123" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOTCZ" name="WOPR Tczew" nation="POL" region="POM">
          <CONTACT name="1" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="3665">
              <RESULTS>
                <RESULT eventid="1179" points="319" swimtime="00:01:16.14" resultid="3666" heatid="7006" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="271" swimtime="00:02:54.46" resultid="3667" heatid="7080" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="356" swimtime="00:00:33.48" resultid="3668" heatid="7119" lane="8" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZWAR" name="AZS-AWF Warszawa" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="ydiss@o2.pl" internet="www.azsawf.com" name="Kaczyński Jaczek" phone="698695042" state="MAZ" street="Marymoncka 34" zip="01-813" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" license="S00114100002" athleteid="3416">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. B /30-34/" eventid="1179" points="585" swimtime="00:01:02.25" resultid="3417" heatid="7008" lane="4" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="586" swimtime="00:00:29.95" resultid="3418" heatid="7034" lane="4" entrytime="00:00:29.80" />
                <RESULT comment="Rekord Polski Masters w kat. B /30-34/" eventid="1361" points="535" swimtime="00:02:19.11" resultid="3419" heatid="7081" lane="4" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:07.61" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat B /30-34/" eventid="1422" points="568" swimtime="00:01:07.67" resultid="3420" heatid="7105" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="543" swimtime="00:00:29.07" resultid="3421" heatid="7120" lane="5" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-16" firstname="Jacek" gender="M" lastname="Kaczyński" nation="POL" license="S00114200017" athleteid="3670">
              <RESULTS>
                <RESULT eventid="1256" points="626" swimtime="00:00:26.22" resultid="3671" heatid="7046" lane="5" entrytime="00:00:25.88" />
                <RESULT comment="Rekord Polski Masters w kat A /25-29/" eventid="1468" points="658" swimtime="00:00:24.03" resultid="3672" heatid="7136" lane="5" entrytime="00:00:24.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-14" firstname="Bartasz" gender="M" lastname="Krawczak" nation="POL" athleteid="5146" />
            <ATHLETE birthdate="1987-01-28" firstname="Jan" gender="M" lastname="Chmura" nation="POL" athleteid="5147" />
            <ATHLETE birthdate="1987-07-18" firstname="Damian" gender="M" lastname="Iwaniuk" nation="POL" athleteid="5148" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. A /100-119/" eventid="1346" points="642" swimtime="00:01:38.31" resultid="5149" heatid="7076" lane="4" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.05" />
                    <SPLIT distance="100" swimtime="00:00:50.05" />
                    <SPLIT distance="150" swimtime="00:01:14.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5146" number="1" />
                    <RELAYPOSITION athleteid="5147" number="2" />
                    <RELAYPOSITION athleteid="5148" number="3" />
                    <RELAYPOSITION athleteid="3670" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ORRAD" name="Orka Masters Radlin" nation="POL" region="SLA">
          <CONTACT city="Rydułtowy" email="zurekt@poczta.onet.pl" name="Żurczak Tomasz" state="ŚLĄSK" street="Gen.Maczka  12" zip="44-280" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="RUDOLF" gender="M" lastname="BUGLA" nation="POL" athleteid="3680">
              <RESULTS>
                <RESULT eventid="1134" points="97" swimtime="00:00:52.32" resultid="3681" heatid="6988" lane="4" entrytime="00:00:53.00" />
                <RESULT eventid="1224" points="68" swimtime="00:04:32.87" resultid="3682" heatid="7026" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.27" />
                    <SPLIT distance="100" swimtime="00:02:06.57" />
                    <SPLIT distance="150" swimtime="00:03:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="84" swimtime="00:01:58.19" resultid="3683" heatid="7067" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="81" swimtime="00:04:23.01" resultid="3684" heatid="7097" lane="8" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.46" />
                    <SPLIT distance="100" swimtime="00:02:08.59" />
                    <SPLIT distance="150" swimtime="00:03:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="83" swimtime="00:04:16.15" resultid="3685" heatid="7141" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.71" />
                    <SPLIT distance="100" swimtime="00:02:07.59" />
                    <SPLIT distance="150" swimtime="00:03:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="56" swimtime="00:09:32.52" resultid="3686" heatid="7168" lane="7" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.46" />
                    <SPLIT distance="100" swimtime="00:02:06.11" />
                    <SPLIT distance="150" swimtime="00:03:16.91" />
                    <SPLIT distance="200" swimtime="00:04:31.22" />
                    <SPLIT distance="250" swimtime="00:05:47.29" />
                    <SPLIT distance="300" swimtime="00:07:02.89" />
                    <SPLIT distance="350" swimtime="00:08:20.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-06-30" firstname="JAN" gender="M" lastname="KLAPSIA" nation="POL" athleteid="3687">
              <RESULTS>
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="3688" heatid="6988" lane="0" entrytime="00:01:04.00" />
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="3689" heatid="7009" lane="5" entrytime="00:02:45.00" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3690" heatid="7052" lane="3" entrytime="00:01:04.00" />
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="3691" heatid="7066" lane="1" entrytime="00:03:20.00" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="3692" heatid="7121" lane="2" entrytime="00:01:03.00" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="3693" heatid="7155" lane="2" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="JERZY" gender="M" lastname="CIECIOR" nation="POL" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="3695" heatid="6991" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="3696" heatid="7013" lane="9" entrytime="00:01:16.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3697" heatid="7039" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="3698" heatid="7085" lane="2" entrytime="00:02:47.00" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="3699" heatid="7108" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="3700" heatid="7143" lane="8" entrytime="00:03:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="MARIAN" gender="M" lastname="OTLIK" nation="POL" athleteid="3701">
              <RESULTS>
                <RESULT eventid="1134" points="210" swimtime="00:00:40.43" resultid="3702" heatid="6990" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1194" points="315" swimtime="00:01:08.88" resultid="3703" heatid="7010" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="226" swimtime="00:00:36.79" resultid="3704" heatid="7040" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1406" points="218" swimtime="00:03:09.30" resultid="3705" heatid="7098" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:32.99" />
                    <SPLIT distance="150" swimtime="00:02:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="296" swimtime="00:00:31.37" resultid="3706" heatid="7129" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1543" points="231" swimtime="00:01:35.47" resultid="3707" heatid="7158" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="LEON" gender="M" lastname="IRCZYK" nation="POL" athleteid="3708">
              <RESULTS>
                <RESULT eventid="1104" points="167" swimtime="00:03:50.96" resultid="3709" heatid="6975" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                    <SPLIT distance="100" swimtime="00:01:51.38" />
                    <SPLIT distance="150" swimtime="00:02:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="61" swimtime="00:04:43.22" resultid="3710" heatid="7025" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.45" />
                    <SPLIT distance="100" swimtime="00:02:15.20" />
                    <SPLIT distance="150" swimtime="00:03:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="93" swimtime="00:03:44.80" resultid="3711" heatid="7083" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.19" />
                    <SPLIT distance="100" swimtime="00:01:46.42" />
                    <SPLIT distance="150" swimtime="00:02:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="96" swimtime="00:04:08.71" resultid="3712" heatid="7096" lane="0" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.18" />
                    <SPLIT distance="100" swimtime="00:02:06.40" />
                    <SPLIT distance="150" swimtime="00:03:12.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="65" swimtime="00:02:03.72" resultid="3713" heatid="7106" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="147" swimtime="00:01:50.96" resultid="3714" heatid="7158" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="3715" heatid="6999" lane="4" entrytime="00:02:52.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3680" number="1" />
                    <RELAYPOSITION athleteid="3708" number="2" />
                    <RELAYPOSITION athleteid="3694" number="3" />
                    <RELAYPOSITION athleteid="3701" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="3716" heatid="7074" lane="5" entrytime="00:02:28.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3680" number="1" />
                    <RELAYPOSITION athleteid="3708" number="2" />
                    <RELAYPOSITION athleteid="3694" number="3" />
                    <RELAYPOSITION athleteid="3701" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SOKOL" name="Sokół Kolbuszowa" nation="POL" region="MAZ">
          <CONTACT name="Pietryka" phone="604620876" />
          <ATHLETES>
            <ATHLETE birthdate="1972-02-11" firstname="Witold" gender="M" lastname="Rado" nation="POL" athleteid="3725">
              <RESULTS>
                <RESULT eventid="1134" points="329" swimtime="00:00:34.79" resultid="3726" heatid="6995" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1194" points="348" swimtime="00:01:06.65" resultid="3727" heatid="7018" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="347" swimtime="00:00:31.89" resultid="3728" heatid="7043" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1406" points="315" swimtime="00:02:47.50" resultid="3729" heatid="7102" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:14.84" />
                    <SPLIT distance="150" swimtime="00:02:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="339" swimtime="00:01:11.40" resultid="3730" heatid="7110" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="310" swimtime="00:05:24.98" resultid="3731" heatid="7172" lane="9" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:56.63" />
                    <SPLIT distance="200" swimtime="00:02:38.87" />
                    <SPLIT distance="250" swimtime="00:03:21.57" />
                    <SPLIT distance="300" swimtime="00:04:03.32" />
                    <SPLIT distance="350" swimtime="00:04:44.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PIWAR" name="Uczniowski Klub Sportowy PINGWINY" nation="POL" region="MAZ" shortname="Uks Pingwiny">
          <CONTACT city="Warszawa" name="Perl Karol" />
          <ATHLETES>
            <ATHLETE birthdate="1959-07-30" firstname="Andrzej" gender="M" lastname="Błocki" nation="POL" athleteid="3733">
              <RESULTS>
                <RESULT eventid="1286" points="182" swimtime="00:00:47.06" resultid="3734" heatid="7055" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1468" points="164" swimtime="00:00:38.16" resultid="3735" heatid="7124" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-02" firstname="Grzegorz" gender="M" lastname="Krawczyk" nation="POL" athleteid="3736">
              <RESULTS>
                <RESULT eventid="1376" points="184" swimtime="00:02:59.02" resultid="3737" heatid="7084" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:25.26" />
                    <SPLIT distance="150" swimtime="00:02:13.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-18" firstname="Maciej" gender="M" lastname="Leszczyński" nation="POL" athleteid="3738">
              <RESULTS>
                <RESULT eventid="1104" points="165" swimtime="00:03:51.95" resultid="3739" heatid="6974" lane="4" entrytime="00:04:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:44.23" />
                    <SPLIT distance="150" swimtime="00:02:46.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="3740" heatid="7054" lane="3" entrytime="00:00:44.97" />
                <RESULT eventid="1543" points="165" swimtime="00:01:46.75" resultid="3741" heatid="7156" lane="2" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-09" firstname="Władysław" gender="M" lastname="Pawłowski" nation="POL" athleteid="3742">
              <RESULTS>
                <RESULT comment="K-12 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie" eventid="1104" status="DSQ" swimtime="00:04:11.43" resultid="3743" heatid="6974" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.68" />
                    <SPLIT distance="100" swimtime="00:02:03.24" />
                    <SPLIT distance="150" swimtime="00:03:08.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="168" swimtime="00:01:24.96" resultid="3744" heatid="7011" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="137" swimtime="00:00:43.41" resultid="3745" heatid="7037" lane="1" entrytime="00:00:41.00" />
                <RESULT comment="K-11 - Praca nóg w płaszczyźnie pionowej w dół" eventid="1286" status="DSQ" swimtime="00:00:49.64" resultid="3746" heatid="7054" lane="8" entrytime="00:00:46.00" />
                <RESULT eventid="1468" points="176" swimtime="00:00:37.31" resultid="3747" heatid="7123" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1543" points="149" swimtime="00:01:50.28" resultid="3748" heatid="7156" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-11-03" firstname="Karol" gender="M" lastname="Perl" nation="POL" athleteid="3749">
              <RESULTS>
                <RESULT eventid="1256" points="379" swimtime="00:00:30.97" resultid="3750" heatid="7040" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1376" points="334" swimtime="00:02:26.88" resultid="3751" heatid="7087" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="234" swimtime="00:03:04.96" resultid="3752" heatid="7101" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="150" swimtime="00:02:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="380" swimtime="00:00:28.86" resultid="3753" heatid="7129" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1573" points="315" swimtime="00:05:23.39" resultid="3754" heatid="7171" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:51.48" />
                    <SPLIT distance="200" swimtime="00:02:33.12" />
                    <SPLIT distance="250" swimtime="00:03:15.38" />
                    <SPLIT distance="300" swimtime="00:03:58.77" />
                    <SPLIT distance="350" swimtime="00:04:43.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-16" firstname="Małgorzata" gender="F" lastname="Sawicka" nation="POL" athleteid="3755">
              <RESULTS>
                <RESULT eventid="1119" points="243" swimtime="00:00:43.34" resultid="3756" heatid="6985" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1240" points="209" swimtime="00:00:42.19" resultid="3757" heatid="7033" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1301" points="207" swimtime="00:01:38.25" resultid="3758" heatid="7065" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="199" swimtime="00:03:33.58" resultid="3759" heatid="7139" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.18" />
                    <SPLIT distance="100" swimtime="00:01:41.34" />
                    <SPLIT distance="150" swimtime="00:02:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1346" points="236" swimtime="00:02:17.19" resultid="7595" heatid="7075" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:48.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3736" number="1" />
                    <RELAYPOSITION athleteid="3733" number="2" />
                    <RELAYPOSITION athleteid="3742" number="3" />
                    <RELAYPOSITION athleteid="3749" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MIELE" name="Mielec" nation="POL" region="PDK">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" athleteid="3761">
              <RESULTS>
                <RESULT eventid="1224" points="546" swimtime="00:02:16.35" resultid="3762" heatid="7029" lane="4" entrytime="00:02:16.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="458" swimtime="00:02:12.25" resultid="3763" heatid="7090" lane="8" entrytime="00:02:08.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="400" swimtime="00:02:34.65" resultid="3764" heatid="7103" lane="1" entrytime="00:02:26.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:02:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="456" swimtime="00:01:04.71" resultid="3765" heatid="7111" lane="4" entrytime="00:01:02.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="497" swimtime="00:04:37.82" resultid="3766" heatid="7174" lane="5" entrytime="00:04:29.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:42.26" />
                    <SPLIT distance="200" swimtime="00:02:17.61" />
                    <SPLIT distance="250" swimtime="00:02:53.72" />
                    <SPLIT distance="300" swimtime="00:03:29.48" />
                    <SPLIT distance="350" swimtime="00:04:04.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPLO" name="Płońsk Masters" nation="POL" region="MAZ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Alina" gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="3805">
              <RESULTS>
                <RESULT eventid="1119" points="42" swimtime="00:01:17.53" resultid="3806" heatid="6982" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1179" points="21" swimtime="00:03:06.37" resultid="3807" heatid="7003" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="16" swimtime="00:01:39.11" resultid="3808" heatid="7030" lane="2" entrytime="00:01:38.00" />
                <RESULT eventid="1301" points="38" swimtime="00:02:52.02" resultid="3809" heatid="7063" lane="9" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="39" swimtime="00:06:06.85" resultid="3810" heatid="7137" lane="1" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.38" />
                    <SPLIT distance="100" swimtime="00:03:01.39" />
                    <SPLIT distance="150" swimtime="00:04:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="34" swimtime="00:03:18.90" resultid="3811" heatid="7151" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SATCZ" name="Sambor Tczew" nation="POL" region="POM">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Kamila" gender="F" lastname="Ormianin" nation="POL" athleteid="3813">
              <RESULTS>
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="3814" heatid="7008" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1361" status="DNS" swimtime="00:00:00.00" resultid="3815" heatid="7081" lane="2" entrytime="00:02:25.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="3816" heatid="7120" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1558" status="DNS" swimtime="00:00:00.00" resultid="3817" heatid="7167" lane="6" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WORAD" name="Wodnik Radom" nation="POL" region="MAZ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Sebastian" gender="M" lastname="Pajdzik" nation="POL" athleteid="3819">
              <RESULTS>
                <RESULT eventid="1134" points="437" swimtime="00:00:31.66" resultid="3820" heatid="6997" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1316" points="441" swimtime="00:01:08.20" resultid="3821" heatid="7072" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3822" heatid="7102" lane="7" entrytime="00:02:35.00" />
                <RESULT eventid="1573" points="414" swimtime="00:04:55.21" resultid="3823" heatid="7173" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                    <SPLIT distance="200" swimtime="00:02:24.90" />
                    <SPLIT distance="250" swimtime="00:03:02.16" />
                    <SPLIT distance="300" swimtime="00:03:40.34" />
                    <SPLIT distance="350" swimtime="00:04:18.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKUT" name="WOPR Kutno" nation="POL" region="KUJ">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1932-01-01" firstname="Kazimierz" gender="M" lastname="From" nation="POL" athleteid="3825">
              <RESULTS>
                <RESULT eventid="1134" points="26" swimtime="00:01:20.78" resultid="3826" heatid="6987" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1194" points="39" swimtime="00:02:18.01" resultid="3827" heatid="7010" lane="0" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="26" swimtime="00:02:55.22" resultid="3828" heatid="7066" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="29" swimtime="00:05:28.84" resultid="3829" heatid="7082" lane="3" entrytime="00:04:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.34" />
                    <SPLIT distance="100" swimtime="00:02:32.80" />
                    <SPLIT distance="150" swimtime="00:04:02.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="45" swimtime="00:00:58.59" resultid="3830" heatid="7121" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1498" points="22" swimtime="00:06:37.31" resultid="3831" heatid="7140" lane="5" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.62" />
                    <SPLIT distance="100" swimtime="00:03:08.66" />
                    <SPLIT distance="150" swimtime="00:04:55.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASOP" name="Sopot Masters" nation="POL" region="POM">
          <CONTACT city="Gdańsk" email="puchalskaasia@wp.pl" name="Puchalska Joanna" phone="607035439" state="POMOR" street="Chłopska 10H/9" zip="80-399" />
          <ATHLETES>
            <ATHLETE birthdate="1964-08-04" firstname="Joanna" gender="F" lastname="Puchalska" nation="POL" athleteid="3835">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat E /45-49/" eventid="1058" points="416" swimtime="00:03:07.61" resultid="3836" heatid="6973" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:32.14" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1209" points="371" swimtime="00:02:49.48" resultid="3837" heatid="7024" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:18.78" />
                    <SPLIT distance="150" swimtime="00:02:02.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="383" swimtime="00:00:34.50" resultid="3838" heatid="7034" lane="9" entrytime="00:00:35.00" />
                <RESULT comment="Rekord Polski Masters w kat. E /45-49/" eventid="1391" points="420" swimtime="00:02:48.43" resultid="3839" heatid="7094" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:02:09.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat E /45-49/" eventid="1422" points="425" swimtime="00:01:14.53" resultid="3840" heatid="7105" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat E /45-49/" eventid="1528" points="410" swimtime="00:01:26.75" resultid="3841" heatid="7154" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TOTOR" name="Toruńczyk Masters Toruń" nation="POL" region="KUJ">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ -" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="3843">
              <RESULTS>
                <RESULT eventid="1194" points="498" swimtime="00:00:59.17" resultid="3844" heatid="7020" lane="5" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="384" swimtime="00:02:20.26" resultid="3845" heatid="7089" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="448" swimtime="00:00:27.32" resultid="3846" heatid="7133" lane="6" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="3847">
              <RESULTS>
                <RESULT eventid="1134" points="58" swimtime="00:01:02.03" resultid="3848" heatid="6988" lane="7" entrytime="00:00:56.52" />
                <RESULT eventid="1194" points="102" swimtime="00:01:40.13" resultid="3849" heatid="7010" lane="3" entrytime="00:01:34.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="3850" heatid="7067" lane="0" entrytime="00:02:07.42" />
                <RESULT eventid="1376" points="71" swimtime="00:04:06.05" resultid="3851" heatid="7083" lane="9" entrytime="00:03:51.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                    <SPLIT distance="100" swimtime="00:01:52.25" />
                    <SPLIT distance="150" swimtime="00:03:01.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="123" swimtime="00:00:41.96" resultid="3852" heatid="7123" lane="0" entrytime="00:00:39.54" />
                <RESULT eventid="1498" points="46" swimtime="00:05:11.93" resultid="3853" heatid="7141" lane="1" entrytime="00:04:45.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.87" />
                    <SPLIT distance="100" swimtime="00:02:33.74" />
                    <SPLIT distance="150" swimtime="00:03:55.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="3854">
              <RESULTS>
                <RESULT eventid="1119" points="306" swimtime="00:00:40.14" resultid="3855" heatid="6986" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1179" points="365" swimtime="00:01:12.84" resultid="3856" heatid="7008" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="282" swimtime="00:02:52.20" resultid="3857" heatid="7081" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:20.60" />
                    <SPLIT distance="150" swimtime="00:02:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="288" swimtime="00:03:10.93" resultid="3858" heatid="7094" lane="3" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="150" swimtime="00:02:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="255" swimtime="00:03:16.73" resultid="3859" heatid="7139" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:37.29" />
                    <SPLIT distance="150" swimtime="00:02:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="304" swimtime="00:05:55.65" resultid="3860" heatid="7167" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                    <SPLIT distance="150" swimtime="00:02:08.53" />
                    <SPLIT distance="200" swimtime="00:02:54.24" />
                    <SPLIT distance="250" swimtime="00:03:39.83" />
                    <SPLIT distance="300" swimtime="00:04:25.73" />
                    <SPLIT distance="350" swimtime="00:05:11.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-03" firstname="Artur" gender="M" lastname="Kłosiński" nation="POL" athleteid="3861">
              <RESULTS>
                <RESULT eventid="1134" points="318" swimtime="00:00:35.21" resultid="3862" heatid="6990" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1194" points="434" swimtime="00:01:01.94" resultid="3863" heatid="7021" lane="0" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="383" swimtime="00:00:36.70" resultid="3864" heatid="7059" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1376" points="356" swimtime="00:02:23.82" resultid="3865" heatid="7089" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="445" swimtime="00:00:27.38" resultid="3866" heatid="7135" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1543" points="326" swimtime="00:01:25.05" resultid="3867" heatid="7161" lane="9" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="3868">
              <RESULTS>
                <RESULT eventid="1134" points="206" swimtime="00:00:40.64" resultid="3869" heatid="6991" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1194" points="257" swimtime="00:01:13.69" resultid="3870" heatid="7014" lane="3" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="250" swimtime="00:00:35.59" resultid="3871" heatid="7040" lane="6" entrytime="00:00:34.50" />
                <RESULT eventid="1406" points="182" swimtime="00:03:20.80" resultid="3872" heatid="7097" lane="6" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:41.62" />
                    <SPLIT distance="150" swimtime="00:02:39.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="164" swimtime="00:01:30.94" resultid="3873" heatid="7108" lane="8" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="268" swimtime="00:00:32.43" resultid="3874" heatid="7128" lane="0" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-04" firstname="Karol" gender="M" lastname="Twarowski" nation="POL" athleteid="3875">
              <RESULTS>
                <RESULT eventid="1104" points="395" swimtime="00:02:53.48" resultid="3876" heatid="6980" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="501" swimtime="00:00:59.03" resultid="3877" heatid="7022" lane="0" entrytime="00:00:57.49" />
                <RESULT eventid="1376" points="453" swimtime="00:02:12.73" resultid="3878" heatid="7090" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="444" swimtime="00:02:29.36" resultid="3879" heatid="7103" lane="8" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:10.41" />
                    <SPLIT distance="150" swimtime="00:01:55.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="372" swimtime="00:02:35.61" resultid="3880" heatid="7146" lane="0" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="441" swimtime="00:04:49.12" resultid="3881" heatid="7173" lane="3" entrytime="00:04:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                    <SPLIT distance="150" swimtime="00:01:41.66" />
                    <SPLIT distance="200" swimtime="00:02:19.07" />
                    <SPLIT distance="250" swimtime="00:02:56.80" />
                    <SPLIT distance="300" swimtime="00:03:34.95" />
                    <SPLIT distance="350" swimtime="00:04:13.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="3882">
              <RESULTS>
                <RESULT eventid="1134" points="183" swimtime="00:00:42.32" resultid="3883" heatid="6992" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1224" points="205" swimtime="00:03:09.05" resultid="3884" heatid="7028" lane="0" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="325" swimtime="00:00:32.62" resultid="3885" heatid="7041" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="7099" lane="1" entrytime="00:02:55.00" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="3887" heatid="7110" lane="1" entrytime="00:01:14.50" />
                <RESULT eventid="1573" points="278" swimtime="00:05:36.95" resultid="3888" heatid="7171" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:05.16" />
                    <SPLIT distance="200" swimtime="00:02:49.23" />
                    <SPLIT distance="250" swimtime="00:03:33.38" />
                    <SPLIT distance="300" swimtime="00:04:15.03" />
                    <SPLIT distance="350" swimtime="00:04:56.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="3889">
              <RESULTS>
                <RESULT eventid="1104" points="150" swimtime="00:03:59.37" resultid="3890" heatid="6976" lane="0" entrytime="00:03:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="100" swimtime="00:01:50.50" />
                    <SPLIT distance="150" swimtime="00:02:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="96" swimtime="00:00:52.50" resultid="3891" heatid="6989" lane="2" entrytime="00:00:49.50" />
                <RESULT eventid="1286" points="182" swimtime="00:00:47.05" resultid="3892" heatid="7054" lane="1" entrytime="00:00:45.50" />
                <RESULT eventid="1316" points="88" swimtime="00:01:56.53" resultid="3893" heatid="7067" lane="7" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="93" swimtime="00:01:49.90" resultid="3894" heatid="7107" lane="6" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="150" swimtime="00:01:50.15" resultid="3895" heatid="7157" lane="9" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-08" firstname="Maciej" gender="M" lastname="Kuras" nation="POL" athleteid="3896">
              <RESULTS>
                <RESULT eventid="1134" points="284" swimtime="00:00:36.54" resultid="3897" heatid="6994" lane="7" entrytime="00:00:35.10" />
                <RESULT eventid="1256" points="348" swimtime="00:00:31.86" resultid="3898" heatid="7042" lane="6" entrytime="00:00:30.63" />
                <RESULT eventid="1316" points="293" swimtime="00:01:18.12" resultid="3899" heatid="7070" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="280" swimtime="00:02:51.03" resultid="3900" heatid="7145" lane="1" entrytime="00:02:43.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:02:06.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="3901">
              <RESULTS>
                <RESULT eventid="1104" points="114" swimtime="00:04:21.83" resultid="3902" heatid="6974" lane="5" entrytime="00:04:15.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                    <SPLIT distance="100" swimtime="00:02:00.66" />
                    <SPLIT distance="150" swimtime="00:03:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="105" swimtime="00:00:50.88" resultid="3903" heatid="6989" lane="0" entrytime="00:00:51.03" />
                <RESULT eventid="1286" points="140" swimtime="00:00:51.28" resultid="3904" heatid="7053" lane="5" entrytime="00:00:48.02" />
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="3905" heatid="7067" lane="2" entrytime="00:01:56.23" />
                <RESULT eventid="1543" points="124" swimtime="00:01:57.36" resultid="3906" heatid="7156" lane="7" entrytime="00:01:54.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="3907">
              <RESULTS>
                <RESULT eventid="1194" points="122" swimtime="00:01:34.40" resultid="6691" heatid="7012" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="6692" heatid="7037" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="6693" heatid="7107" lane="4" entrytime="00:01:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-27" firstname="Magdalena" gender="F" lastname="Rogozińska" nation="POL" athleteid="3911">
              <RESULTS>
                <RESULT eventid="1058" points="287" swimtime="00:03:32.37" resultid="3912" heatid="6972" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="100" swimtime="00:01:42.65" />
                    <SPLIT distance="150" swimtime="00:02:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="307" swimtime="00:00:40.09" resultid="3913" heatid="6985" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1240" points="275" swimtime="00:00:38.55" resultid="3914" heatid="7033" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1271" points="364" swimtime="00:00:41.72" resultid="3915" heatid="7050" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1453" points="339" swimtime="00:00:34.00" resultid="3916" heatid="7119" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1528" points="305" swimtime="00:01:35.65" resultid="3917" heatid="7153" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Maciej" gender="M" lastname="Walenta" nation="POL" athleteid="3918">
              <RESULTS>
                <RESULT eventid="1134" points="402" swimtime="00:00:32.57" resultid="3919" heatid="6994" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1194" points="456" swimtime="00:01:00.91" resultid="3920" heatid="7018" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="420" swimtime="00:00:29.93" resultid="3921" heatid="7042" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1286" points="442" swimtime="00:00:35.01" resultid="3922" heatid="7060" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1468" points="428" swimtime="00:00:27.74" resultid="3923" heatid="7134" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1543" points="364" swimtime="00:01:21.98" resultid="3924" heatid="7162" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="3925" heatid="6999" lane="3" entrytime="00:03:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3901" number="1" />
                    <RELAYPOSITION athleteid="3889" number="2" />
                    <RELAYPOSITION athleteid="3868" number="3" />
                    <RELAYPOSITION athleteid="3847" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1346" points="455" swimtime="00:01:50.30" resultid="3926" heatid="7076" lane="2" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                    <SPLIT distance="100" swimtime="00:00:53.08" />
                    <SPLIT distance="150" swimtime="00:01:22.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3843" number="1" />
                    <RELAYPOSITION athleteid="3875" number="2" />
                    <RELAYPOSITION athleteid="3882" number="3" />
                    <RELAYPOSITION athleteid="3861" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MACHE" name="Masters Chełm" nation="POL" region="LBL">
          <CONTACT city="Chełm" email="elzbietadz@gmail.com" name="Dziwisz Elżbieta" state="LUB" street="Lubelska 139 D/13" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1941-11-10" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="3936">
              <RESULTS>
                <RESULT eventid="1104" points="118" swimtime="00:04:19.39" resultid="3937" heatid="6975" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.19" />
                    <SPLIT distance="100" swimtime="00:02:07.10" />
                    <SPLIT distance="150" swimtime="00:03:15.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="54" swimtime="00:04:53.89" resultid="3938" heatid="7025" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.76" />
                    <SPLIT distance="100" swimtime="00:02:24.36" />
                    <SPLIT distance="150" swimtime="00:03:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="96" swimtime="00:00:48.91" resultid="3939" heatid="7036" lane="8" entrytime="00:00:56.00" />
                <RESULT eventid="1286" points="188" swimtime="00:00:46.52" resultid="3940" heatid="7055" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="1438" points="74" swimtime="00:01:58.50" resultid="3941" heatid="7106" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="140" swimtime="00:01:52.74" resultid="3942" heatid="7156" lane="5" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Wiesław" gender="M" lastname="Wepa" nation="POL" athleteid="3943">
              <RESULTS>
                <RESULT eventid="1104" points="127" swimtime="00:04:13.14" resultid="3944" heatid="6975" lane="0" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.20" />
                    <SPLIT distance="100" swimtime="00:01:53.21" />
                    <SPLIT distance="150" swimtime="00:03:02.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="114" swimtime="00:01:36.57" resultid="3945" heatid="7009" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="80" swimtime="00:00:51.94" resultid="3946" heatid="7036" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1286" points="155" swimtime="00:00:49.64" resultid="3947" heatid="7054" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1468" points="136" swimtime="00:00:40.59" resultid="3948" heatid="7123" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1543" points="144" swimtime="00:01:51.60" resultid="3949" heatid="7156" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1926-01-01" firstname="Barbara" gender="F" lastname="Korol" nation="POL" athleteid="3950">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat.M /85-89/" eventid="1119" points="15" swimtime="00:01:47.61" resultid="3951" heatid="6981" lane="3" />
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="3952" heatid="7002" lane="7" />
                <RESULT eventid="1301" points="12" swimtime="00:04:08.41" resultid="3953" heatid="7062" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="7" swimtime="00:01:58.72" resultid="3954" heatid="7113" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Hanna" gender="F" lastname="Wepa" nation="POL" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1058" points="77" swimtime="00:05:28.97" resultid="3956" heatid="6970" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.78" />
                    <SPLIT distance="100" swimtime="00:02:38.82" />
                    <SPLIT distance="150" swimtime="00:04:03.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="3957" heatid="6981" lane="7" />
                <RESULT eventid="1271" points="65" swimtime="00:01:13.85" resultid="3958" heatid="7047" lane="3" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3959" heatid="7062" lane="3" />
                <RESULT eventid="1453" points="29" swimtime="00:01:16.55" resultid="3960" heatid="7113" lane="4" />
                <RESULT eventid="1528" points="64" swimtime="00:02:40.69" resultid="7625" heatid="7150" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Elżbieta" gender="F" lastname="Dziwisz" nation="POL" athleteid="3961">
              <RESULTS>
                <RESULT eventid="1058" points="105" swimtime="00:04:56.72" resultid="3962" heatid="6971" lane="9" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.30" />
                    <SPLIT distance="100" swimtime="00:02:22.13" />
                    <SPLIT distance="150" swimtime="00:03:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="97" swimtime="00:00:58.88" resultid="3963" heatid="6982" lane="7" entrytime="00:01:03.00" />
                <RESULT eventid="1271" points="101" swimtime="00:01:03.83" resultid="3964" heatid="7048" lane="3" entrytime="00:00:58.00" />
                <RESULT eventid="1301" points="91" swimtime="00:02:09.08" resultid="3965" heatid="7063" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="100" swimtime="00:04:28.86" resultid="3966" heatid="7137" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.64" />
                    <SPLIT distance="100" swimtime="00:02:11.48" />
                    <SPLIT distance="150" swimtime="00:03:19.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="97" swimtime="00:02:19.84" resultid="3967" heatid="7152" lane="9" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Alicja" gender="F" lastname="Wątrobińska" nation="POL" athleteid="3968">
              <RESULTS>
                <RESULT eventid="1119" points="42" swimtime="00:01:17.77" resultid="3969" heatid="6981" lane="2" />
                <RESULT eventid="1179" points="55" swimtime="00:02:16.65" resultid="3970" heatid="7002" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="75" swimtime="00:01:10.46" resultid="3971" heatid="7047" lane="5" />
                <RESULT eventid="1301" points="37" swimtime="00:02:53.44" resultid="3972" heatid="7062" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="66" swimtime="00:00:58.47" resultid="3973" heatid="7113" lane="5" />
                <RESULT eventid="1528" points="63" swimtime="00:02:41.59" resultid="3974" heatid="7150" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1149" points="40" swimtime="00:05:08.26" resultid="3975" heatid="6998" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:52.14" />
                    <SPLIT distance="100" swimtime="00:03:03.32" />
                    <SPLIT distance="150" swimtime="00:04:17.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3950" number="1" />
                    <RELAYPOSITION athleteid="3955" number="2" />
                    <RELAYPOSITION athleteid="3968" number="3" />
                    <RELAYPOSITION athleteid="3961" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1513" points="57" swimtime="00:04:01.69" resultid="3976" heatid="7147" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.44" />
                    <SPLIT distance="100" swimtime="00:02:11.23" />
                    <SPLIT distance="150" swimtime="00:03:05.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3943" number="1" />
                    <RELAYPOSITION athleteid="3955" number="2" />
                    <RELAYPOSITION athleteid="3936" number="3" />
                    <RELAYPOSITION athleteid="3968" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAGDY" name="Gdynia Masters" nation="POL" region="POM">
          <CONTACT email="misiek@am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1944-01-01" firstname="Stefania" gender="F" lastname="Kowalska" nation="POL" athleteid="3980">
              <RESULTS>
                <RESULT eventid="1058" points="98" swimtime="00:05:03.74" resultid="3981" heatid="6970" lane="4" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.94" />
                    <SPLIT distance="100" swimtime="00:02:27.73" />
                    <SPLIT distance="150" swimtime="00:03:48.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="61" swimtime="00:02:12.13" resultid="3982" heatid="7003" lane="0" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="53" swimtime="00:01:06.66" resultid="3983" heatid="7030" lane="5" entrytime="00:01:02.00" />
                <RESULT eventid="1391" points="55" swimtime="00:05:31.67" resultid="3984" heatid="7091" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.36" />
                    <SPLIT distance="100" swimtime="00:02:50.73" />
                    <SPLIT distance="150" swimtime="00:04:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="73" swimtime="00:00:56.66" resultid="3985" heatid="7115" lane="8" entrytime="00:00:53.00" />
                <RESULT eventid="1528" points="99" swimtime="00:02:19.09" resultid="3986" heatid="7151" lane="2" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-01-01" firstname="Danuta" gender="F" lastname="Szczepańska" nation="POL" athleteid="3987">
              <RESULTS>
                <RESULT eventid="1119" points="186" swimtime="00:00:47.35" resultid="3988" heatid="6983" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="1453" points="197" swimtime="00:00:40.72" resultid="3989" heatid="7115" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="3990">
              <RESULTS>
                <RESULT eventid="1119" points="227" swimtime="00:00:44.30" resultid="3991" heatid="6985" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1179" points="206" swimtime="00:01:28.14" resultid="3992" heatid="7004" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="175" swimtime="00:00:44.79" resultid="3993" heatid="7032" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1301" points="184" swimtime="00:01:42.14" resultid="3994" heatid="7064" lane="9" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="248" swimtime="00:00:37.73" resultid="3995" heatid="7117" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1483" points="170" swimtime="00:03:44.93" resultid="3996" heatid="7138" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="150" swimtime="00:02:48.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="3997">
              <RESULTS>
                <RESULT eventid="1104" points="158" swimtime="00:03:55.32" resultid="3998" heatid="6976" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:49.52" />
                    <SPLIT distance="150" swimtime="00:02:53.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="138" swimtime="00:01:30.63" resultid="3999" heatid="7012" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="240" swimtime="00:00:42.91" resultid="4000" heatid="7055" lane="3" entrytime="00:00:42.30" />
                <RESULT eventid="1406" points="128" swimtime="00:03:45.75" resultid="4001" heatid="7097" lane="9" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:48.13" />
                    <SPLIT distance="150" swimtime="00:02:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="162" swimtime="00:00:38.32" resultid="4002" heatid="7124" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1543" points="185" swimtime="00:01:42.77" resultid="4003" heatid="7157" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Władysław" gender="M" lastname="Kurylczyk" nation="POL" athleteid="4004">
              <RESULTS>
                <RESULT eventid="1134" points="111" swimtime="00:00:49.88" resultid="4005" heatid="6991" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1194" points="145" swimtime="00:01:29.26" resultid="4006" heatid="7011" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4007" heatid="7037" lane="3" entrytime="00:00:40.00" />
                <RESULT comment="K-14 - Dotknięcie ściany jedną ręką przy nawrocie" eventid="1406" status="DSQ" swimtime="00:04:08.68" resultid="4008" heatid="7097" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:50.96" />
                    <SPLIT distance="150" swimtime="00:03:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="179" swimtime="00:00:37.05" resultid="4009" heatid="7124" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1543" points="187" swimtime="00:01:42.35" resultid="4010" heatid="7157" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Maja" gender="F" lastname="Szaduro" nation="POL" athleteid="4011">
              <RESULTS>
                <RESULT eventid="1058" points="248" swimtime="00:03:42.85" resultid="4012" heatid="6972" lane="0" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:41.41" />
                    <SPLIT distance="150" swimtime="00:02:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="268" swimtime="00:00:46.22" resultid="4013" heatid="7049" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1391" points="135" swimtime="00:04:05.89" resultid="4014" heatid="7092" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:53.92" />
                    <SPLIT distance="150" swimtime="00:02:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="276" swimtime="00:01:38.98" resultid="4015" heatid="7152" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="4016">
              <RESULTS>
                <RESULT eventid="1119" points="151" swimtime="00:00:50.71" resultid="4017" heatid="6982" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="1209" points="77" swimtime="00:04:45.34" resultid="4018" heatid="7023" lane="5" entrytime="00:04:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.67" />
                    <SPLIT distance="100" swimtime="00:02:15.47" />
                    <SPLIT distance="150" swimtime="00:03:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="72" swimtime="00:01:00.24" resultid="4019" heatid="7030" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1391" points="98" swimtime="00:04:33.38" resultid="4020" heatid="7091" lane="4" entrytime="00:04:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.68" />
                    <SPLIT distance="100" swimtime="00:02:11.75" />
                    <SPLIT distance="150" swimtime="00:03:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="68" swimtime="00:02:16.71" resultid="4021" heatid="7104" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="114" swimtime="00:02:12.65" resultid="4022" heatid="7152" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Renata" gender="F" lastname="Polańczyk" nation="POL" athleteid="4023">
              <RESULTS>
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="4024" heatid="7004" lane="1" entrytime="00:01:29.95" />
                <RESULT eventid="1209" points="120" swimtime="00:04:06.62" resultid="4025" heatid="7024" lane="8" entrytime="00:03:59.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                    <SPLIT distance="100" swimtime="00:01:54.38" />
                    <SPLIT distance="150" swimtime="00:03:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="193" swimtime="00:01:40.56" resultid="4026" heatid="7064" lane="8" entrytime="00:01:36.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="199" swimtime="00:03:33.62" resultid="4028" heatid="7138" lane="2" entrytime="00:03:25.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                    <SPLIT distance="100" swimtime="00:01:45.02" />
                    <SPLIT distance="150" swimtime="00:02:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="186" swimtime="00:06:58.57" resultid="4029" heatid="7165" lane="3" entrytime="00:06:46.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:35.71" />
                    <SPLIT distance="150" swimtime="00:02:29.45" />
                    <SPLIT distance="200" swimtime="00:03:23.68" />
                    <SPLIT distance="250" swimtime="00:04:18.10" />
                    <SPLIT distance="300" swimtime="00:05:13.15" />
                    <SPLIT distance="350" swimtime="00:06:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="160" swimtime="00:03:52.22" resultid="5650" heatid="7092" lane="1" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="100" swimtime="00:01:45.64" />
                    <SPLIT distance="150" swimtime="00:03:02.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="4030">
              <RESULTS>
                <RESULT eventid="1104" points="157" swimtime="00:03:55.71" resultid="4031" heatid="6975" lane="7" entrytime="00:03:53.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                    <SPLIT distance="100" swimtime="00:01:54.30" />
                    <SPLIT distance="150" swimtime="00:02:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="188" swimtime="00:00:46.49" resultid="4032" heatid="7054" lane="0" entrytime="00:00:46.04" />
                <RESULT eventid="1543" points="149" swimtime="00:01:50.47" resultid="4033" heatid="7156" lane="4" entrytime="00:01:46.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="Mazurek" nation="POL" athleteid="4034">
              <RESULTS>
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="4035" heatid="6984" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1179" points="253" swimtime="00:01:22.27" resultid="4036" heatid="7005" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="239" swimtime="00:00:40.39" resultid="4037" heatid="7032" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1271" points="338" swimtime="00:00:42.77" resultid="4038" heatid="7050" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1422" points="168" swimtime="00:01:41.55" resultid="4039" heatid="7105" lane="0" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="266" swimtime="00:01:40.17" resultid="4040" heatid="7153" lane="8" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Zuzanna" gender="F" lastname="Drążkiewicz" nation="POL" athleteid="4041">
              <RESULTS>
                <RESULT eventid="1179" status="DNF" swimtime="00:00:00.00" resultid="4042" heatid="7002" lane="6" entrytime="00:02:26.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="57" swimtime="00:01:17.36" resultid="4043" heatid="7048" lane="8" entrytime="00:01:18.67" />
                <RESULT eventid="1453" points="48" swimtime="00:01:05.24" resultid="4044" heatid="7114" lane="4" entrytime="00:00:58.56" />
                <RESULT eventid="1528" points="58" swimtime="00:02:45.70" resultid="4045" heatid="7151" lane="8" entrytime="00:02:56.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="4046">
              <RESULTS>
                <RESULT eventid="1058" points="202" swimtime="00:03:58.65" resultid="4047" heatid="6971" lane="6" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.60" />
                    <SPLIT distance="100" swimtime="00:01:56.16" />
                    <SPLIT distance="150" swimtime="00:02:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="167" swimtime="00:01:34.44" resultid="4048" heatid="7004" lane="0" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="144" swimtime="00:00:47.77" resultid="4049" heatid="7031" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1422" points="114" swimtime="00:01:55.40" resultid="4051" heatid="7104" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="170" swimtime="00:01:56.23" resultid="4052" heatid="7152" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Anna" gender="F" lastname="Krzysztofik" nation="POL" athleteid="4053">
              <RESULTS>
                <RESULT eventid="1058" points="212" swimtime="00:03:54.81" resultid="4054" heatid="6971" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.69" />
                    <SPLIT distance="100" swimtime="00:01:53.22" />
                    <SPLIT distance="150" swimtime="00:02:54.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="4055" heatid="6984" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1301" points="162" swimtime="00:01:46.60" resultid="4056" heatid="7063" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="160" swimtime="00:03:49.86" resultid="4057" heatid="7138" lane="9" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                    <SPLIT distance="100" swimtime="00:01:53.74" />
                    <SPLIT distance="150" swimtime="00:02:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="184" swimtime="00:01:53.26" resultid="4058" heatid="7152" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Magdalena" gender="F" lastname="Majewska" nation="POL" athleteid="4059">
              <RESULTS>
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="4060" heatid="6984" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1453" points="164" swimtime="00:00:43.28" resultid="4061" heatid="7116" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1149" points="184" swimtime="00:03:06.34" resultid="7591" heatid="6998" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:42.86" />
                    <SPLIT distance="150" swimtime="00:02:24.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3990" number="1" />
                    <RELAYPOSITION athleteid="3980" number="2" />
                    <RELAYPOSITION athleteid="4034" number="3" />
                    <RELAYPOSITION athleteid="4023" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="146" swimtime="00:03:03.57" resultid="4063" heatid="7073" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:41.03" />
                    <SPLIT distance="150" swimtime="00:02:25.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4034" number="1" />
                    <RELAYPOSITION athleteid="4023" number="2" />
                    <RELAYPOSITION athleteid="3987" number="3" />
                    <RELAYPOSITION athleteid="3980" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1513" points="104" swimtime="00:03:18.23" resultid="4062" heatid="7148" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.95" />
                    <SPLIT distance="100" swimtime="00:01:37.10" />
                    <SPLIT distance="150" swimtime="00:02:23.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3987" number="1" />
                    <RELAYPOSITION athleteid="4030" number="2" />
                    <RELAYPOSITION athleteid="3997" number="3" />
                    <RELAYPOSITION athleteid="3980" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" name="TS Olimpia Poznań" nation="POL" region="WIE">
          <CONTACT name="Pieteraszewski Zbigniew" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="4076">
              <RESULTS>
                <RESULT eventid="1179" points="194" swimtime="00:01:29.94" resultid="4077" heatid="7004" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="156" swimtime="00:00:46.51" resultid="4078" heatid="7031" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1391" points="156" swimtime="00:03:54.16" resultid="4079" heatid="7092" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                    <SPLIT distance="100" swimtime="00:01:54.80" />
                    <SPLIT distance="150" swimtime="00:03:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="238" swimtime="00:00:38.25" resultid="4080" heatid="7116" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1558" points="205" swimtime="00:06:45.52" resultid="4081" heatid="7165" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="150" swimtime="00:02:30.14" />
                    <SPLIT distance="200" swimtime="00:03:22.92" />
                    <SPLIT distance="250" swimtime="00:04:13.90" />
                    <SPLIT distance="300" swimtime="00:05:05.42" />
                    <SPLIT distance="350" swimtime="00:05:56.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="4082">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat G /55-59/" eventid="1058" points="332" swimtime="00:03:22.22" resultid="4083" heatid="6972" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:37.23" />
                    <SPLIT distance="150" swimtime="00:02:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. G /55-59/" eventid="1271" points="319" swimtime="00:00:43.59" resultid="4084" heatid="7050" lane="8" entrytime="00:00:43.00" />
                <RESULT comment="Rekord Polski Masters w kat. G /55-59/" eventid="1391" points="292" swimtime="00:03:10.13" resultid="4085" heatid="7093" lane="3" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:24.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat G /55-59/" eventid="1528" points="306" swimtime="00:01:35.64" resultid="4086" heatid="7153" lane="2" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="4087">
              <RESULTS>
                <RESULT eventid="1134" points="197" swimtime="00:00:41.25" resultid="4088" heatid="6991" lane="2" entrytime="00:00:41.50" />
                <RESULT eventid="1316" points="164" swimtime="00:01:34.77" resultid="4089" heatid="7068" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="141" swimtime="00:03:34.61" resultid="4090" heatid="7142" lane="3" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                    <SPLIT distance="100" swimtime="00:01:47.85" />
                    <SPLIT distance="150" swimtime="00:02:44.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="4091">
              <RESULTS>
                <RESULT eventid="1224" points="130" swimtime="00:03:40.08" resultid="4092" heatid="7026" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:45.32" />
                    <SPLIT distance="150" swimtime="00:02:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="283" swimtime="00:00:40.61" resultid="4093" heatid="7057" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1406" points="224" swimtime="00:03:07.60" resultid="4094" heatid="7098" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:24.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="205" swimtime="00:03:09.68" resultid="4095" heatid="7143" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:32.65" />
                    <SPLIT distance="150" swimtime="00:02:21.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Ryszard" gender="M" lastname="Nowak" nation="POL" athleteid="4096">
              <RESULTS>
                <RESULT eventid="1134" points="246" swimtime="00:00:38.33" resultid="4097" heatid="6993" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="1316" points="218" swimtime="00:01:26.27" resultid="4098" heatid="7069" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="227" swimtime="00:00:34.27" resultid="4099" heatid="7125" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1498" status="DNS" swimtime="00:00:00.00" resultid="4100" heatid="7143" lane="6" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="4101">
              <RESULTS>
                <RESULT eventid="1104" points="351" swimtime="00:03:00.43" resultid="4102" heatid="6979" lane="1" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:26.03" />
                    <SPLIT distance="150" swimtime="00:02:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="419" swimtime="00:00:35.63" resultid="4103" heatid="7058" lane="3" entrytime="00:00:36.50" />
                <RESULT eventid="1376" points="331" swimtime="00:02:27.38" resultid="4104" heatid="7087" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="385" swimtime="00:01:20.46" resultid="4105" heatid="7161" lane="1" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="229" swimtime="00:02:32.53" resultid="4106" heatid="7000" lane="0" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                    <SPLIT distance="150" swimtime="00:01:59.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4096" number="1" />
                    <RELAYPOSITION athleteid="4091" number="2" />
                    <RELAYPOSITION athleteid="4101" number="3" />
                    <RELAYPOSITION athleteid="4087" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="GRKOZ" name="Grot Koziegłowy" nation="POL" region="WIE">
          <CONTACT name="Ewa Szała" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="4111">
              <RESULTS>
                <RESULT eventid="1119" points="293" swimtime="00:00:40.73" resultid="4112" heatid="6984" lane="4" entrytime="00:00:41.20" />
                <RESULT eventid="1179" points="293" swimtime="00:01:18.31" resultid="4113" heatid="7005" lane="3" entrytime="00:01:22.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="303" swimtime="00:01:26.49" resultid="4114" heatid="7064" lane="1" entrytime="00:01:33.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="278" swimtime="00:02:53.08" resultid="4115" heatid="7080" lane="2" entrytime="00:02:48.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="150" swimtime="00:02:09.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="294" swimtime="00:03:07.57" resultid="4116" heatid="7138" lane="4" entrytime="00:03:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="150" swimtime="00:02:20.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="273" swimtime="00:06:08.21" resultid="4117" heatid="7166" lane="3" entrytime="00:06:09.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:13.05" />
                    <SPLIT distance="200" swimtime="00:03:01.48" />
                    <SPLIT distance="250" swimtime="00:03:49.47" />
                    <SPLIT distance="300" swimtime="00:04:37.13" />
                    <SPLIT distance="350" swimtime="00:05:24.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" name="Steef Wrocław" nation="POL">
          <CONTACT name="Skrzypek Stefan" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="4119">
              <RESULTS>
                <RESULT eventid="1224" points="153" swimtime="00:03:28.36" resultid="4120" heatid="7026" lane="4" entrytime="00:03:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                    <SPLIT distance="150" swimtime="00:02:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="238" swimtime="00:02:44.59" resultid="4121" heatid="7086" lane="1" entrytime="00:02:38.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="150" swimtime="00:02:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="145" swimtime="00:01:34.64" resultid="4122" heatid="7108" lane="1" entrytime="00:01:25.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="252" swimtime="00:05:48.27" resultid="4123" heatid="7170" lane="5" entrytime="00:05:44.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:06.92" />
                    <SPLIT distance="200" swimtime="00:02:52.25" />
                    <SPLIT distance="250" swimtime="00:03:37.07" />
                    <SPLIT distance="300" swimtime="00:04:22.26" />
                    <SPLIT distance="350" swimtime="00:05:05.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMSZC" name="Smt Szczecin" nation="POL" region="ZAC">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Kamila" gender="F" lastname="Wojdak" nation="POL" athleteid="4141">
              <RESULTS>
                <RESULT eventid="1453" points="534" swimtime="00:00:29.24" resultid="7618" heatid="7113" lane="6" />
                <RESULT eventid="1058" points="560" swimtime="00:02:49.96" resultid="4142" heatid="6973" lane="4" entrytime="00:02:44.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:21.84" />
                    <SPLIT distance="150" swimtime="00:02:05.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="544" swimtime="00:00:36.49" resultid="4143" heatid="7051" lane="4" entrytime="00:00:35.17" />
                <RESULT eventid="1391" points="523" swimtime="00:02:36.48" resultid="4144" heatid="7094" lane="5" entrytime="00:02:36.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:59.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" status="DNS" swimtime="00:00:00.00" resultid="4145" heatid="7154" lane="4" entrytime="00:01:16.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Michał" gender="M" lastname="Zaremba" nation="POL" athleteid="4146">
              <RESULTS>
                <RESULT eventid="1406" points="349" swimtime="00:02:41.83" resultid="4147" heatid="7103" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                    <SPLIT distance="150" swimtime="00:02:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M-9 - Niejednoczesne dotknięcie ściany w czasie wykonywania  nawrotu" eventid="1438" status="DSQ" swimtime="00:01:11.22" resultid="4148" heatid="7110" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Piotr" gender="M" lastname="Zaremba" nation="POL" athleteid="4149">
              <RESULTS>
                <RESULT eventid="1406" points="428" swimtime="00:02:31.20" resultid="4150" heatid="7102" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="438" swimtime="00:01:05.58" resultid="4151" heatid="7110" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Rafał" gender="M" lastname="Lisiecki" nation="POL" athleteid="4152">
              <RESULTS>
                <RESULT eventid="1134" points="384" swimtime="00:00:33.06" resultid="4153" heatid="6997" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1316" points="370" swimtime="00:01:12.32" resultid="4154" heatid="7071" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="409" swimtime="00:00:28.15" resultid="4155" heatid="7131" lane="3" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIPOZ" name="Wielkopolski Klub Bałtycki - Poznań" nation="POL" region="WIE">
          <CONTACT name="q" />
          <ATHLETES>
            <ATHLETE birthdate="1946-01-01" firstname="Teresa" gender="F" lastname="Zarzeczańska-Różańska" nation="POL" athleteid="4157">
              <RESULTS>
                <RESULT eventid="1058" points="144" swimtime="00:04:27.01" resultid="4158" heatid="6971" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                    <SPLIT distance="100" swimtime="00:02:08.53" />
                    <SPLIT distance="150" swimtime="00:03:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="188" swimtime="00:00:51.95" resultid="4159" heatid="7049" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1558" points="78" swimtime="00:09:19.45" resultid="4160" heatid="7164" lane="7" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.24" />
                    <SPLIT distance="100" swimtime="00:02:02.27" />
                    <SPLIT distance="150" swimtime="00:03:11.59" />
                    <SPLIT distance="200" swimtime="00:04:23.65" />
                    <SPLIT distance="250" swimtime="00:05:38.37" />
                    <SPLIT distance="300" swimtime="00:06:51.83" />
                    <SPLIT distance="350" swimtime="00:08:07.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIRZE" name="Rzeszów niezrzeszony" nation="POL" region="PDK">
          <CONTACT city="Rzeszów" email="wieslawcieklinski@wp.pl" name="Ciekliński" phone="602682904" state="PODKA" street="Jagiellońska 7/3" zip="35-025" />
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="4167">
              <RESULTS>
                <RESULT eventid="1194" points="277" swimtime="00:01:11.92" resultid="4168" heatid="7015" lane="0" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="186" swimtime="00:00:39.23" resultid="4169" heatid="7038" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1376" points="212" swimtime="00:02:51.05" resultid="4170" heatid="7085" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="301" swimtime="00:00:31.20" resultid="4171" heatid="7127" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1573" points="200" swimtime="00:06:16.09" resultid="4172" heatid="7170" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:14.69" />
                    <SPLIT distance="200" swimtime="00:03:04.19" />
                    <SPLIT distance="250" swimtime="00:03:54.06" />
                    <SPLIT distance="300" swimtime="00:04:43.74" />
                    <SPLIT distance="350" swimtime="00:05:32.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLSTR" name="Olimpic Strawczynek" nation="POL" region="SWI">
          <CONTACT city="Kielce" email="lipskakatarzyna@wp.pl" fax="-" name="Janusz Lipski" phone="600154761" state="ŚWIĘT" street="Słowackiego 11/1" zip="25-365" />
          <ATHLETES>
            <ATHLETE birthdate="1952-01-27" firstname="Janusz" gender="M" lastname="Lipski" nation="POL" athleteid="4174">
              <RESULTS>
                <RESULT eventid="1194" points="239" swimtime="00:01:15.56" resultid="4175" heatid="7014" lane="5" entrytime="00:01:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4176" heatid="7039" lane="0" entrytime="00:00:36.20" />
                <RESULT eventid="1376" status="DNS" swimtime="00:00:00.00" resultid="4177" heatid="7086" lane="7" entrytime="00:02:38.40" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="4178" heatid="7125" lane="9" entrytime="00:00:34.10" />
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="4179" heatid="7170" lane="4" entrytime="00:05:42.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CIPOZ" name="CityZen Poznań" nation="POL" region="WIE">
          <CONTACT email="uks@ukscityzen.pl" internet="www.ukscityzen.pl" name="Roszak" />
          <ATHLETES>
            <ATHLETE birthdate="1985-01-01" firstname="Tadeusz" gender="M" lastname="Gołembiewski" nation="POL" athleteid="4181">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="4182" heatid="7022" lane="1" entrytime="00:00:57.00" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="4183" heatid="7028" lane="3" entrytime="00:02:44.00" />
                <RESULT eventid="1256" points="452" swimtime="00:00:29.22" resultid="4184" heatid="7045" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1376" points="446" swimtime="00:02:13.42" resultid="4185" heatid="7090" lane="0" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.45" />
                    <SPLIT distance="150" swimtime="00:01:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="365" swimtime="00:01:09.69" resultid="4186" heatid="7112" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="399" swimtime="00:04:58.89" resultid="4187" heatid="7172" lane="0" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:49.21" />
                    <SPLIT distance="200" swimtime="00:02:27.65" />
                    <SPLIT distance="250" swimtime="00:03:06.26" />
                    <SPLIT distance="300" swimtime="00:03:44.99" />
                    <SPLIT distance="350" swimtime="00:04:23.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKAT" name="UKS Wodnik 29 Katowice" nation="POL" region="SLA">
          <CONTACT city="Katowice" name="Mrozińska Bożena" phone="502013302" state="ŚLĄSK" street="Barbary 14/9" />
          <ATHLETES>
            <ATHLETE birthdate="1932-01-01" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="4189">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat.L /80-84/" eventid="1119" points="86" swimtime="00:01:01.14" resultid="4190" heatid="6982" lane="2" entrytime="00:01:01.80" />
                <RESULT comment="Rekord Polski Masters w kat. L /80-84/" eventid="1301" points="55" swimtime="00:02:32.10" resultid="4191" heatid="7063" lane="8" entrytime="00:02:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="53" swimtime="00:01:02.88" resultid="4192" heatid="7114" lane="3" entrytime="00:01:00.00" />
                <RESULT comment="Rekord Polski Masters w kat L /80-84/" eventid="1558" points="45" swimtime="00:11:11.29" resultid="4193" heatid="7164" lane="1" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.73" />
                    <SPLIT distance="100" swimtime="00:02:32.50" />
                    <SPLIT distance="150" swimtime="00:03:57.74" />
                    <SPLIT distance="200" swimtime="00:05:25.57" />
                    <SPLIT distance="250" swimtime="00:06:52.45" />
                    <SPLIT distance="300" swimtime="00:08:19.42" />
                    <SPLIT distance="350" swimtime="00:09:45.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Maria" gender="F" lastname="ŚMIGLEWSKA" nation="POL" athleteid="4194">
              <RESULTS>
                <RESULT eventid="1058" points="36" swimtime="00:07:03.35" resultid="4195" heatid="6970" lane="6" entrytime="00:06:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.95" />
                    <SPLIT distance="100" swimtime="00:03:22.08" />
                    <SPLIT distance="150" swimtime="00:05:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="39" swimtime="00:01:19.16" resultid="4196" heatid="6983" lane="0" />
                <RESULT eventid="1271" points="31" swimtime="00:01:34.74" resultid="4197" heatid="7048" lane="9" entrytime="00:01:35.00" />
                <RESULT eventid="1528" points="30" swimtime="00:03:25.52" resultid="4198" heatid="7151" lane="9" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:42.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Marcin" gender="M" lastname="SZCZYPIŃSKI" nation="POL" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1194" points="597" swimtime="00:00:55.69" resultid="4200" heatid="7022" lane="2" entrytime="00:00:56.00" />
                <RESULT eventid="1256" points="542" swimtime="00:00:27.50" resultid="4201" heatid="7045" lane="8" entrytime="00:00:27.80" />
                <RESULT eventid="1376" points="521" swimtime="00:02:06.74" resultid="4202" heatid="7090" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="547" swimtime="00:01:00.89" resultid="4203" heatid="7111" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. A /25-29/" eventid="1573" points="533" swimtime="00:04:31.32" resultid="4204" heatid="7174" lane="1" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:02.83" />
                    <SPLIT distance="150" swimtime="00:01:36.78" />
                    <SPLIT distance="200" swimtime="00:02:11.52" />
                    <SPLIT distance="250" swimtime="00:02:46.04" />
                    <SPLIT distance="300" swimtime="00:03:21.22" />
                    <SPLIT distance="350" swimtime="00:03:56.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Michał" gender="M" lastname="Spławiński" nation="POL" athleteid="4205">
              <RESULTS>
                <RESULT eventid="1104" points="348" swimtime="00:03:00.96" resultid="4206" heatid="6979" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:29.12" />
                    <SPLIT distance="150" swimtime="00:02:17.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="426" swimtime="00:00:31.94" resultid="4207" heatid="6997" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1256" points="558" swimtime="00:00:27.23" resultid="4208" heatid="7045" lane="3" entrytime="00:00:27.36" />
                <RESULT eventid="1286" points="594" swimtime="00:00:31.72" resultid="4209" heatid="7061" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1468" points="503" swimtime="00:00:26.28" resultid="4210" heatid="7136" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1543" points="515" swimtime="00:01:13.06" resultid="4211" heatid="7160" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-01-01" firstname="Wiktoria" gender="F" lastname="Skrzesińska - Gabryś" nation="POL" athleteid="4212">
              <RESULTS>
                <RESULT eventid="1119" points="31" swimtime="00:01:25.52" resultid="4213" heatid="6982" lane="9" entrytime="00:01:24.00" />
                <RESULT eventid="1271" points="43" swimtime="00:01:24.64" resultid="4214" heatid="7048" lane="0" entrytime="00:01:24.00" />
                <RESULT eventid="1453" points="35" swimtime="00:01:12.46" resultid="4215" heatid="7114" lane="2" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4216">
              <RESULTS>
                <RESULT eventid="1134" points="335" swimtime="00:00:34.60" resultid="4217" heatid="6994" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1194" points="414" swimtime="00:01:02.94" resultid="4218" heatid="7019" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="293" swimtime="00:01:18.14" resultid="4219" heatid="7070" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="340" swimtime="00:02:26.07" resultid="4220" heatid="7088" lane="0" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="248" swimtime="00:02:58.01" resultid="4221" heatid="7144" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                    <SPLIT distance="150" swimtime="00:02:13.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="330" swimtime="00:05:18.21" resultid="4222" heatid="7172" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                    <SPLIT distance="200" swimtime="00:02:33.70" />
                    <SPLIT distance="250" swimtime="00:03:16.05" />
                    <SPLIT distance="300" swimtime="00:03:58.03" />
                    <SPLIT distance="350" swimtime="00:04:39.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Edyta" gender="F" lastname="Mróz" nation="POL" athleteid="4223">
              <RESULTS>
                <RESULT eventid="1119" points="337" swimtime="00:00:38.86" resultid="4224" heatid="6985" lane="4" entrytime="00:00:38.40" />
                <RESULT eventid="1301" points="354" swimtime="00:01:22.09" resultid="4225" heatid="7065" lane="8" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="344" swimtime="00:02:41.19" resultid="4226" heatid="7080" lane="4" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                    <SPLIT distance="150" swimtime="00:02:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1483" points="347" swimtime="00:02:57.56" resultid="4227" heatid="7139" lane="3" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:02:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1558" points="349" swimtime="00:05:39.55" resultid="4228" heatid="7167" lane="9" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:04.69" />
                    <SPLIT distance="200" swimtime="00:02:48.15" />
                    <SPLIT distance="250" swimtime="00:03:32.08" />
                    <SPLIT distance="300" swimtime="00:04:15.71" />
                    <SPLIT distance="350" swimtime="00:04:59.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="4229">
              <RESULTS>
                <RESULT eventid="1194" points="561" swimtime="00:00:56.86" resultid="4230" heatid="7021" lane="3" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="539" swimtime="00:00:27.56" resultid="4231" heatid="7045" lane="2" entrytime="00:00:27.40" />
                <RESULT eventid="1376" points="472" swimtime="00:02:10.96" resultid="4232" heatid="7089" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="100" swimtime="00:01:04.21" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="489" swimtime="00:00:26.54" resultid="4233" heatid="7136" lane="1" entrytime="00:00:25.55" />
                <RESULT eventid="1573" points="433" swimtime="00:04:50.73" resultid="4234" heatid="7172" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:46.47" />
                    <SPLIT distance="200" swimtime="00:02:23.69" />
                    <SPLIT distance="250" swimtime="00:03:01.09" />
                    <SPLIT distance="300" swimtime="00:03:38.81" />
                    <SPLIT distance="350" swimtime="00:04:16.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4235">
              <RESULTS>
                <RESULT eventid="1104" points="287" swimtime="00:03:12.82" resultid="4236" heatid="6978" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:31.01" />
                    <SPLIT distance="150" swimtime="00:02:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="276" swimtime="00:01:12.04" resultid="4237" heatid="7015" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="432" swimtime="00:00:35.27" resultid="4238" heatid="7058" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1376" points="228" swimtime="00:02:46.73" resultid="4239" heatid="7085" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="352" swimtime="00:01:22.96" resultid="4240" heatid="7160" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="4241">
              <RESULTS>
                <RESULT eventid="1194" points="224" swimtime="00:01:17.18" resultid="4242" heatid="7009" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="123" swimtime="00:03:44.03" resultid="4243" heatid="7026" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:44.28" />
                    <SPLIT distance="150" swimtime="00:02:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="293" swimtime="00:00:33.77" resultid="4244" heatid="7041" lane="9" entrytime="00:00:33.50" />
                <RESULT eventid="1406" points="177" swimtime="00:03:22.85" resultid="4245" heatid="7097" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:29.20" />
                    <SPLIT distance="150" swimtime="00:02:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="182" swimtime="00:01:27.79" resultid="4246" heatid="7108" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="253" swimtime="00:00:33.03" resultid="4247" heatid="7122" lane="9" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Tomasz" gender="M" lastname="Kozioł" nation="POL" athleteid="4248">
              <RESULTS>
                <RESULT eventid="1104" points="369" swimtime="00:02:57.34" resultid="4249" heatid="6978" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:25.23" />
                    <SPLIT distance="150" swimtime="00:02:11.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="449" swimtime="00:01:01.24" resultid="4250" heatid="7017" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="388" swimtime="00:02:19.73" resultid="4251" heatid="7087" lane="4" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                    <SPLIT distance="150" swimtime="00:01:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="403" swimtime="00:02:34.25" resultid="4252" heatid="7101" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:58.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4253" heatid="7158" lane="3" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Tomasz" gender="M" lastname="Gruszka" nation="POL" athleteid="4254">
              <RESULTS>
                <RESULT eventid="1134" points="427" swimtime="00:00:31.91" resultid="4255" heatid="6997" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1194" points="445" swimtime="00:01:01.44" resultid="4256" heatid="7021" lane="8" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="385" swimtime="00:01:11.34" resultid="4257" heatid="7072" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="440" swimtime="00:00:27.48" resultid="4258" heatid="7136" lane="9" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Michał" gender="M" lastname="Gorazdowski" nation="POL" athleteid="4259">
              <RESULTS>
                <RESULT eventid="1194" points="295" swimtime="00:01:10.42" resultid="4260" heatid="7016" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="240" swimtime="00:00:42.91" resultid="4261" heatid="7056" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1468" points="325" swimtime="00:00:30.40" resultid="4262" heatid="7131" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1543" points="194" swimtime="00:01:41.04" resultid="4263" heatid="7160" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="4264">
              <RESULTS>
                <RESULT eventid="1179" points="405" swimtime="00:01:10.34" resultid="4265" heatid="7008" lane="2" entrytime="00:01:06.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="478" swimtime="00:00:32.05" resultid="4266" heatid="7034" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1391" points="357" swimtime="00:02:57.72" resultid="4267" heatid="7094" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:24.20" />
                    <SPLIT distance="150" swimtime="00:02:16.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="477" swimtime="00:00:30.35" resultid="4268" heatid="7120" lane="3" entrytime="00:00:28.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. B /120-159/" eventid="1164" points="504" swimtime="00:01:57.36" resultid="4269" heatid="7001" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:32.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4216" number="1" />
                    <RELAYPOSITION athleteid="4205" number="2" />
                    <RELAYPOSITION athleteid="4229" number="3" />
                    <RELAYPOSITION athleteid="4199" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters w kat. B /120-159/" eventid="1346" points="521" swimtime="00:01:45.42" resultid="4352" heatid="7075" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:00:54.61" />
                    <SPLIT distance="150" swimtime="00:01:20.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4216" number="1" />
                    <RELAYPOSITION athleteid="4205" number="2" />
                    <RELAYPOSITION athleteid="4229" number="3" />
                    <RELAYPOSITION athleteid="4199" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat B /120-159/" eventid="1513" points="397" swimtime="00:02:07.11" resultid="4270" heatid="7149" lane="4" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="150" swimtime="00:01:37.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4223" number="1" />
                    <RELAYPOSITION athleteid="4205" number="2" />
                    <RELAYPOSITION athleteid="4229" number="3" />
                    <RELAYPOSITION athleteid="4264" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TORPE" name="Torpedos" nation="LTU">
          <CONTACT city="MARIJAMPOLE" email="vilmantasenator@gmail.com" internet="www.torpedos.puslapiai.lt" name="VILMANTAS KRASAUSKAS" phone="+370 687 46068" street="JUKNEVICIAUS 78-10" zip="68198" />
          <ATHLETES>
            <ATHLETE birthdate="1964-07-31" firstname="VILMANTAS" gender="M" lastname="KRASAUSKAS" nation="LTU" license="Marijampole" athleteid="4284">
              <RESULTS>
                <RESULT eventid="1194" points="371" swimtime="00:01:05.23" resultid="4285" heatid="7019" lane="1" entrytime="00:01:02.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="374" swimtime="00:02:21.47" resultid="4286" heatid="7088" lane="8" entrytime="00:02:20.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="350" swimtime="00:00:29.65" resultid="4287" heatid="7129" lane="5" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="1573" points="389" swimtime="00:05:01.37" resultid="4288" heatid="7173" lane="0" entrytime="00:04:58.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                    <SPLIT distance="200" swimtime="00:02:30.95" />
                    <SPLIT distance="250" swimtime="00:03:08.48" />
                    <SPLIT distance="300" swimtime="00:03:46.67" />
                    <SPLIT distance="350" swimtime="00:04:24.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-04" firstname="JURATE" gender="F" lastname="PRANCKEVICIENE" nation="LTU" license="Marijampole" athleteid="4289">
              <RESULTS>
                <RESULT eventid="1179" points="343" swimtime="00:01:14.32" resultid="4290" heatid="7007" lane="8" entrytime="00:01:14.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="361" swimtime="00:00:33.32" resultid="4291" heatid="7119" lane="7" entrytime="00:00:32.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-03-14" firstname="STASYS" gender="M" lastname="GRIGAS" nation="LTU" license="Marijampole" athleteid="4292">
              <RESULTS>
                <RESULT eventid="1104" points="63" swimtime="00:05:18.37" resultid="4293" heatid="6974" lane="1" entrytime="00:05:08.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.83" />
                    <SPLIT distance="100" swimtime="00:02:23.75" />
                    <SPLIT distance="150" swimtime="00:03:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="49" swimtime="00:01:05.59" resultid="4294" heatid="6987" lane="3" entrytime="00:01:10.26" entrycourse="SCM" />
                <RESULT eventid="1286" points="105" swimtime="00:00:56.40" resultid="4295" heatid="7053" lane="8" entrytime="00:00:55.74" entrycourse="LCM" />
                <RESULT eventid="1316" points="48" swimtime="00:02:22.40" resultid="4296" heatid="7067" lane="9" entrytime="00:02:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="47" swimtime="00:05:09.77" resultid="4297" heatid="7140" lane="4" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.69" />
                    <SPLIT distance="100" swimtime="00:02:28.91" />
                    <SPLIT distance="150" swimtime="00:03:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="63" swimtime="00:02:26.59" resultid="4298" heatid="7155" lane="5" entrytime="00:02:12.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQWRO" name="Aquapark Wrocław" nation="POL" region="DOL">
          <CONTACT name="Kujat" street="Borowska 99" />
          <ATHLETES>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="Stasiaczek" nation="POL" athleteid="4300">
              <RESULTS>
                <RESULT eventid="1104" points="451" swimtime="00:02:45.94" resultid="4301" heatid="6980" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="522" swimtime="00:00:33.11" resultid="4302" heatid="7061" lane="7" entrytime="00:00:31.99" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="4303" heatid="7102" lane="2" entrytime="00:02:35.00" />
                <RESULT eventid="1543" points="493" swimtime="00:01:14.12" resultid="4304" heatid="7163" lane="2" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-09" firstname="Michał" gender="M" lastname="Witkowski" nation="POL" athleteid="4305">
              <RESULTS>
                <RESULT eventid="1194" points="541" swimtime="00:00:57.56" resultid="4306" heatid="7022" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1256" points="502" swimtime="00:00:28.21" resultid="4307" heatid="7046" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="1468" points="515" swimtime="00:00:26.08" resultid="4308" heatid="7136" lane="4" entrytime="00:00:23.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-01" firstname="Tomasz" gender="M" lastname="Cimicki" nation="POL" athleteid="4309">
              <RESULTS>
                <RESULT eventid="1104" points="343" swimtime="00:03:01.73" resultid="4310" heatid="6980" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                    <SPLIT distance="150" swimtime="00:02:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="419" swimtime="00:00:35.62" resultid="4311" heatid="7060" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1543" points="377" swimtime="00:01:21.04" resultid="4312" heatid="7163" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-09" firstname="Paweł" gender="M" lastname="Handke" nation="POL" athleteid="4313">
              <RESULTS>
                <RESULT eventid="1104" points="436" swimtime="00:02:47.84" resultid="4314" heatid="6980" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:04.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="504" swimtime="00:00:58.94" resultid="4315" heatid="7021" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="4316" heatid="7061" lane="0" entrytime="00:00:32.57" />
                <RESULT eventid="1376" points="470" swimtime="00:02:11.18" resultid="4317" heatid="7090" lane="5" entrytime="00:02:03.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="430" swimtime="00:00:27.69" resultid="4318" heatid="7135" lane="9" entrytime="00:00:26.42" />
                <RESULT eventid="1543" points="416" swimtime="00:01:18.44" resultid="4319" heatid="7163" lane="9" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-24" firstname="Krystian" gender="M" lastname="Młyński" nation="POL" athleteid="4320">
              <RESULTS>
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="4321" heatid="6997" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1468" points="407" swimtime="00:00:28.20" resultid="4322" heatid="7133" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1498" points="247" swimtime="00:02:58.27" resultid="4323" heatid="7145" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:23.73" />
                    <SPLIT distance="150" swimtime="00:02:09.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-29" firstname="Łukasz" gender="M" lastname="Lesiewicz" nation="POL" athleteid="4324">
              <RESULTS>
                <RESULT eventid="1134" points="396" swimtime="00:00:32.71" resultid="4325" heatid="6994" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1316" points="382" swimtime="00:01:11.58" resultid="4326" heatid="7070" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="420" swimtime="00:00:27.90" resultid="4327" heatid="7129" lane="1" entrytime="00:00:30.00" />
                <RESULT comment="G-1 - Nieutrzymanie pozycji na plecach " eventid="1498" status="DSQ" swimtime="00:02:44.61" resultid="4328" heatid="7145" lane="9" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                    <SPLIT distance="150" swimtime="00:02:00.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="4329">
              <RESULTS>
                <RESULT eventid="1104" points="436" swimtime="00:02:47.89" resultid="4330" heatid="6980" lane="4" entrytime="00:02:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:03.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="536" swimtime="00:00:32.83" resultid="4331" heatid="7061" lane="1" entrytime="00:00:31.99" />
                <RESULT eventid="1543" points="474" swimtime="00:01:15.09" resultid="4332" heatid="7163" lane="6" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="4333" heatid="7001" lane="1" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4320" number="1" />
                    <RELAYPOSITION athleteid="4300" number="2" />
                    <RELAYPOSITION athleteid="4305" number="3" />
                    <RELAYPOSITION athleteid="4313" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="4334" heatid="7076" lane="9" entrytime="00:01:54.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4313" number="1" />
                    <RELAYPOSITION athleteid="4300" number="2" />
                    <RELAYPOSITION athleteid="4305" number="3" />
                    <RELAYPOSITION athleteid="4309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="433" swimtime="00:02:03.47" resultid="4466" heatid="7001" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:36.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4309" number="1" />
                    <RELAYPOSITION athleteid="4300" number="2" />
                    <RELAYPOSITION athleteid="4305" number="3" />
                    <RELAYPOSITION athleteid="4313" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="447" swimtime="00:01:50.93" resultid="4467" heatid="7075" lane="4" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                    <SPLIT distance="100" swimtime="00:00:54.61" />
                    <SPLIT distance="150" swimtime="00:01:22.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4313" number="1" />
                    <RELAYPOSITION athleteid="4300" number="2" />
                    <RELAYPOSITION athleteid="4305" number="3" />
                    <RELAYPOSITION athleteid="4309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KOOLS" name="Masters Kormoran Olsztyn" nation="POL" region="WAR">
          <CONTACT city="Olsztyn/Łupstych" email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" phone="501372846" state="WARM-" street="Leśna 1" zip="11-041" />
          <ATHLETES>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="4816">
              <RESULTS>
                <RESULT eventid="1058" points="291" swimtime="00:03:31.32" resultid="4817" heatid="6972" lane="5" entrytime="00:03:28.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.80" />
                    <SPLIT distance="100" swimtime="00:01:42.23" />
                    <SPLIT distance="150" swimtime="00:02:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="325" swimtime="00:01:15.72" resultid="4818" heatid="7006" lane="4" entrytime="00:01:15.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="303" swimtime="00:02:48.05" resultid="4819" heatid="7080" lane="3" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="150" swimtime="00:02:05.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1391" points="266" swimtime="00:03:16.05" resultid="4820" heatid="7093" lane="7" entrytime="00:03:15.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:01:34.70" />
                    <SPLIT distance="150" swimtime="00:02:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="314" swimtime="00:00:34.88" resultid="4821" heatid="7118" lane="2" entrytime="00:00:34.50" entrycourse="LCM" />
                <RESULT eventid="1558" points="290" swimtime="00:06:00.93" resultid="4822" heatid="7167" lane="0" entrytime="00:05:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:10.23" />
                    <SPLIT distance="200" swimtime="00:02:56.91" />
                    <SPLIT distance="250" swimtime="00:03:43.45" />
                    <SPLIT distance="300" swimtime="00:04:30.18" />
                    <SPLIT distance="350" swimtime="00:05:16.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-14" firstname="Dariusz" gender="M" lastname="Poziemski" nation="POL" athleteid="4823">
              <RESULTS>
                <RESULT eventid="1134" points="351" swimtime="00:00:34.07" resultid="4824" heatid="6995" lane="4" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="374" swimtime="00:00:31.13" resultid="4825" heatid="7042" lane="8" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1316" points="327" swimtime="00:01:15.39" resultid="4826" heatid="7071" lane="7" entrytime="00:01:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="4827">
              <RESULTS>
                <RESULT eventid="1256" points="377" swimtime="00:00:31.04" resultid="4828" heatid="7043" lane="1" entrytime="00:00:30.21" entrycourse="LCM" />
                <RESULT eventid="1376" points="388" swimtime="00:02:19.83" resultid="4829" heatid="7088" lane="4" entrytime="00:02:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="349" swimtime="00:01:10.70" resultid="4830" heatid="7108" lane="3" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-4 - Przedwczwsny start" eventid="1573" status="DSQ" swimtime="00:04:58.09" resultid="4831" heatid="7172" lane="5" entrytime="00:05:01.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="150" swimtime="00:01:49.72" />
                    <SPLIT distance="200" swimtime="00:02:27.90" />
                    <SPLIT distance="250" swimtime="00:03:06.22" />
                    <SPLIT distance="300" swimtime="00:03:44.30" />
                    <SPLIT distance="350" swimtime="00:04:22.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPIA" name="Mks Piaseczno" nation="POL" region="MAZ">
          <CONTACT city="PIASECZNO" name="ANDRZEJ RUBASZKIEWICZ" />
          <ATHLETES>
            <ATHLETE birthdate="1949-04-10" firstname="ANDRZEJ" gender="M" lastname="RUBASZKIEWICZ" nation="POL" athleteid="4833">
              <RESULTS>
                <RESULT eventid="1134" points="250" swimtime="00:00:38.15" resultid="4834" heatid="6993" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1194" points="342" swimtime="00:01:07.04" resultid="4835" heatid="7017" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="284" swimtime="00:00:34.10" resultid="4836" heatid="7040" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1376" points="256" swimtime="00:02:40.58" resultid="4837" heatid="7085" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="157" swimtime="00:01:32.34" resultid="4838" heatid="7108" lane="5" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="319" swimtime="00:00:30.58" resultid="4839" heatid="7128" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SUPOL" name="Śródmiejski Uczniowski Klub Sportowy" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="suks.polna@gmail.com" internet="www.sukspolna.pl" name="Gapińska Agnieszka" street="Polna 7a" zip="00-625" />
          <ATHLETES>
            <ATHLETE birthdate="1984-12-19" firstname="Agnieszka" gender="F" lastname="Gapińska" nation="POL" athleteid="4841">
              <RESULTS>
                <RESULT eventid="1179" points="330" swimtime="00:01:15.33" resultid="4842" heatid="7007" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="364" swimtime="00:00:35.08" resultid="4843" heatid="7034" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1453" points="381" swimtime="00:00:32.71" resultid="4844" heatid="7118" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-08-12" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="4845">
              <RESULTS>
                <RESULT eventid="1119" points="187" swimtime="00:00:47.28" resultid="4846" heatid="6983" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1453" points="214" swimtime="00:00:39.63" resultid="4847" heatid="7116" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-21" firstname="Elżbieta" gender="F" lastname="Mzyk" nation="POL" athleteid="4848">
              <RESULTS>
                <RESULT eventid="1179" points="188" swimtime="00:01:30.82" resultid="4849" heatid="7004" lane="3" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="217" swimtime="00:00:41.71" resultid="4850" heatid="7032" lane="7" entrytime="00:00:42.00" />
                <RESULT comment="O-4 - Przedwczwsny start" eventid="1391" status="DSQ" swimtime="00:03:49.16" resultid="4851" heatid="7092" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:56.33" />
                    <SPLIT distance="150" swimtime="00:02:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" points="156" swimtime="00:01:43.98" resultid="4852" heatid="7105" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-02" firstname="Piotr" gender="M" lastname="Przybylski" nation="POL" athleteid="4853">
              <RESULTS>
                <RESULT eventid="1224" points="194" swimtime="00:03:12.54" resultid="4854" heatid="7027" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:28.61" />
                    <SPLIT distance="150" swimtime="00:02:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="370" swimtime="00:00:29.12" resultid="4855" heatid="7129" lane="0" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-12-24" firstname="Justyna" gender="F" lastname="Tarnowska" nation="POL" athleteid="4856">
              <RESULTS>
                <RESULT eventid="1558" points="245" swimtime="00:06:21.94" resultid="4857" heatid="7166" lane="2" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:16.38" />
                    <SPLIT distance="200" swimtime="00:03:05.65" />
                    <SPLIT distance="250" swimtime="00:03:55.72" />
                    <SPLIT distance="300" swimtime="00:04:46.14" />
                    <SPLIT distance="350" swimtime="00:05:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="4858">
              <RESULTS>
                <RESULT eventid="1134" points="273" swimtime="00:00:37.05" resultid="4859" heatid="6993" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1286" points="380" swimtime="00:00:36.80" resultid="4860" heatid="7057" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1468" points="399" swimtime="00:00:28.38" resultid="4861" heatid="7131" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1543" points="318" swimtime="00:01:25.75" resultid="4862" heatid="7160" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="295" swimtime="00:02:25.26" resultid="4864" heatid="7073" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:47.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4841" number="1" />
                    <RELAYPOSITION athleteid="4856" number="2" />
                    <RELAYPOSITION athleteid="4845" number="3" />
                    <RELAYPOSITION athleteid="4848" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1149" points="279" swimtime="00:02:42.29" resultid="4865" heatid="6998" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:33.26" />
                    <SPLIT distance="150" swimtime="00:02:07.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4845" number="1" />
                    <RELAYPOSITION athleteid="4848" number="2" />
                    <RELAYPOSITION athleteid="4841" number="3" />
                    <RELAYPOSITION athleteid="4856" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1513" points="253" swimtime="00:02:27.69" resultid="4863" heatid="7148" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:01:59.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4845" number="1" />
                    <RELAYPOSITION athleteid="4858" number="2" />
                    <RELAYPOSITION athleteid="4841" number="3" />
                    <RELAYPOSITION athleteid="4853" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KAPRU" name="UKS Kapry-Armexim Pruszków" nation="POL" region="MAZ">
          <CONTACT name="borkowski" />
          <ATHLETES>
            <ATHLETE birthdate="1987-09-16" firstname="Mariusz" gender="M" lastname="Winogrodzki" nation="POL" athleteid="4873">
              <RESULTS>
                <RESULT eventid="1256" points="574" swimtime="00:00:26.98" resultid="4874" heatid="7046" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="1286" points="679" swimtime="00:00:30.33" resultid="4875" heatid="7061" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1543" points="628" swimtime="00:01:08.38" resultid="4876" heatid="7163" lane="4" entrytime="00:01:06.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPFIG" name="WOPR Warszawa SPORT-Figielski" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="sport-figielski@o2.pl" fax="224032788" internet="www.sport-figielski.pl" name="Grzegorz Figielski" phone="501294477" state="MAZ" street="Sarmacka 21 m. 41" zip="02-594" />
          <ATHLETES>
            <ATHLETE birthdate="1965-02-05" firstname="Agata" gender="F" lastname="Figielska" nation="POL" athleteid="4878">
              <RESULTS>
                <RESULT eventid="1271" points="111" swimtime="00:01:01.99" resultid="4879" heatid="7048" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1528" points="92" swimtime="00:02:22.49" resultid="4880" heatid="7151" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-12-27" firstname="Grzegorz" gender="M" lastname="Figielski" nation="POL" athleteid="4881">
              <RESULTS>
                <RESULT eventid="1376" points="171" swimtime="00:03:03.64" resultid="4882" heatid="7084" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:25.62" />
                    <SPLIT distance="150" swimtime="00:02:14.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="123" swimtime="00:03:48.81" resultid="4883" heatid="7096" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.91" />
                    <SPLIT distance="100" swimtime="00:01:55.27" />
                    <SPLIT distance="150" swimtime="00:03:01.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-25" firstname="Fabian" gender="M" lastname="Filipiak" nation="POL" athleteid="4884">
              <RESULTS>
                <RESULT eventid="1104" points="87" swimtime="00:04:46.86" resultid="4885" heatid="6974" lane="7" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.35" />
                    <SPLIT distance="100" swimtime="00:02:18.43" />
                    <SPLIT distance="150" swimtime="00:03:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="51" swimtime="00:04:59.56" resultid="4886" heatid="7025" lane="6" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.47" />
                    <SPLIT distance="100" swimtime="00:02:18.52" />
                    <SPLIT distance="150" swimtime="00:03:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="68" swimtime="00:02:06.76" resultid="4887" heatid="7067" lane="1" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="83" swimtime="00:04:21.07" resultid="4888" heatid="7095" lane="4" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.90" />
                    <SPLIT distance="100" swimtime="00:02:08.78" />
                    <SPLIT distance="150" swimtime="00:03:24.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="47" swimtime="00:02:17.28" resultid="4889" heatid="7106" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="83" swimtime="00:04:16.32" resultid="4890" heatid="7141" lane="6" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.30" />
                    <SPLIT distance="100" swimtime="00:02:05.44" />
                    <SPLIT distance="150" swimtime="00:03:12.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-19" firstname="Andrzej" gender="M" lastname="Gryboś" nation="POL" athleteid="4891">
              <RESULTS>
                <RESULT eventid="1376" points="203" swimtime="00:02:53.28" resultid="4892" heatid="7083" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:02:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" status="DNS" swimtime="00:00:00.00" resultid="4893" heatid="7169" lane="6" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-03-13" firstname="Alina" gender="F" lastname="Kraśniewska" nation="POL" athleteid="4894">
              <RESULTS>
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="4895" heatid="7002" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="4896" heatid="7030" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="1391" status="DNS" swimtime="00:00:00.00" resultid="4897" heatid="7091" lane="6" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:05:10.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1422" status="DNS" swimtime="00:00:00.00" resultid="4898" heatid="7104" lane="0" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="4899" heatid="7114" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-09-01" firstname="Maja" gender="F" lastname="Lipniacka" nation="POL" athleteid="4900">
              <RESULTS>
                <RESULT eventid="1119" points="14" swimtime="00:01:51.32" resultid="4901" heatid="6981" lane="4" entrytime="00:01:50.00" />
                <RESULT eventid="1301" points="13" swimtime="00:04:04.22" resultid="4902" heatid="7062" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:56.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1528" points="13" swimtime="00:04:31.93" resultid="4903" heatid="7150" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:15.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-08-25" firstname="Stanisława" gender="F" lastname="Połczyńska" nation="POL" athleteid="4904">
              <RESULTS>
                <RESULT eventid="1271" points="4" swimtime="00:02:58.62" resultid="4905" heatid="7047" lane="4" entrytime="00:03:00.00" />
                <RESULT eventid="1453" status="DNS" swimtime="00:00:00.00" resultid="4906" heatid="7114" lane="0" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-25" firstname="Artur" gender="M" lastname="Ilgner" nation="POL" athleteid="4907">
              <RESULTS>
                <RESULT eventid="1468" points="149" swimtime="00:00:39.39" resultid="7620" heatid="7131" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-29" firstname="Michał" gender="M" lastname="Chojecki" nation="POL" athleteid="4909">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="4910" heatid="7013" lane="6" entrytime="00:01:15.00" />
                <RESULT eventid="1468" points="279" swimtime="00:00:32.00" resultid="4911" heatid="7126" lane="8" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Tadeusz" gender="M" lastname="Vorbrodt" nation="POL" athleteid="4912">
              <RESULTS>
                <RESULT eventid="1134" points="106" swimtime="00:00:50.70" resultid="4913" heatid="6989" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1194" points="144" swimtime="00:01:29.36" resultid="4914" heatid="7011" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="130" swimtime="00:07:13.99" resultid="4915" heatid="7169" lane="0" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:27.59" />
                    <SPLIT distance="200" swimtime="00:03:21.96" />
                    <SPLIT distance="250" swimtime="00:04:18.99" />
                    <SPLIT distance="300" swimtime="00:05:18.10" />
                    <SPLIT distance="350" swimtime="00:06:18.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-04-28" firstname="Joanna" gender="F" lastname="Szczepańska" nation="POL" athleteid="4916">
              <RESULTS>
                <RESULT eventid="1271" points="122" swimtime="00:00:59.93" resultid="4917" heatid="7049" lane="0" entrytime="00:00:53.00" />
                <RESULT eventid="1361" points="66" swimtime="00:04:39.54" resultid="4918" heatid="7077" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.13" />
                    <SPLIT distance="100" swimtime="00:02:09.27" />
                    <SPLIT distance="150" swimtime="00:03:25.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-07-03" firstname="Marcin" gender="M" lastname="Korzycki" nation="POL" athleteid="4919">
              <RESULTS>
                <RESULT eventid="1104" points="185" swimtime="00:03:43.16" resultid="4920" heatid="6976" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                    <SPLIT distance="100" swimtime="00:01:43.08" />
                    <SPLIT distance="150" swimtime="00:02:42.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="231" swimtime="00:00:43.46" resultid="4921" heatid="7056" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="4922" heatid="7158" lane="8" entrytime="00:01:35.00" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="7594" heatid="7121" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-01" firstname="Robert" gender="M" lastname="Zieliński" nation="POL" athleteid="4923">
              <RESULTS>
                <RESULT eventid="1134" points="196" swimtime="00:00:41.34" resultid="4924" heatid="6991" lane="7" entrytime="00:00:41.55" />
                <RESULT eventid="1194" points="224" swimtime="00:01:17.14" resultid="4925" heatid="7013" lane="4" entrytime="00:01:14.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="141" swimtime="00:01:39.72" resultid="4926" heatid="7068" lane="1" entrytime="00:01:35.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="171" swimtime="00:03:03.59" resultid="4927" heatid="7084" lane="3" entrytime="00:02:57.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:02:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="225" swimtime="00:00:34.35" resultid="4928" heatid="7127" lane="1" entrytime="00:00:31.46" />
                <RESULT eventid="1498" points="127" swimtime="00:03:42.27" resultid="4929" heatid="7142" lane="0" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                    <SPLIT distance="100" swimtime="00:01:48.81" />
                    <SPLIT distance="150" swimtime="00:02:47.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-05" firstname="Anna" gender="F" lastname="Zielińska" nation="POL" athleteid="4930">
              <RESULTS>
                <RESULT eventid="1058" points="41" swimtime="00:06:45.63" resultid="4931" heatid="6970" lane="3" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.60" />
                    <SPLIT distance="100" swimtime="00:03:21.58" />
                    <SPLIT distance="150" swimtime="00:05:06.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="34" swimtime="00:02:39.22" resultid="4932" heatid="7002" lane="2" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="35" swimtime="00:01:31.02" resultid="4933" heatid="7048" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1301" points="40" swimtime="00:02:49.55" resultid="4934" heatid="7062" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="32" swimtime="00:01:14.35" resultid="4935" heatid="7114" lane="7" entrytime="00:01:09.00" />
                <RESULT eventid="1528" points="35" swimtime="00:03:15.99" resultid="4936" heatid="7151" lane="1" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-04" firstname="Wiktor" gender="M" lastname="Dębski" nation="BLR" athleteid="4937">
              <RESULTS>
                <RESULT eventid="1286" points="469" swimtime="00:00:34.32" resultid="4938" heatid="7059" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1543" points="398" swimtime="00:01:19.63" resultid="4939" heatid="7161" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-03-07" firstname="Barbara" gender="F" lastname="Czabańska" nation="POL" athleteid="4940">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="4941" heatid="6970" lane="7" />
                <RESULT eventid="1179" points="45" swimtime="00:02:26.37" resultid="4942" heatid="7002" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="4943" heatid="7030" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="1391" points="35" swimtime="00:06:24.35" resultid="4944" heatid="7092" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:49.45" />
                    <SPLIT distance="100" swimtime="00:03:29.81" />
                    <SPLIT distance="150" swimtime="00:05:04.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="4948" heatid="6999" lane="5" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4884" number="1" />
                    <RELAYPOSITION athleteid="4909" number="2" />
                    <RELAYPOSITION athleteid="4912" number="3" />
                    <RELAYPOSITION athleteid="4891" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kat. F /280 i starsi/" eventid="1149" points="10" swimtime="00:07:58.41" resultid="4945" heatid="6998" lane="8" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:51.19" />
                    <SPLIT distance="100" swimtime="00:05:05.66" />
                    <SPLIT distance="150" swimtime="00:06:46.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4900" number="1" />
                    <RELAYPOSITION athleteid="4904" number="2" />
                    <RELAYPOSITION athleteid="4940" number="3" />
                    <RELAYPOSITION athleteid="4930" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters w kat. F /280 i starsi/" eventid="1331" points="8" swimtime="00:07:55.38" resultid="4946" heatid="7073" lane="8" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:23.68" />
                    <SPLIT distance="100" swimtime="00:05:29.99" />
                    <SPLIT distance="150" swimtime="00:06:40.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4900" number="1" />
                    <RELAYPOSITION athleteid="4904" number="2" />
                    <RELAYPOSITION athleteid="4940" number="3" />
                    <RELAYPOSITION athleteid="4930" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1513" points="12" swimtime="00:06:47.52" resultid="4947" heatid="7147" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:06:09.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4900" number="1" />
                    <RELAYPOSITION athleteid="4904" number="2" />
                    <RELAYPOSITION athleteid="4884" number="3" />
                    <RELAYPOSITION athleteid="4907" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAGOR" name="Masters Gorzów" nation="POL" region="LBS">
          <CONTACT city="Kłodawa" name="Łopaciński" state="LUBUS" street="Dębowa" zip="66-415" />
          <ATHLETES>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="Wojciechowicz" nation="POL" athleteid="4960">
              <RESULTS>
                <RESULT eventid="1194" points="428" swimtime="00:01:02.24" resultid="4961" heatid="7018" lane="3" entrytime="00:01:03.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1376" points="347" swimtime="00:02:25.06" resultid="4962" heatid="7083" lane="4" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="316" swimtime="00:02:47.23" resultid="4963" heatid="7099" lane="5" entrytime="00:02:50.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="150" swimtime="00:02:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="395" swimtime="00:00:28.49" resultid="4964" heatid="7132" lane="9" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1573" points="330" swimtime="00:05:18.34" resultid="4965" heatid="7172" lane="2" entrytime="00:05:15.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                    <SPLIT distance="200" swimtime="00:02:33.67" />
                    <SPLIT distance="250" swimtime="00:03:15.67" />
                    <SPLIT distance="300" swimtime="00:03:58.41" />
                    <SPLIT distance="350" swimtime="00:04:40.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" athleteid="4966">
              <RESULTS>
                <RESULT eventid="1134" points="371" swimtime="00:00:33.44" resultid="4967" heatid="6995" lane="2" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1316" points="351" swimtime="00:01:13.59" resultid="4968" heatid="7071" lane="0" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="296" swimtime="00:02:50.97" resultid="4969" heatid="7101" lane="2" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:09.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="388" swimtime="00:00:28.65" resultid="4970" heatid="7131" lane="6" entrytime="00:00:28.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-22" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" athleteid="4971">
              <RESULTS>
                <RESULT eventid="1134" points="272" swimtime="00:00:37.10" resultid="4972" heatid="6993" lane="5" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1224" points="243" swimtime="00:02:58.58" resultid="4973" heatid="7028" lane="8" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="345" swimtime="00:00:31.97" resultid="4974" heatid="7042" lane="0" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1406" points="306" swimtime="00:02:49.14" resultid="4975" heatid="7099" lane="8" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:19.79" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="262" swimtime="00:01:17.81" resultid="4976" heatid="7110" lane="6" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1573" points="306" swimtime="00:05:26.43" resultid="4977" heatid="7172" lane="1" entrytime="00:05:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:55.55" />
                    <SPLIT distance="200" swimtime="00:02:38.09" />
                    <SPLIT distance="250" swimtime="00:03:21.17" />
                    <SPLIT distance="300" swimtime="00:04:04.11" />
                    <SPLIT distance="350" swimtime="00:04:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-11" firstname="Artur" gender="M" lastname="Łopacinski" nation="POL" athleteid="4978">
              <RESULTS>
                <RESULT eventid="1224" points="208" swimtime="00:03:07.99" resultid="4979" heatid="7027" lane="3" entrytime="00:03:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:13.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="336" swimtime="00:00:32.26" resultid="4980" heatid="7042" lane="9" entrytime="00:00:31.63" entrycourse="LCM" />
                <RESULT eventid="1406" points="276" swimtime="00:02:55.03" resultid="4981" heatid="7100" lane="6" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:21.19" />
                    <SPLIT distance="150" swimtime="00:02:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="347" swimtime="00:00:29.73" resultid="4982" heatid="7129" lane="2" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="1543" points="250" swimtime="00:01:32.97" resultid="4983" heatid="7157" lane="6" entrytime="00:01:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="359" swimtime="00:02:11.40" resultid="4984" heatid="7000" lane="6" entrytime="00:02:10.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:44.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4960" number="1" />
                    <RELAYPOSITION athleteid="4966" number="2" />
                    <RELAYPOSITION athleteid="4978" number="3" />
                    <RELAYPOSITION athleteid="4971" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="407" swimtime="00:01:54.49" resultid="4985" heatid="7075" lane="5" entrytime="00:01:54.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="100" swimtime="00:00:57.09" />
                    <SPLIT distance="150" swimtime="00:01:26.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4960" number="1" />
                    <RELAYPOSITION athleteid="4971" number="2" />
                    <RELAYPOSITION athleteid="4978" number="3" />
                    <RELAYPOSITION athleteid="4966" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LEWAR" name="SKT Legia Warszawa" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="sekcja@plywanielegia.pl" internet="www.plywanielegia.pl" name="Drzewiński Łukasz" phone="509268321" state="MAZ" street="ul. Myśliwiecka 4a" zip="00-459" />
          <ATHLETES>
            <ATHLETE birthdate="1984-04-09" firstname="Łukasz" gender="M" lastname="Drzewiński" nation="POL" license="066/14" athleteid="5029">
              <RESULTS>
                <RESULT eventid="1224" points="499" swimtime="00:02:20.54" resultid="5030" heatid="7029" lane="5" entrytime="00:02:18.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="582" swimtime="00:00:26.85" resultid="5031" heatid="7046" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1438" points="537" swimtime="00:01:01.27" resultid="5032" heatid="7112" lane="3" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" license="066/14" athleteid="5033">
              <RESULTS>
                <RESULT eventid="1194" points="512" swimtime="00:00:58.63" resultid="5034" heatid="7021" lane="9" entrytime="00:00:59.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="461" swimtime="00:00:27.06" resultid="5035" heatid="7135" lane="0" entrytime="00:00:26.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-17" firstname="Bartosz" gender="M" lastname="Korsak" nation="POL" license="066/14" athleteid="5036">
              <RESULTS>
                <RESULT eventid="1194" points="557" swimtime="00:00:56.99" resultid="5037" heatid="7022" lane="9" entrytime="00:00:57.50" />
                <RESULT eventid="1376" points="492" swimtime="00:02:09.16" resultid="5038" heatid="7090" lane="4" entrytime="00:02:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:05.58" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-16" firstname="Maciej" gender="M" lastname="Drzewiński" nation="POL" license="066/14" athleteid="5040">
              <RESULTS>
                <RESULT eventid="1468" points="434" swimtime="00:00:27.60" resultid="5041" heatid="7132" lane="7" entrytime="00:00:27.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-09" firstname="Tomasz" gender="M" lastname="Drzewiński" nation="POL" license="066/14" athleteid="5042">
              <RESULTS>
                <RESULT eventid="1468" points="265" swimtime="00:00:32.53" resultid="5043" heatid="7132" lane="2" entrytime="00:00:27.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-25" firstname="Andrzej" gender="M" lastname="Drzewiński" nation="POL" license="066/14" athleteid="5044">
              <RESULTS>
                <RESULT eventid="1286" points="106" swimtime="00:00:56.28" resultid="5045" heatid="7054" lane="7" entrytime="00:00:45.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-24" firstname="Maciej" gender="M" lastname="Grzelak" nation="POL" license="066/14" athleteid="5046">
              <RESULTS>
                <RESULT eventid="1194" points="250" swimtime="00:01:14.38" resultid="5047" heatid="7013" lane="1" entrytime="00:01:15.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="173" swimtime="00:03:19.74" resultid="5048" heatid="7026" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="150" swimtime="00:02:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="270" swimtime="00:00:34.69" resultid="5049" heatid="7039" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="5050" heatid="7097" lane="3" entrytime="00:03:15.00" />
                <RESULT eventid="1438" points="208" swimtime="00:01:24.02" resultid="5051" heatid="7108" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="257" swimtime="00:00:32.87" resultid="5052" heatid="7124" lane="5" entrytime="00:00:34.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" license="066/14" athleteid="5053">
              <RESULTS>
                <RESULT eventid="1468" points="450" swimtime="00:00:27.28" resultid="5054" heatid="7134" lane="3" entrytime="00:00:26.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-08-28" firstname="Krzesimir" gender="M" lastname="Sieczych" nation="POL" license="066/14" athleteid="5055">
              <RESULTS>
                <RESULT eventid="1194" points="393" swimtime="00:01:04.00" resultid="5056" heatid="7019" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="373" swimtime="00:00:31.14" resultid="5057" heatid="7043" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1468" points="404" swimtime="00:00:28.27" resultid="5058" heatid="7134" lane="8" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-11" firstname="Marta" gender="F" lastname="Sadomska" nation="POL" license="066/14" athleteid="5059">
              <RESULTS>
                <RESULT eventid="1453" points="467" swimtime="00:00:30.58" resultid="5060" heatid="7120" lane="6" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-22" firstname="Paweł" gender="M" lastname="Kozak" nation="POL" license="066/14" athleteid="5061">
              <RESULTS>
                <RESULT eventid="1194" status="DNS" swimtime="00:00:00.00" resultid="5062" heatid="7022" lane="7" entrytime="00:00:56.20" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="5063" heatid="7045" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1438" status="DNS" swimtime="00:00:00.00" resultid="5064" heatid="7112" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="5065" heatid="7135" lane="8" entrytime="00:00:26.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" license="066/14" athleteid="5066">
              <RESULTS>
                <RESULT eventid="1134" points="568" swimtime="00:00:29.02" resultid="5067" heatid="6997" lane="4" entrytime="00:00:27.49" />
                <RESULT eventid="1256" points="565" swimtime="00:00:27.13" resultid="5068" heatid="7046" lane="7" entrytime="00:00:26.30" />
                <RESULT eventid="1316" points="558" swimtime="00:01:03.06" resultid="5069" heatid="7072" lane="4" entrytime="00:00:59.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="550" swimtime="00:01:00.79" resultid="5071" heatid="7112" lane="6" entrytime="00:00:59.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="522" swimtime="00:02:18.93" resultid="5492" heatid="7146" lane="4" entrytime="00:02:14.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="6963" heatid="7103" lane="4" entrytime="00:02:14.81" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-21" firstname="Maciej" gender="M" lastname="Bień" nation="POL" license="066/14" athleteid="5072">
              <RESULTS>
                <RESULT eventid="1194" points="294" swimtime="00:01:10.51" resultid="5073" heatid="7015" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="346" swimtime="00:00:37.98" resultid="5074" heatid="7059" lane="9" entrytime="00:00:36.20" />
                <RESULT eventid="1468" points="297" swimtime="00:00:31.31" resultid="5075" heatid="7128" lane="5" entrytime="00:00:30.11" />
                <RESULT eventid="1543" points="291" swimtime="00:01:28.33" resultid="5076" heatid="7161" lane="7" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-20" firstname="Piotr" gender="M" lastname="Gęgotek" nation="POL" license="066/14" athleteid="5077">
              <RESULTS>
                <RESULT eventid="1468" points="498" swimtime="00:00:26.37" resultid="5078" heatid="7133" lane="5" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Piotr" gender="M" lastname="Krzakowski" nation="POL" athleteid="5500">
              <RESULTS>
                <RESULT eventid="1286" points="223" swimtime="00:00:43.92" resultid="5501" heatid="7058" lane="9" entrytime="00:00:37.20" />
                <RESULT eventid="1543" status="DNS" swimtime="00:00:00.00" resultid="5502" heatid="7159" lane="2" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" gender="M" lastname="Krzakowski" nation="POL" athleteid="6964" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1164" points="240" swimtime="00:02:30.25" resultid="6965" heatid="7001" lane="0" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:26.00" />
                    <SPLIT distance="150" swimtime="00:01:56.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5029" number="1" />
                    <RELAYPOSITION athleteid="5044" number="2" />
                    <RELAYPOSITION athleteid="5040" number="3" />
                    <RELAYPOSITION athleteid="5042" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1346" points="546" swimtime="00:01:43.80" resultid="6968" heatid="7076" lane="3" entrytime="00:01:46.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                    <SPLIT distance="100" swimtime="00:00:52.65" />
                    <SPLIT distance="150" swimtime="00:01:17.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5066" number="1" />
                    <RELAYPOSITION athleteid="5029" number="2" />
                    <RELAYPOSITION athleteid="5053" number="3" />
                    <RELAYPOSITION athleteid="5033" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1164" points="266" swimtime="00:02:25.11" resultid="6966" heatid="7001" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5055" number="1" />
                    <RELAYPOSITION athleteid="5072" number="2" />
                    <RELAYPOSITION athleteid="5046" number="3" />
                    <RELAYPOSITION athleteid="6964" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1346" points="458" swimtime="00:01:50.07" resultid="6969" heatid="7076" lane="7" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:00:57.16" />
                    <SPLIT distance="150" swimtime="00:01:24.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5072" number="1" />
                    <RELAYPOSITION athleteid="5040" number="2" />
                    <RELAYPOSITION athleteid="5055" number="3" />
                    <RELAYPOSITION athleteid="5077" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1164" points="491" swimtime="00:01:58.35" resultid="6967" heatid="7001" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:04.37" />
                    <SPLIT distance="150" swimtime="00:01:32.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5066" number="1" />
                    <RELAYPOSITION athleteid="5053" number="2" />
                    <RELAYPOSITION athleteid="5077" number="3" />
                    <RELAYPOSITION athleteid="5033" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAPAB" name="WOPR Masters Pabianice" nation="POL" region="LOD">
          <CONTACT city="Pabianice" email="jarowyrwa@onet.pl" name="Wyrwa Jarosław" phone="503574455" state="ŁÓDZK" street="St.Moniuszki 94 a m 6" zip="95-200" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-21" firstname="Jarosław" gender="M" lastname="Wyrwa" nation="POL" athleteid="5084">
              <RESULTS>
                <RESULT eventid="1286" points="312" swimtime="00:00:39.32" resultid="5085" heatid="7056" lane="5" entrytime="00:00:39.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIEDL" name="Siedlce" nation="POL">
          <CONTACT name="Jedrychowski" />
          <ATHLETES>
            <ATHLETE birthdate="1989-06-11" firstname="Adam" gender="M" lastname="Jędrychowski" nation="POL" athleteid="5087">
              <RESULTS>
                <RESULT eventid="1286" points="578" swimtime="00:00:32.01" resultid="5088" heatid="7061" lane="2" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1543" points="488" swimtime="00:01:14.39" resultid="5089" heatid="7163" lane="0" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASUW" name="Suwałki" nation="POL" region="PDL">
          <CONTACT name="Obukowicz" />
          <ATHLETES>
            <ATHLETE birthdate="1985-09-23" firstname="Marcin" gender="M" lastname="Obukowicz" nation="POL" athleteid="5091">
              <RESULTS>
                <RESULT eventid="1256" points="354" swimtime="00:00:31.69" resultid="5092" heatid="7035" lane="4" entrytime="00:00:58.00" entrycourse="LCM" />
                <RESULT eventid="1286" points="411" swimtime="00:00:35.85" resultid="5093" heatid="7060" lane="2" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="5094" heatid="7099" lane="4" entrytime="00:02:50.00" entrycourse="LCM" />
                <RESULT eventid="1573" points="199" swimtime="00:06:16.85" resultid="5095" heatid="7171" lane="6" entrytime="00:05:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:20.98" />
                    <SPLIT distance="150" swimtime="00:02:07.92" />
                    <SPLIT distance="200" swimtime="00:02:57.68" />
                    <SPLIT distance="250" swimtime="00:03:47.68" />
                    <SPLIT distance="300" swimtime="00:04:38.44" />
                    <SPLIT distance="350" swimtime="00:05:28.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-24" firstname="Michał" gender="M" lastname="Choiński" nation="POL" athleteid="5096">
              <RESULTS>
                <RESULT eventid="1256" points="563" swimtime="00:00:27.16" resultid="5097" heatid="7046" lane="1" entrytime="00:00:26.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UCWAR" name="UCSiR Warszawa" nation="POL" region="MAZ">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-03" firstname="ALICJA" gender="F" lastname="CICHA-MIKOŁAJCZYK" nation="POL" athleteid="5099">
              <RESULTS>
                <RESULT eventid="1119" points="64" swimtime="00:01:07.58" resultid="5100" heatid="6982" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1179" points="85" swimtime="00:01:58.29" resultid="5101" heatid="7003" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="55" swimtime="00:02:32.05" resultid="5102" heatid="7063" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="77" swimtime="00:04:24.77" resultid="5103" heatid="7077" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.42" />
                    <SPLIT distance="100" swimtime="00:02:07.03" />
                    <SPLIT distance="150" swimtime="00:03:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="115" swimtime="00:00:48.66" resultid="5104" heatid="7115" lane="7" entrytime="00:00:49.00" />
                <RESULT eventid="1483" points="57" swimtime="00:05:23.11" resultid="5105" heatid="7137" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.91" />
                    <SPLIT distance="100" swimtime="00:02:41.61" />
                    <SPLIT distance="150" swimtime="00:04:02.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-26" firstname="MAŁGORZATA" gender="F" lastname="KOTAŃSKA" nation="POL" athleteid="5106">
              <RESULTS>
                <RESULT eventid="1058" points="237" swimtime="00:03:46.14" resultid="5107" heatid="6972" lane="7" entrytime="00:03:31.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                    <SPLIT distance="100" swimtime="00:01:46.10" />
                    <SPLIT distance="150" swimtime="00:02:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="165" swimtime="00:01:34.85" resultid="5108" heatid="7004" lane="5" entrytime="00:01:25.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="261" swimtime="00:00:46.63" resultid="5109" heatid="7050" lane="0" entrytime="00:00:44.06" />
                <RESULT eventid="1361" status="DNS" swimtime="00:00:00.00" resultid="5110" heatid="7078" lane="4" entrytime="00:03:16.00" />
                <RESULT eventid="1453" points="209" swimtime="00:00:39.93" resultid="5111" heatid="7116" lane="3" entrytime="00:00:38.39" />
                <RESULT eventid="1528" points="241" swimtime="00:01:43.46" resultid="5112" heatid="7153" lane="9" entrytime="00:01:37.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-16" firstname="MONIKA" gender="F" lastname="KURYŁOWICZ" nation="POL" athleteid="5113">
              <RESULTS>
                <RESULT eventid="1179" points="208" swimtime="00:01:27.78" resultid="5114" heatid="7005" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="193" swimtime="00:03:15.50" resultid="5115" heatid="7079" lane="8" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:35.91" />
                    <SPLIT distance="150" swimtime="00:02:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="231" swimtime="00:00:38.63" resultid="5116" heatid="7116" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1558" points="194" swimtime="00:06:53.00" resultid="5117" heatid="7165" lane="7" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                    <SPLIT distance="100" swimtime="00:01:37.47" />
                    <SPLIT distance="150" swimtime="00:02:30.84" />
                    <SPLIT distance="200" swimtime="00:03:24.76" />
                    <SPLIT distance="250" swimtime="00:04:18.26" />
                    <SPLIT distance="300" swimtime="00:05:11.90" />
                    <SPLIT distance="350" swimtime="00:06:05.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="MICHAŁ" gender="M" lastname="NOWAK" nation="POL" athleteid="5118">
              <RESULTS>
                <RESULT eventid="1104" points="272" swimtime="00:03:16.44" resultid="5119" heatid="6978" lane="0" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:30.71" />
                    <SPLIT distance="150" swimtime="00:02:22.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="369" swimtime="00:00:37.17" resultid="5120" heatid="7058" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1406" points="212" swimtime="00:03:10.90" resultid="5121" heatid="7098" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:35.82" />
                    <SPLIT distance="150" swimtime="00:02:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1438" points="142" swimtime="00:01:35.43" resultid="5122" heatid="7108" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1543" points="331" swimtime="00:01:24.64" resultid="5123" heatid="7159" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="MICHAŁ" gender="M" lastname="RYBARCZYK" nation="POL" athleteid="5124">
              <RESULTS>
                <RESULT eventid="1134" points="168" swimtime="00:00:43.54" resultid="5125" heatid="6991" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1194" points="368" swimtime="00:01:05.43" resultid="5126" heatid="7018" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="287" swimtime="00:00:33.99" resultid="5127" heatid="7041" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1376" points="286" swimtime="00:02:34.76" resultid="5128" heatid="7087" lane="8" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:54.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="376" swimtime="00:00:28.95" resultid="5129" heatid="7130" lane="5" entrytime="00:00:28.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="RYSZARD" gender="M" lastname="RYBARCZYK" nation="POL" athleteid="5130">
              <RESULTS>
                <RESULT eventid="1286" points="199" swimtime="00:00:45.65" resultid="5131" heatid="7055" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1468" points="154" swimtime="00:00:38.99" resultid="5132" heatid="7122" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="MACIEJ" gender="M" lastname="RYBICKI" nation="POL" athleteid="5133">
              <RESULTS>
                <RESULT eventid="1468" status="DNS" swimtime="00:00:00.00" resultid="5134" heatid="7127" lane="8" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-16" firstname="OLGA" gender="F" lastname="SCHAAF" nation="POL" athleteid="5135">
              <RESULTS>
                <RESULT eventid="1179" points="355" swimtime="00:01:13.52" resultid="5136" heatid="7007" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="357" swimtime="00:00:33.45" resultid="5137" heatid="7118" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1558" points="270" swimtime="00:06:09.84" resultid="5138" heatid="7166" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                    <SPLIT distance="200" swimtime="00:02:55.42" />
                    <SPLIT distance="250" swimtime="00:03:44.17" />
                    <SPLIT distance="300" swimtime="00:04:33.41" />
                    <SPLIT distance="350" swimtime="00:05:23.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-26" firstname="URSZULA" gender="F" lastname="BIELAWSKA" nation="POL" athleteid="5139">
              <RESULTS>
                <RESULT eventid="1058" points="280" swimtime="00:03:34.18" resultid="5140" heatid="6972" lane="1" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="100" swimtime="00:01:41.93" />
                    <SPLIT distance="150" swimtime="00:02:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="379" swimtime="00:01:11.91" resultid="5141" heatid="7007" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="304" swimtime="00:00:44.29" resultid="5142" heatid="7050" lane="9" entrytime="00:00:44.50" />
                <RESULT eventid="1361" points="332" swimtime="00:02:43.00" resultid="5143" heatid="7080" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="373" swimtime="00:00:32.95" resultid="5144" heatid="7118" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1558" points="313" swimtime="00:05:52.01" resultid="5145" heatid="7166" lane="4" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:05.92" />
                    <SPLIT distance="200" swimtime="00:02:51.12" />
                    <SPLIT distance="250" swimtime="00:03:37.17" />
                    <SPLIT distance="300" swimtime="00:04:23.55" />
                    <SPLIT distance="350" swimtime="00:05:09.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STSWI" name="Stowarzyszenie Pływackie &quot;Swimmers&quot;" nation="POL" region="14">
          <ATHLETES>
            <ATHLETE birthdate="1976-01-01" firstname="Remigiusz" gender="M" lastname="Gołebiowski " nation="POL" athleteid="5488">
              <RESULTS>
                <RESULT eventid="1256" points="402" swimtime="00:00:30.38" resultid="5490" heatid="7045" lane="9" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWWAR" name="AZS SWPS Warszawa" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" name="Mroczek" phone="500 231 093" street="Malwowa" />
          <ATHLETES>
            <ATHLETE birthdate="1991-12-15" firstname="Antoni" gender="M" lastname="Kląskała-Mroczek" nation="POL" athleteid="5684">
              <RESULTS>
                <RESULT eventid="1134" points="439" swimtime="00:00:31.62" resultid="5685" heatid="6997" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1316" points="375" swimtime="00:01:11.97" resultid="5686" heatid="7072" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="325" swimtime="00:02:42.76" resultid="5687" heatid="7146" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="150" swimtime="00:02:02.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

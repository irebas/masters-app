<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SMS SwimArt Myślenice" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Łódź" name="Zimowe Mistrzostwa Polskiw Pływaniu Masters" course="SCM" deadline="2019-10-30" hostclub="UTW Masters Zgierz" hostclub.url="https://www.swimart.pl" organizer="Masters Łódź" reservecount="2" result.url="https://www.megatiming.pl" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2019-11-17" type="YEAR" />
      <POOL name="Zatoka Sportu Politechniki Łódzkiej" lanemax="9" />
      <FACILITY city="Łódź" name="Zatoka Sportu Politechniki Łódzkiej" nation="POL" street="Aleja Politechniki 10" zip="93-590" />
      <POINTTABLE pointtableid="3012" name="FINA Point Scoring" version="2019" />
      <CONTACT email="zawody@swimart.pl" name="Artur Żak" phone="501 689 458" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="15500" />
      </FEES>
      <SESSIONS>
        <SESSION date="2019-11-15" daytime="14:00" endtime="19:55" name="Zimowe Mistrzostwa Polskiw Pływaniu Masters BLOK I" number="1" warmupfrom="13:00" warmupuntil="13:45">
          <EVENTS>
            <EVENT eventid="1059" daytime="14:00" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="1062" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="1064" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3777" />
                    <RANKING order="2" place="2" resultid="4096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4121" />
                    <RANKING order="2" place="2" resultid="4235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3787" />
                    <RANKING order="2" place="2" resultid="5662" />
                    <RANKING order="3" place="3" resultid="5960" />
                    <RANKING order="4" place="4" resultid="4130" />
                    <RANKING order="5" place="5" resultid="4164" />
                    <RANKING order="6" place="6" resultid="3771" />
                    <RANKING order="7" place="-1" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4821" />
                    <RANKING order="2" place="2" resultid="2470" />
                    <RANKING order="3" place="3" resultid="4114" />
                    <RANKING order="4" place="4" resultid="3807" />
                    <RANKING order="5" place="5" resultid="4146" />
                    <RANKING order="6" place="6" resultid="2307" />
                    <RANKING order="7" place="7" resultid="3907" />
                    <RANKING order="8" place="8" resultid="2589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3103" />
                    <RANKING order="2" place="2" resultid="4770" />
                    <RANKING order="3" place="3" resultid="5797" />
                    <RANKING order="4" place="4" resultid="4057" />
                    <RANKING order="5" place="5" resultid="4073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3987" />
                    <RANKING order="2" place="2" resultid="4268" />
                    <RANKING order="3" place="3" resultid="2368" />
                    <RANKING order="4" place="4" resultid="6201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3154" />
                    <RANKING order="2" place="2" resultid="5803" />
                    <RANKING order="3" place="3" resultid="4701" />
                    <RANKING order="4" place="4" resultid="2079" />
                    <RANKING order="5" place="5" resultid="5088" />
                    <RANKING order="6" place="6" resultid="3916" />
                    <RANKING order="7" place="7" resultid="4372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3173" />
                    <RANKING order="2" place="2" resultid="4987" />
                    <RANKING order="3" place="3" resultid="3691" />
                    <RANKING order="4" place="4" resultid="2932" />
                    <RANKING order="5" place="5" resultid="6163" />
                    <RANKING order="6" place="6" resultid="5108" />
                    <RANKING order="7" place="7" resultid="5508" />
                    <RANKING order="8" place="8" resultid="5261" />
                    <RANKING order="9" place="9" resultid="3525" />
                    <RANKING order="10" place="10" resultid="5735" />
                    <RANKING order="11" place="11" resultid="3275" />
                    <RANKING order="12" place="12" resultid="5641" />
                    <RANKING order="13" place="13" resultid="3301" />
                    <RANKING order="14" place="14" resultid="5947" />
                    <RANKING order="15" place="-1" resultid="3956" />
                    <RANKING order="16" place="-1" resultid="6410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3379" />
                    <RANKING order="2" place="2" resultid="2439" />
                    <RANKING order="3" place="3" resultid="2815" />
                    <RANKING order="4" place="4" resultid="4946" />
                    <RANKING order="5" place="5" resultid="4416" />
                    <RANKING order="6" place="6" resultid="6224" />
                    <RANKING order="7" place="7" resultid="5600" />
                    <RANKING order="8" place="8" resultid="4012" />
                    <RANKING order="9" place="9" resultid="5609" />
                    <RANKING order="10" place="10" resultid="3386" />
                    <RANKING order="11" place="11" resultid="2652" />
                    <RANKING order="12" place="-1" resultid="4023" />
                    <RANKING order="13" place="-1" resultid="5646" />
                    <RANKING order="14" place="-1" resultid="6390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1060" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5808" />
                    <RANKING order="2" place="2" resultid="5242" />
                    <RANKING order="3" place="3" resultid="4037" />
                    <RANKING order="4" place="4" resultid="3701" />
                    <RANKING order="5" place="5" resultid="2827" />
                    <RANKING order="6" place="6" resultid="2645" />
                    <RANKING order="7" place="7" resultid="3877" />
                    <RANKING order="8" place="8" resultid="3469" />
                    <RANKING order="9" place="9" resultid="5575" />
                    <RANKING order="10" place="10" resultid="5019" />
                    <RANKING order="11" place="11" resultid="3391" />
                    <RANKING order="12" place="12" resultid="6459" />
                    <RANKING order="13" place="13" resultid="4338" />
                    <RANKING order="14" place="14" resultid="4473" />
                    <RANKING order="15" place="15" resultid="3592" />
                    <RANKING order="16" place="-1" resultid="2990" />
                    <RANKING order="17" place="-1" resultid="3111" />
                    <RANKING order="18" place="-1" resultid="3515" />
                    <RANKING order="19" place="-1" resultid="4538" />
                    <RANKING order="20" place="-1" resultid="4660" />
                    <RANKING order="21" place="-1" resultid="5209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6335" />
                    <RANKING order="2" place="2" resultid="2980" />
                    <RANKING order="3" place="3" resultid="2034" />
                    <RANKING order="4" place="4" resultid="2777" />
                    <RANKING order="5" place="5" resultid="4523" />
                    <RANKING order="6" place="6" resultid="5836" />
                    <RANKING order="7" place="7" resultid="3868" />
                    <RANKING order="8" place="8" resultid="4685" />
                    <RANKING order="9" place="9" resultid="3328" />
                    <RANKING order="10" place="10" resultid="3464" />
                    <RANKING order="11" place="11" resultid="5842" />
                    <RANKING order="12" place="12" resultid="3483" />
                    <RANKING order="13" place="13" resultid="3293" />
                    <RANKING order="14" place="14" resultid="2744" />
                    <RANKING order="15" place="15" resultid="5119" />
                    <RANKING order="16" place="16" resultid="2228" />
                    <RANKING order="17" place="17" resultid="4383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2618" />
                    <RANKING order="2" place="2" resultid="3735" />
                    <RANKING order="3" place="3" resultid="4015" />
                    <RANKING order="4" place="4" resultid="2770" />
                    <RANKING order="5" place="5" resultid="3537" />
                    <RANKING order="6" place="6" resultid="2674" />
                    <RANKING order="7" place="-1" resultid="3833" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7234" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7235" daytime="14:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7236" daytime="14:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7237" daytime="14:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7238" daytime="14:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7239" daytime="14:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7240" daytime="14:09" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7241" daytime="14:11" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7242" daytime="14:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7243" daytime="14:13" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7244" daytime="14:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7245" daytime="14:16" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="17:15" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7647" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7648" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7649" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7650" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7651" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3096" />
                    <RANKING order="2" place="2" resultid="5165" />
                    <RANKING order="3" place="3" resultid="4780" />
                    <RANKING order="4" place="4" resultid="2420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7652" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3925" />
                    <RANKING order="2" place="2" resultid="2089" />
                    <RANKING order="3" place="3" resultid="2103" />
                    <RANKING order="4" place="4" resultid="2763" />
                    <RANKING order="5" place="-1" resultid="3649" />
                    <RANKING order="6" place="-1" resultid="5677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7653" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5694" />
                    <RANKING order="2" place="2" resultid="2837" />
                    <RANKING order="3" place="3" resultid="4653" />
                    <RANKING order="4" place="4" resultid="2604" />
                    <RANKING order="5" place="-1" resultid="3212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7654" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4393" />
                    <RANKING order="2" place="2" resultid="6098" />
                    <RANKING order="3" place="3" resultid="6035" />
                    <RANKING order="4" place="4" resultid="2567" />
                    <RANKING order="5" place="-1" resultid="2218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7655" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2290" />
                    <RANKING order="2" place="2" resultid="5991" />
                    <RANKING order="3" place="3" resultid="2806" />
                    <RANKING order="4" place="4" resultid="5521" />
                    <RANKING order="5" place="5" resultid="6248" />
                    <RANKING order="6" place="6" resultid="4806" />
                    <RANKING order="7" place="-1" resultid="2002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7656" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4254" />
                    <RANKING order="2" place="2" resultid="3324" />
                    <RANKING order="3" place="3" resultid="6107" />
                    <RANKING order="4" place="4" resultid="6193" />
                    <RANKING order="5" place="5" resultid="5703" />
                    <RANKING order="6" place="6" resultid="5722" />
                    <RANKING order="7" place="7" resultid="2809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7657" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2044" />
                    <RANKING order="2" place="2" resultid="4624" />
                    <RANKING order="3" place="3" resultid="6006" />
                    <RANKING order="4" place="4" resultid="2878" />
                    <RANKING order="5" place="5" resultid="4693" />
                    <RANKING order="6" place="6" resultid="2110" />
                    <RANKING order="7" place="7" resultid="3042" />
                    <RANKING order="8" place="8" resultid="5920" />
                    <RANKING order="9" place="9" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7658" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6024" />
                    <RANKING order="2" place="2" resultid="6181" />
                    <RANKING order="3" place="3" resultid="2541" />
                    <RANKING order="4" place="4" resultid="5787" />
                    <RANKING order="5" place="5" resultid="4503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7659" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5855" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="2584" />
                    <RANKING order="4" place="4" resultid="5913" />
                    <RANKING order="5" place="5" resultid="3265" />
                    <RANKING order="6" place="-1" resultid="6366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7660" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2518" />
                    <RANKING order="2" place="2" resultid="6255" />
                    <RANKING order="3" place="3" resultid="3508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7661" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3822" />
                    <RANKING order="2" place="2" resultid="4512" />
                    <RANKING order="3" place="3" resultid="2317" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7294" daytime="17:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7295" daytime="17:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7296" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7297" daytime="17:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7298" daytime="18:03" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7299" daytime="18:18" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1761" />
                <TIMESTANDARDREF timestandardlistid="1773" />
                <TIMESTANDARDREF timestandardlistid="1779" />
                <TIMESTANDARDREF timestandardlistid="1785" />
                <TIMESTANDARDREF timestandardlistid="1791" />
                <TIMESTANDARDREF timestandardlistid="1797" />
                <TIMESTANDARDREF timestandardlistid="1803" />
                <TIMESTANDARDREF timestandardlistid="1809" />
                <TIMESTANDARDREF timestandardlistid="1815" />
                <TIMESTANDARDREF timestandardlistid="1821" />
                <TIMESTANDARDREF timestandardlistid="1827" />
                <TIMESTANDARDREF timestandardlistid="1833" />
                <TIMESTANDARDREF timestandardlistid="1839" />
                <TIMESTANDARDREF timestandardlistid="1845" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1076" daytime="14:18" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7587" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7588" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2242" />
                    <RANKING order="2" place="-1" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7589" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4099" />
                    <RANKING order="2" place="2" resultid="4563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7590" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5684" />
                    <RANKING order="2" place="2" resultid="4648" />
                    <RANKING order="3" place="3" resultid="4170" />
                    <RANKING order="4" place="4" resultid="3940" />
                    <RANKING order="5" place="5" resultid="4814" />
                    <RANKING order="6" place="6" resultid="2692" />
                    <RANKING order="7" place="7" resultid="2505" />
                    <RANKING order="8" place="8" resultid="2701" />
                    <RANKING order="9" place="-1" resultid="5173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7591" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3794" />
                    <RANKING order="2" place="2" resultid="2199" />
                    <RANKING order="3" place="3" resultid="3125" />
                    <RANKING order="4" place="4" resultid="4779" />
                    <RANKING order="5" place="5" resultid="2096" />
                    <RANKING order="6" place="6" resultid="4065" />
                    <RANKING order="7" place="7" resultid="3814" />
                    <RANKING order="8" place="8" resultid="2683" />
                    <RANKING order="9" place="-1" resultid="3946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7592" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4597" />
                    <RANKING order="2" place="2" resultid="2125" />
                    <RANKING order="3" place="3" resultid="2088" />
                    <RANKING order="4" place="4" resultid="3924" />
                    <RANKING order="5" place="5" resultid="5776" />
                    <RANKING order="6" place="6" resultid="3136" />
                    <RANKING order="7" place="7" resultid="5933" />
                    <RANKING order="8" place="8" resultid="2102" />
                    <RANKING order="9" place="9" resultid="2298" />
                    <RANKING order="10" place="-1" resultid="3648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7593" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5552" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="3184" />
                    <RANKING order="4" place="4" resultid="3764" />
                    <RANKING order="5" place="5" resultid="6499" />
                    <RANKING order="6" place="6" resultid="5812" />
                    <RANKING order="7" place="7" resultid="4155" />
                    <RANKING order="8" place="8" resultid="4652" />
                    <RANKING order="9" place="9" resultid="3239" />
                    <RANKING order="10" place="10" resultid="2756" />
                    <RANKING order="11" place="11" resultid="4843" />
                    <RANKING order="12" place="-1" resultid="2474" />
                    <RANKING order="13" place="-1" resultid="5529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7594" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2411" />
                    <RANKING order="2" place="2" resultid="3852" />
                    <RANKING order="3" place="3" resultid="4615" />
                    <RANKING order="4" place="4" resultid="2429" />
                    <RANKING order="5" place="5" resultid="5181" />
                    <RANKING order="6" place="6" resultid="3411" />
                    <RANKING order="7" place="7" resultid="5727" />
                    <RANKING order="8" place="8" resultid="4797" />
                    <RANKING order="9" place="9" resultid="2972" />
                    <RANKING order="10" place="10" resultid="6115" />
                    <RANKING order="11" place="11" resultid="3289" />
                    <RANKING order="12" place="12" resultid="3118" />
                    <RANKING order="13" place="13" resultid="6482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7595" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6304" />
                    <RANKING order="2" place="2" resultid="5617" />
                    <RANKING order="3" place="3" resultid="5635" />
                    <RANKING order="4" place="4" resultid="5753" />
                    <RANKING order="5" place="5" resultid="2289" />
                    <RANKING order="6" place="6" resultid="3010" />
                    <RANKING order="7" place="7" resultid="5990" />
                    <RANKING order="8" place="8" resultid="4578" />
                    <RANKING order="9" place="9" resultid="5520" />
                    <RANKING order="10" place="10" resultid="2718" />
                    <RANKING order="11" place="11" resultid="3220" />
                    <RANKING order="12" place="12" resultid="3180" />
                    <RANKING order="13" place="13" resultid="4805" />
                    <RANKING order="14" place="14" resultid="4518" />
                    <RANKING order="15" place="15" resultid="2462" />
                    <RANKING order="16" place="16" resultid="2524" />
                    <RANKING order="17" place="17" resultid="3626" />
                    <RANKING order="18" place="18" resultid="5139" />
                    <RANKING order="19" place="19" resultid="4289" />
                    <RANKING order="20" place="20" resultid="2230" />
                    <RANKING order="21" place="21" resultid="4296" />
                    <RANKING order="22" place="22" resultid="3963" />
                    <RANKING order="23" place="23" resultid="5082" />
                    <RANKING order="24" place="-1" resultid="2001" />
                    <RANKING order="25" place="-1" resultid="6468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7596" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6145" />
                    <RANKING order="2" place="2" resultid="4558" />
                    <RANKING order="3" place="3" resultid="4253" />
                    <RANKING order="4" place="4" resultid="2359" />
                    <RANKING order="5" place="5" resultid="4247" />
                    <RANKING order="6" place="6" resultid="3682" />
                    <RANKING order="7" place="7" resultid="3740" />
                    <RANKING order="8" place="8" resultid="2666" />
                    <RANKING order="9" place="9" resultid="6344" />
                    <RANKING order="10" place="10" resultid="4385" />
                    <RANKING order="11" place="11" resultid="3633" />
                    <RANKING order="12" place="12" resultid="3396" />
                    <RANKING order="13" place="13" resultid="3323" />
                    <RANKING order="14" place="14" resultid="3754" />
                    <RANKING order="15" place="15" resultid="5702" />
                    <RANKING order="16" place="16" resultid="4527" />
                    <RANKING order="17" place="17" resultid="3673" />
                    <RANKING order="18" place="18" resultid="6192" />
                    <RANKING order="19" place="19" resultid="5927" />
                    <RANKING order="20" place="20" resultid="3614" />
                    <RANKING order="21" place="21" resultid="3131" />
                    <RANKING order="22" place="22" resultid="5200" />
                    <RANKING order="23" place="23" resultid="5721" />
                    <RANKING order="24" place="24" resultid="6106" />
                    <RANKING order="25" place="25" resultid="3058" />
                    <RANKING order="26" place="26" resultid="3993" />
                    <RANKING order="27" place="27" resultid="5826" />
                    <RANKING order="28" place="-1" resultid="4425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7597" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2993" />
                    <RANKING order="2" place="2" resultid="4928" />
                    <RANKING order="3" place="3" resultid="6371" />
                    <RANKING order="4" place="4" resultid="3199" />
                    <RANKING order="5" place="5" resultid="6042" />
                    <RANKING order="6" place="6" resultid="6380" />
                    <RANKING order="7" place="7" resultid="3019" />
                    <RANKING order="8" place="8" resultid="6005" />
                    <RANKING order="9" place="9" resultid="6341" />
                    <RANKING order="10" place="10" resultid="4692" />
                    <RANKING order="11" place="11" resultid="6136" />
                    <RANKING order="12" place="12" resultid="6377" />
                    <RANKING order="13" place="13" resultid="4959" />
                    <RANKING order="14" place="14" resultid="5713" />
                    <RANKING order="15" place="15" resultid="6186" />
                    <RANKING order="16" place="16" resultid="4314" />
                    <RANKING order="17" place="17" resultid="5013" />
                    <RANKING order="18" place="18" resultid="5095" />
                    <RANKING order="19" place="19" resultid="2053" />
                    <RANKING order="20" place="20" resultid="5626" />
                    <RANKING order="21" place="21" resultid="5038" />
                    <RANKING order="22" place="22" resultid="4881" />
                    <RANKING order="23" place="23" resultid="3253" />
                    <RANKING order="24" place="24" resultid="2490" />
                    <RANKING order="25" place="25" resultid="4908" />
                    <RANKING order="26" place="26" resultid="2985" />
                    <RANKING order="27" place="27" resultid="2066" />
                    <RANKING order="28" place="28" resultid="4830" />
                    <RANKING order="29" place="29" resultid="3141" />
                    <RANKING order="30" place="30" resultid="5254" />
                    <RANKING order="31" place="31" resultid="2737" />
                    <RANKING order="32" place="-1" resultid="2029" />
                    <RANKING order="33" place="-1" resultid="2899" />
                    <RANKING order="34" place="-1" resultid="4706" />
                    <RANKING order="35" place="-1" resultid="4984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7598" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4731" />
                    <RANKING order="2" place="2" resultid="3717" />
                    <RANKING order="3" place="3" resultid="6014" />
                    <RANKING order="4" place="4" resultid="5044" />
                    <RANKING order="5" place="5" resultid="3589" />
                    <RANKING order="6" place="6" resultid="2964" />
                    <RANKING order="7" place="7" resultid="4421" />
                    <RANKING order="8" place="8" resultid="6090" />
                    <RANKING order="9" place="9" resultid="2378" />
                    <RANKING order="10" place="10" resultid="4990" />
                    <RANKING order="11" place="11" resultid="5204" />
                    <RANKING order="12" place="12" resultid="4345" />
                    <RANKING order="13" place="13" resultid="5219" />
                    <RANKING order="14" place="14" resultid="5214" />
                    <RANKING order="15" place="15" resultid="5584" />
                    <RANKING order="16" place="16" resultid="6023" />
                    <RANKING order="17" place="17" resultid="4965" />
                    <RANKING order="18" place="18" resultid="5786" />
                    <RANKING order="19" place="19" resultid="3429" />
                    <RANKING order="20" place="20" resultid="4886" />
                    <RANKING order="21" place="21" resultid="2540" />
                    <RANKING order="22" place="22" resultid="2239" />
                    <RANKING order="23" place="23" resultid="5051" />
                    <RANKING order="24" place="24" resultid="4999" />
                    <RANKING order="25" place="25" resultid="2445" />
                    <RANKING order="26" place="26" resultid="6863" />
                    <RANKING order="27" place="27" resultid="4460" />
                    <RANKING order="28" place="28" resultid="2459" />
                    <RANKING order="29" place="-1" resultid="2024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7599" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4283" />
                    <RANKING order="2" place="2" resultid="2956" />
                    <RANKING order="3" place="3" resultid="2853" />
                    <RANKING order="4" place="4" resultid="4395" />
                    <RANKING order="5" place="5" resultid="3487" />
                    <RANKING order="6" place="6" resultid="2951" />
                    <RANKING order="7" place="7" resultid="2974" />
                    <RANKING order="8" place="8" resultid="3860" />
                    <RANKING order="9" place="9" resultid="2212" />
                    <RANKING order="10" place="10" resultid="4241" />
                    <RANKING order="11" place="11" resultid="5248" />
                    <RANKING order="12" place="12" resultid="6233" />
                    <RANKING order="13" place="13" resultid="4994" />
                    <RANKING order="14" place="14" resultid="2150" />
                    <RANKING order="15" place="15" resultid="4310" />
                    <RANKING order="16" place="16" resultid="3264" />
                    <RANKING order="17" place="17" resultid="2845" />
                    <RANKING order="18" place="-1" resultid="2987" />
                    <RANKING order="19" place="-1" resultid="3434" />
                    <RANKING order="20" place="-1" resultid="3542" />
                    <RANKING order="21" place="-1" resultid="3546" />
                    <RANKING order="22" place="-1" resultid="4469" />
                    <RANKING order="23" place="-1" resultid="4674" />
                    <RANKING order="24" place="-1" resultid="6365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7600" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2146" />
                    <RANKING order="2" place="2" resultid="3727" />
                    <RANKING order="3" place="3" resultid="4630" />
                    <RANKING order="4" place="4" resultid="5145" />
                    <RANKING order="5" place="5" resultid="2579" />
                    <RANKING order="6" place="6" resultid="5230" />
                    <RANKING order="7" place="7" resultid="2402" />
                    <RANKING order="8" place="8" resultid="3507" />
                    <RANKING order="9" place="9" resultid="6051" />
                    <RANKING order="10" place="10" resultid="6350" />
                    <RANKING order="11" place="11" resultid="2907" />
                    <RANKING order="12" place="12" resultid="3015" />
                    <RANKING order="13" place="13" resultid="2175" />
                    <RANKING order="14" place="14" resultid="5225" />
                    <RANKING order="15" place="15" resultid="6439" />
                    <RANKING order="16" place="16" resultid="3581" />
                    <RANKING order="17" place="17" resultid="3473" />
                    <RANKING order="18" place="18" resultid="2513" />
                    <RANKING order="19" place="19" resultid="3578" />
                    <RANKING order="20" place="20" resultid="3574" />
                    <RANKING order="21" place="21" resultid="2405" />
                    <RANKING order="22" place="22" resultid="2208" />
                    <RANKING order="23" place="23" resultid="3535" />
                    <RANKING order="24" place="24" resultid="3576" />
                    <RANKING order="25" place="25" resultid="3533" />
                    <RANKING order="26" place="26" resultid="3531" />
                    <RANKING order="27" place="-1" resultid="2183" />
                    <RANKING order="28" place="-1" resultid="2188" />
                    <RANKING order="29" place="-1" resultid="2335" />
                    <RANKING order="30" place="-1" resultid="2959" />
                    <RANKING order="31" place="-1" resultid="3452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7601" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4200" />
                    <RANKING order="2" place="2" resultid="6360" />
                    <RANKING order="3" place="3" resultid="2609" />
                    <RANKING order="4" place="4" resultid="3821" />
                    <RANKING order="5" place="5" resultid="2316" />
                    <RANKING order="6" place="6" resultid="3477" />
                    <RANKING order="7" place="7" resultid="4511" />
                    <RANKING order="8" place="8" resultid="3893" />
                    <RANKING order="9" place="9" resultid="2659" />
                    <RANKING order="10" place="10" resultid="3585" />
                    <RANKING order="11" place="11" resultid="3975" />
                    <RANKING order="12" place="12" resultid="2154" />
                    <RANKING order="13" place="-1" resultid="2627" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7246" daytime="14:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7247" daytime="14:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7248" daytime="14:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7249" daytime="14:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7250" daytime="14:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7251" daytime="14:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7252" daytime="14:27" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7253" daytime="14:29" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7254" daytime="14:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7255" daytime="14:31" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7256" daytime="14:32" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7257" daytime="14:34" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7258" daytime="14:35" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7259" daytime="14:36" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7260" daytime="14:38" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7261" daytime="14:39" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7262" daytime="14:40" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7263" daytime="14:41" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7264" daytime="14:42" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="7265" daytime="14:44" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="7266" daytime="14:45" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="7267" daytime="14:46" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="7268" daytime="14:47" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="7269" daytime="14:48" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="7270" daytime="14:50" number="25" order="25" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="19:42" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7677" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7678" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7679" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7680" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2636" />
                    <RANKING order="2" place="2" resultid="4815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7681" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7682" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="2" resultid="5777" />
                    <RANKING order="3" place="3" resultid="4108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7683" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5282" />
                    <RANKING order="2" place="2" resultid="3259" />
                    <RANKING order="3" place="3" resultid="6500" />
                    <RANKING order="4" place="4" resultid="5862" />
                    <RANKING order="5" place="-1" resultid="6494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7684" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5182" />
                    <RANKING order="2" place="2" resultid="6116" />
                    <RANKING order="3" place="3" resultid="2885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7685" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5818" />
                    <RANKING order="2" place="2" resultid="2386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7686" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6146" />
                    <RANKING order="2" place="2" resultid="3397" />
                    <RANKING order="3" place="3" resultid="3755" />
                    <RANKING order="4" place="4" resultid="3674" />
                    <RANKING order="5" place="5" resultid="5075" />
                    <RANKING order="6" place="6" resultid="4001" />
                    <RANKING order="7" place="-1" resultid="2529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7687" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6137" />
                    <RANKING order="2" place="2" resultid="3233" />
                    <RANKING order="3" place="3" resultid="5714" />
                    <RANKING order="4" place="4" resultid="5006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7688" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6416" />
                    <RANKING order="2" place="-1" resultid="4329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7689" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2975" />
                    <RANKING order="2" place="-1" resultid="6432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7690" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7691" agemax="24" agemin="20" name="0" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7302" daytime="19:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7303" daytime="20:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7304" daytime="20:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7305" daytime="20:59" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1884" />
                <TIMESTANDARDREF timestandardlistid="1890" />
                <TIMESTANDARDREF timestandardlistid="1896" />
                <TIMESTANDARDREF timestandardlistid="1902" />
                <TIMESTANDARDREF timestandardlistid="1908" />
                <TIMESTANDARDREF timestandardlistid="1914" />
                <TIMESTANDARDREF timestandardlistid="1920" />
                <TIMESTANDARDREF timestandardlistid="1926" />
                <TIMESTANDARDREF timestandardlistid="1932" />
                <TIMESTANDARDREF timestandardlistid="1938" />
                <TIMESTANDARDREF timestandardlistid="1944" />
                <TIMESTANDARDREF timestandardlistid="1950" />
                <TIMESTANDARDREF timestandardlistid="1956" />
                <TIMESTANDARDREF timestandardlistid="1962" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1092" daytime="14:51" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7602" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7603" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7604" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7605" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7606" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7607" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4082" />
                    <RANKING order="2" place="2" resultid="3284" />
                    <RANKING order="3" place="3" resultid="5663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7608" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3444" />
                    <RANKING order="2" place="2" resultid="6484" />
                    <RANKING order="3" place="3" resultid="4822" />
                    <RANKING order="4" place="4" resultid="2308" />
                    <RANKING order="5" place="5" resultid="2262" />
                    <RANKING order="6" place="6" resultid="5290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7609" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4222" />
                    <RANKING order="2" place="2" resultid="2798" />
                    <RANKING order="3" place="3" resultid="5125" />
                    <RANKING order="4" place="4" resultid="5972" />
                    <RANKING order="5" place="5" resultid="4074" />
                    <RANKING order="6" place="6" resultid="4788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7610" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2938" />
                    <RANKING order="2" place="2" resultid="2369" />
                    <RANKING order="3" place="3" resultid="6239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7611" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3161" />
                    <RANKING order="2" place="2" resultid="5501" />
                    <RANKING order="3" place="3" resultid="4320" />
                    <RANKING order="4" place="4" resultid="2080" />
                    <RANKING order="5" place="5" resultid="5114" />
                    <RANKING order="6" place="6" resultid="6209" />
                    <RANKING order="7" place="7" resultid="5887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7612" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2481" />
                    <RANKING order="2" place="2" resultid="3167" />
                    <RANKING order="3" place="3" resultid="4495" />
                    <RANKING order="4" place="4" resultid="3665" />
                    <RANKING order="5" place="5" resultid="5509" />
                    <RANKING order="6" place="6" resultid="4432" />
                    <RANKING order="7" place="7" resultid="4975" />
                    <RANKING order="8" place="-1" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7613" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2440" />
                    <RANKING order="2" place="2" resultid="2822" />
                    <RANKING order="3" place="3" resultid="4951" />
                    <RANKING order="4" place="4" resultid="4483" />
                    <RANKING order="5" place="5" resultid="3708" />
                    <RANKING order="6" place="-1" resultid="2862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7614" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4038" />
                    <RANKING order="2" place="2" resultid="3878" />
                    <RANKING order="3" place="3" resultid="6154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7615" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2035" />
                    <RANKING order="2" place="2" resultid="3869" />
                    <RANKING order="3" place="3" resultid="4717" />
                    <RANKING order="4" place="4" resultid="4463" />
                    <RANKING order="5" place="-1" resultid="2912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7616" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5981" />
                    <RANKING order="2" place="2" resultid="2619" />
                    <RANKING order="3" place="3" resultid="3834" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7271" daytime="14:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7272" daytime="14:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7273" daytime="15:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7274" daytime="15:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7275" daytime="15:09" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" daytime="18:37" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7662" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7663" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7664" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7665" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7666" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7667" agemax="69" agemin="65" name="I" />
                <AGEGROUP agegroupid="7668" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3445" />
                    <RANKING order="2" place="2" resultid="3908" />
                    <RANKING order="3" place="3" resultid="5291" />
                    <RANKING order="4" place="4" resultid="2263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7669" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5126" />
                    <RANKING order="2" place="2" resultid="5973" />
                    <RANKING order="3" place="3" resultid="4789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7670" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6240" />
                    <RANKING order="2" place="2" resultid="3406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7671" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6445" />
                    <RANKING order="2" place="2" resultid="3917" />
                    <RANKING order="3" place="3" resultid="6395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7672" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7673" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3709" />
                    <RANKING order="2" place="2" resultid="2395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7674" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6155" />
                    <RANKING order="2" place="2" resultid="5134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7675" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7676" agemax="24" agemin="20" name="0" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7300" daytime="18:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7301" daytime="19:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1886" />
                <TIMESTANDARDREF timestandardlistid="1892" />
                <TIMESTANDARDREF timestandardlistid="1898" />
                <TIMESTANDARDREF timestandardlistid="1904" />
                <TIMESTANDARDREF timestandardlistid="1910" />
                <TIMESTANDARDREF timestandardlistid="1916" />
                <TIMESTANDARDREF timestandardlistid="1922" />
                <TIMESTANDARDREF timestandardlistid="1928" />
                <TIMESTANDARDREF timestandardlistid="1934" />
                <TIMESTANDARDREF timestandardlistid="1940" />
                <TIMESTANDARDREF timestandardlistid="1946" />
                <TIMESTANDARDREF timestandardlistid="1952" />
                <TIMESTANDARDREF timestandardlistid="1958" />
                <TIMESTANDARDREF timestandardlistid="1847" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1108" daytime="15:13" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7617" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7618" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7619" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7620" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5685" />
                    <RANKING order="2" place="2" resultid="2635" />
                    <RANKING order="3" place="-1" resultid="2693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7621" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2200" />
                    <RANKING order="2" place="2" resultid="3126" />
                    <RANKING order="3" place="3" resultid="5164" />
                    <RANKING order="4" place="4" resultid="2419" />
                    <RANKING order="5" place="5" resultid="3932" />
                    <RANKING order="6" place="6" resultid="2684" />
                    <RANKING order="7" place="7" resultid="2728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7622" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4598" />
                    <RANKING order="2" place="2" resultid="5103" />
                    <RANKING order="3" place="3" resultid="4724" />
                    <RANKING order="4" place="4" resultid="2560" />
                    <RANKING order="5" place="5" resultid="2709" />
                    <RANKING order="6" place="6" resultid="2299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7623" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5281" />
                    <RANKING order="2" place="2" resultid="3185" />
                    <RANKING order="3" place="3" resultid="2116" />
                    <RANKING order="4" place="4" resultid="5693" />
                    <RANKING order="5" place="5" resultid="2836" />
                    <RANKING order="6" place="6" resultid="4603" />
                    <RANKING order="7" place="7" resultid="4156" />
                    <RANKING order="8" place="8" resultid="2603" />
                    <RANKING order="9" place="9" resultid="2749" />
                    <RANKING order="10" place="10" resultid="2757" />
                    <RANKING order="11" place="11" resultid="3240" />
                    <RANKING order="12" place="12" resultid="3148" />
                    <RANKING order="13" place="-1" resultid="3211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7624" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3853" />
                    <RANKING order="2" place="2" resultid="4616" />
                    <RANKING order="3" place="3" resultid="2430" />
                    <RANKING order="4" place="4" resultid="5593" />
                    <RANKING order="5" place="5" resultid="6030" />
                    <RANKING order="6" place="-1" resultid="2566" />
                    <RANKING order="7" place="-1" resultid="5728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7625" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5636" />
                    <RANKING order="2" place="2" resultid="4579" />
                    <RANKING order="3" place="3" resultid="2803" />
                    <RANKING order="4" place="4" resultid="2385" />
                    <RANKING order="5" place="5" resultid="5817" />
                    <RANKING order="6" place="6" resultid="6122" />
                    <RANKING order="7" place="7" resultid="2719" />
                    <RANKING order="8" place="8" resultid="2231" />
                    <RANKING order="9" place="-1" resultid="2277" />
                    <RANKING order="10" place="-1" resultid="5618" />
                    <RANKING order="11" place="-1" resultid="6469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7626" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="2360" />
                    <RANKING order="3" place="3" resultid="3659" />
                    <RANKING order="4" place="4" resultid="3741" />
                    <RANKING order="5" place="5" resultid="2667" />
                    <RANKING order="6" place="6" resultid="4363" />
                    <RANKING order="7" place="7" resultid="3683" />
                    <RANKING order="8" place="8" resultid="5827" />
                    <RANKING order="9" place="-1" resultid="5074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7627" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6043" />
                    <RANKING order="2" place="2" resultid="2043" />
                    <RANKING order="3" place="3" resultid="3200" />
                    <RANKING order="4" place="4" resultid="2054" />
                    <RANKING order="5" place="5" resultid="5627" />
                    <RANKING order="6" place="6" resultid="3527" />
                    <RANKING order="7" place="-1" resultid="2999" />
                    <RANKING order="8" place="-1" resultid="5023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7628" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3718" />
                    <RANKING order="2" place="2" resultid="6015" />
                    <RANKING order="3" place="3" resultid="6091" />
                    <RANKING order="4" place="4" resultid="4176" />
                    <RANKING order="5" place="5" resultid="5585" />
                    <RANKING order="6" place="6" resultid="4966" />
                    <RANKING order="7" place="-1" resultid="2446" />
                    <RANKING order="8" place="-1" resultid="5032" />
                    <RANKING order="9" place="-1" resultid="6218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7629" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3225" />
                    <RANKING order="2" place="2" resultid="4396" />
                    <RANKING order="3" place="3" resultid="2854" />
                    <RANKING order="4" place="4" resultid="3495" />
                    <RANKING order="5" place="5" resultid="3861" />
                    <RANKING order="6" place="6" resultid="3488" />
                    <RANKING order="7" place="7" resultid="5912" />
                    <RANKING order="8" place="-1" resultid="5249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7630" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6172" />
                    <RANKING order="2" place="2" resultid="5146" />
                    <RANKING order="3" place="3" resultid="2517" />
                    <RANKING order="4" place="4" resultid="2281" />
                    <RANKING order="5" place="5" resultid="6254" />
                    <RANKING order="6" place="-1" resultid="3453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7631" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2628" />
                    <RANKING order="2" place="2" resultid="2610" />
                    <RANKING order="3" place="3" resultid="3843" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7276" daytime="15:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7277" daytime="15:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7278" daytime="15:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7279" daytime="15:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7280" daytime="15:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7281" daytime="15:39" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7282" daytime="15:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7283" daytime="15:46" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7284" daytime="15:49" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7285" daytime="15:52" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="16:10" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7632" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7633" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7634" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7635" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7636" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4122" />
                    <RANKING order="2" place="2" resultid="4739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7637" agemax="69" agemin="65" name="I" />
                <AGEGROUP agegroupid="7638" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7639" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4771" />
                    <RANKING order="2" place="2" resultid="4229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7640" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2554" />
                    <RANKING order="2" place="2" resultid="5952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7641" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3800" />
                    <RANKING order="2" place="2" resultid="5502" />
                    <RANKING order="3" place="3" resultid="4321" />
                    <RANKING order="4" place="4" resultid="5888" />
                    <RANKING order="5" place="5" resultid="6210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7642" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5557" />
                    <RANKING order="2" place="2" resultid="3072" />
                    <RANKING order="3" place="3" resultid="6164" />
                    <RANKING order="4" place="4" resultid="4976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7643" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4484" />
                    <RANKING order="2" place="2" resultid="5601" />
                    <RANKING order="3" place="3" resultid="4024" />
                    <RANKING order="4" place="4" resultid="4013" />
                    <RANKING order="5" place="5" resultid="6355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7644" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2831" />
                    <RANKING order="2" place="2" resultid="5576" />
                    <RANKING order="3" place="3" resultid="5869" />
                    <RANKING order="4" place="4" resultid="4474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7645" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6129" />
                    <RANKING order="2" place="2" resultid="5837" />
                    <RANKING order="3" place="3" resultid="3329" />
                    <RANKING order="4" place="-1" resultid="3024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7646" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5982" />
                    <RANKING order="2" place="2" resultid="2771" />
                    <RANKING order="3" place="-1" resultid="4016" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7290" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7291" daytime="16:23" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7292" daytime="16:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7293" daytime="16:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1763" />
                <TIMESTANDARDREF timestandardlistid="1775" />
                <TIMESTANDARDREF timestandardlistid="1781" />
                <TIMESTANDARDREF timestandardlistid="1787" />
                <TIMESTANDARDREF timestandardlistid="1793" />
                <TIMESTANDARDREF timestandardlistid="1799" />
                <TIMESTANDARDREF timestandardlistid="1805" />
                <TIMESTANDARDREF timestandardlistid="1811" />
                <TIMESTANDARDREF timestandardlistid="1817" />
                <TIMESTANDARDREF timestandardlistid="1823" />
                <TIMESTANDARDREF timestandardlistid="1829" />
                <TIMESTANDARDREF timestandardlistid="1835" />
                <TIMESTANDARDREF timestandardlistid="1841" />
                <TIMESTANDARDREF timestandardlistid="1847" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1124" daytime="15:56" gender="X" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3819" />
                    <RANKING order="2" place="2" resultid="4137" />
                    <RANKING order="3" place="3" resultid="2325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="4139" />
                    <RANKING order="3" place="3" resultid="4182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3314" />
                    <RANKING order="2" place="2" resultid="6869" />
                    <RANKING order="3" place="3" resultid="4850" />
                    <RANKING order="4" place="4" resultid="6065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5059" />
                    <RANKING order="2" place="2" resultid="4752" />
                    <RANKING order="3" place="3" resultid="2832" />
                    <RANKING order="4" place="4" resultid="6262" />
                    <RANKING order="5" place="5" resultid="3697" />
                    <RANKING order="6" place="6" resultid="3312" />
                    <RANKING order="7" place="7" resultid="5058" />
                    <RANKING order="8" place="8" resultid="6409" />
                    <RANKING order="9" place="9" resultid="4454" />
                    <RANKING order="10" place="10" resultid="4544" />
                    <RANKING order="11" place="11" resultid="4031" />
                    <RANKING order="12" place="12" resultid="5154" />
                    <RANKING order="13" place="-1" resultid="3034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="5276" />
                    <RANKING order="3" place="3" resultid="5153" />
                    <RANKING order="4" place="4" resultid="5057" />
                    <RANKING order="5" place="5" resultid="6263" />
                    <RANKING order="6" place="6" resultid="4347" />
                    <RANKING order="7" place="7" resultid="3595" />
                    <RANKING order="8" place="-1" resultid="5654" />
                    <RANKING order="9" place="-1" resultid="6877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6261" />
                    <RANKING order="2" place="2" resultid="3593" />
                    <RANKING order="3" place="3" resultid="3594" />
                    <RANKING order="4" place="4" resultid="2875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="99" agemin="80" name="0" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7286" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7287" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7288" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7289" daytime="16:07" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-11-16" daytime="09:00" endtime="13:56" name="Zimowe Mistrzostwa Polskiw Pływaniu Masters BLOK II" number="2" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1288" daytime="11:02" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7767" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7768" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7769" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7770" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4650" />
                    <RANKING order="2" place="2" resultid="4171" />
                    <RANKING order="3" place="3" resultid="3942" />
                    <RANKING order="4" place="4" resultid="4816" />
                    <RANKING order="5" place="5" resultid="2703" />
                    <RANKING order="6" place="-1" resultid="5175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7771" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4781" />
                    <RANKING order="2" place="2" resultid="3795" />
                    <RANKING order="3" place="3" resultid="2098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7772" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4599" />
                    <RANKING order="2" place="2" resultid="2128" />
                    <RANKING order="3" place="3" resultid="2090" />
                    <RANKING order="4" place="4" resultid="3926" />
                    <RANKING order="5" place="5" resultid="3137" />
                    <RANKING order="6" place="6" resultid="5934" />
                    <RANKING order="7" place="7" resultid="2104" />
                    <RANKING order="8" place="8" resultid="2301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7773" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3214" />
                    <RANKING order="2" place="2" resultid="3260" />
                    <RANKING order="3" place="3" resultid="3766" />
                    <RANKING order="4" place="4" resultid="6501" />
                    <RANKING order="5" place="5" resultid="4158" />
                    <RANKING order="6" place="6" resultid="5863" />
                    <RANKING order="7" place="7" resultid="4654" />
                    <RANKING order="8" place="8" resultid="3241" />
                    <RANKING order="9" place="9" resultid="4845" />
                    <RANKING order="10" place="10" resultid="3149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7774" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4617" />
                    <RANKING order="2" place="2" resultid="6001" />
                    <RANKING order="3" place="3" resultid="5183" />
                    <RANKING order="4" place="4" resultid="2431" />
                    <RANKING order="5" place="5" resultid="5730" />
                    <RANKING order="6" place="6" resultid="6117" />
                    <RANKING order="7" place="7" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7775" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6305" />
                    <RANKING order="2" place="2" resultid="5637" />
                    <RANKING order="3" place="3" resultid="5754" />
                    <RANKING order="4" place="4" resultid="5522" />
                    <RANKING order="5" place="5" resultid="5819" />
                    <RANKING order="6" place="6" resultid="2720" />
                    <RANKING order="7" place="7" resultid="6123" />
                    <RANKING order="8" place="8" resultid="4519" />
                    <RANKING order="9" place="9" resultid="3656" />
                    <RANKING order="10" place="10" resultid="2232" />
                    <RANKING order="11" place="11" resultid="4298" />
                    <RANKING order="12" place="-1" resultid="2166" />
                    <RANKING order="13" place="-1" resultid="2292" />
                    <RANKING order="14" place="-1" resultid="2525" />
                    <RANKING order="15" place="-1" resultid="5084" />
                    <RANKING order="16" place="-1" resultid="5619" />
                    <RANKING order="17" place="-1" resultid="6470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7776" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4559" />
                    <RANKING order="2" place="2" resultid="2361" />
                    <RANKING order="3" place="3" resultid="6147" />
                    <RANKING order="4" place="4" resultid="4255" />
                    <RANKING order="5" place="5" resultid="4248" />
                    <RANKING order="6" place="6" resultid="3684" />
                    <RANKING order="7" place="7" resultid="3398" />
                    <RANKING order="8" place="8" resultid="3757" />
                    <RANKING order="9" place="9" resultid="3325" />
                    <RANKING order="10" place="10" resultid="6195" />
                    <RANKING order="11" place="11" resultid="5705" />
                    <RANKING order="12" place="12" resultid="3675" />
                    <RANKING order="13" place="13" resultid="2530" />
                    <RANKING order="14" place="14" resultid="3132" />
                    <RANKING order="15" place="15" resultid="4528" />
                    <RANKING order="16" place="16" resultid="3616" />
                    <RANKING order="17" place="17" resultid="6109" />
                    <RANKING order="18" place="18" resultid="5723" />
                    <RANKING order="19" place="19" resultid="5928" />
                    <RANKING order="20" place="20" resultid="5196" />
                    <RANKING order="21" place="21" resultid="3059" />
                    <RANKING order="22" place="22" resultid="4306" />
                    <RANKING order="23" place="23" resultid="5201" />
                    <RANKING order="24" place="24" resultid="4426" />
                    <RANKING order="25" place="25" resultid="3995" />
                    <RANKING order="26" place="-1" resultid="4387" />
                    <RANKING order="27" place="-1" resultid="5770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7777" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4929" />
                    <RANKING order="2" place="2" resultid="6045" />
                    <RANKING order="3" place="3" resultid="6007" />
                    <RANKING order="4" place="4" resultid="4695" />
                    <RANKING order="5" place="5" resultid="4625" />
                    <RANKING order="6" place="6" resultid="5715" />
                    <RANKING order="7" place="7" resultid="6139" />
                    <RANKING order="8" place="8" resultid="3020" />
                    <RANKING order="9" place="9" resultid="4708" />
                    <RANKING order="10" place="10" resultid="5008" />
                    <RANKING order="11" place="11" resultid="4315" />
                    <RANKING order="12" place="12" resultid="2009" />
                    <RANKING order="13" place="13" resultid="5097" />
                    <RANKING order="14" place="14" resultid="6188" />
                    <RANKING order="15" place="15" resultid="3421" />
                    <RANKING order="16" place="16" resultid="3047" />
                    <RANKING order="17" place="17" resultid="4882" />
                    <RANKING order="18" place="18" resultid="4909" />
                    <RANKING order="19" place="19" resultid="2067" />
                    <RANKING order="20" place="20" resultid="2491" />
                    <RANKING order="21" place="21" resultid="5255" />
                    <RANKING order="22" place="22" resultid="2739" />
                    <RANKING order="23" place="-1" resultid="2030" />
                    <RANKING order="24" place="-1" resultid="2111" />
                    <RANKING order="25" place="-1" resultid="4960" />
                    <RANKING order="26" place="-1" resultid="5025" />
                    <RANKING order="27" place="-1" resultid="6378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7778" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6017" />
                    <RANKING order="2" place="2" resultid="2965" />
                    <RANKING order="3" place="3" resultid="4422" />
                    <RANKING order="4" place="4" resultid="4588" />
                    <RANKING order="5" place="5" resultid="2379" />
                    <RANKING order="6" place="6" resultid="5205" />
                    <RANKING order="7" place="7" resultid="6182" />
                    <RANKING order="8" place="8" resultid="3430" />
                    <RANKING order="9" place="9" resultid="4682" />
                    <RANKING order="10" place="10" resultid="5215" />
                    <RANKING order="11" place="11" resultid="5221" />
                    <RANKING order="12" place="12" resultid="5788" />
                    <RANKING order="13" place="13" resultid="2543" />
                    <RANKING order="14" place="14" resultid="4887" />
                    <RANKING order="15" place="15" resultid="5237" />
                    <RANKING order="16" place="16" resultid="4504" />
                    <RANKING order="17" place="17" resultid="2448" />
                    <RANKING order="18" place="18" resultid="3549" />
                    <RANKING order="19" place="19" resultid="6864" />
                    <RANKING order="20" place="-1" resultid="2025" />
                    <RANKING order="21" place="-1" resultid="4346" />
                    <RANKING order="22" place="-1" resultid="4330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7779" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4891" />
                    <RANKING order="2" place="2" resultid="2131" />
                    <RANKING order="3" place="3" resultid="2855" />
                    <RANKING order="4" place="4" resultid="3489" />
                    <RANKING order="5" place="5" resultid="2976" />
                    <RANKING order="6" place="6" resultid="4397" />
                    <RANKING order="7" place="7" resultid="3226" />
                    <RANKING order="8" place="8" resultid="4748" />
                    <RANKING order="9" place="9" resultid="2952" />
                    <RANKING order="10" place="10" resultid="3863" />
                    <RANKING order="11" place="11" resultid="6433" />
                    <RANKING order="12" place="12" resultid="6367" />
                    <RANKING order="13" place="13" resultid="4676" />
                    <RANKING order="14" place="14" resultid="6235" />
                    <RANKING order="15" place="15" resultid="4668" />
                    <RANKING order="16" place="16" resultid="2151" />
                    <RANKING order="17" place="17" resultid="5914" />
                    <RANKING order="18" place="18" resultid="3426" />
                    <RANKING order="19" place="19" resultid="2846" />
                    <RANKING order="20" place="-1" resultid="3267" />
                    <RANKING order="21" place="-1" resultid="3435" />
                    <RANKING order="22" place="-1" resultid="3543" />
                    <RANKING order="23" place="-1" resultid="3547" />
                    <RANKING order="24" place="-1" resultid="4311" />
                    <RANKING order="25" place="-1" resultid="4470" />
                    <RANKING order="26" place="-1" resultid="4996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7780" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4896" />
                    <RANKING order="2" place="2" resultid="2147" />
                    <RANKING order="3" place="3" resultid="3728" />
                    <RANKING order="4" place="4" resultid="6872" />
                    <RANKING order="5" place="5" resultid="4632" />
                    <RANKING order="6" place="6" resultid="6053" />
                    <RANKING order="7" place="7" resultid="2580" />
                    <RANKING order="8" place="8" resultid="6256" />
                    <RANKING order="9" place="9" resultid="6351" />
                    <RANKING order="10" place="10" resultid="3509" />
                    <RANKING order="11" place="11" resultid="2176" />
                    <RANKING order="12" place="12" resultid="2908" />
                    <RANKING order="13" place="13" resultid="3016" />
                    <RANKING order="14" place="14" resultid="6440" />
                    <RANKING order="15" place="15" resultid="2514" />
                    <RANKING order="16" place="16" resultid="3474" />
                    <RANKING order="17" place="-1" resultid="2184" />
                    <RANKING order="18" place="-1" resultid="3582" />
                    <RANKING order="19" place="-1" resultid="5148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7781" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4186" />
                    <RANKING order="2" place="2" resultid="5189" />
                    <RANKING order="3" place="3" resultid="3823" />
                    <RANKING order="4" place="4" resultid="2611" />
                    <RANKING order="5" place="5" resultid="2319" />
                    <RANKING order="6" place="6" resultid="3845" />
                    <RANKING order="7" place="7" resultid="3478" />
                    <RANKING order="8" place="8" resultid="3894" />
                    <RANKING order="9" place="9" resultid="2660" />
                    <RANKING order="10" place="10" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7349" daytime="11:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7350" daytime="11:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7351" daytime="11:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7352" daytime="11:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7353" daytime="11:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7354" daytime="11:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7355" daytime="11:17" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7356" daytime="11:19" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7357" daytime="11:21" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7358" daytime="11:23" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7359" daytime="11:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7360" daytime="11:27" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7361" daytime="11:29" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7362" daytime="11:31" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7363" daytime="11:32" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7364" daytime="11:34" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7365" daytime="11:36" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7366" daytime="11:38" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7367" daytime="11:39" number="19" order="19" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1272" daytime="10:42" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7752" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7753" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7754" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7755" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7756" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7757" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5665" />
                    <RANKING order="2" place="2" resultid="5962" />
                    <RANKING order="3" place="3" resultid="2349" />
                    <RANKING order="4" place="4" resultid="4166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7758" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3086" />
                    <RANKING order="2" place="2" resultid="2471" />
                    <RANKING order="3" place="3" resultid="3809" />
                    <RANKING order="4" place="4" resultid="3910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7759" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4772" />
                    <RANKING order="2" place="2" resultid="5799" />
                    <RANKING order="3" place="3" resultid="4059" />
                    <RANKING order="4" place="4" resultid="4231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7760" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2555" />
                    <RANKING order="2" place="2" resultid="4269" />
                    <RANKING order="3" place="3" resultid="6242" />
                    <RANKING order="4" place="4" resultid="5954" />
                    <RANKING order="5" place="5" resultid="6203" />
                    <RANKING order="6" place="6" resultid="3972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7761" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5504" />
                    <RANKING order="2" place="2" resultid="5805" />
                    <RANKING order="3" place="3" resultid="5089" />
                    <RANKING order="4" place="4" resultid="3918" />
                    <RANKING order="5" place="5" resultid="6211" />
                    <RANKING order="6" place="6" resultid="5889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7762" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3693" />
                    <RANKING order="2" place="2" resultid="5559" />
                    <RANKING order="3" place="3" resultid="2933" />
                    <RANKING order="4" place="4" resultid="5110" />
                    <RANKING order="5" place="5" resultid="4301" />
                    <RANKING order="6" place="6" resultid="5642" />
                    <RANKING order="7" place="7" resultid="4492" />
                    <RANKING order="8" place="-1" resultid="6411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7763" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2441" />
                    <RANKING order="2" place="2" resultid="2816" />
                    <RANKING order="3" place="3" resultid="4948" />
                    <RANKING order="4" place="4" resultid="4642" />
                    <RANKING order="5" place="5" resultid="6227" />
                    <RANKING order="6" place="6" resultid="4417" />
                    <RANKING order="7" place="7" resultid="6391" />
                    <RANKING order="8" place="8" resultid="5602" />
                    <RANKING order="9" place="9" resultid="2863" />
                    <RANKING order="10" place="10" resultid="5611" />
                    <RANKING order="11" place="11" resultid="2653" />
                    <RANKING order="12" place="-1" resultid="4335" />
                    <RANKING order="13" place="-1" resultid="5647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7764" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5809" />
                    <RANKING order="2" place="2" resultid="5243" />
                    <RANKING order="3" place="3" resultid="4039" />
                    <RANKING order="4" place="4" resultid="3703" />
                    <RANKING order="5" place="5" resultid="4743" />
                    <RANKING order="6" place="6" resultid="3749" />
                    <RANKING order="7" place="7" resultid="2828" />
                    <RANKING order="8" place="8" resultid="5578" />
                    <RANKING order="9" place="9" resultid="2646" />
                    <RANKING order="10" place="10" resultid="3470" />
                    <RANKING order="11" place="11" resultid="5020" />
                    <RANKING order="12" place="12" resultid="5870" />
                    <RANKING order="13" place="13" resultid="6460" />
                    <RANKING order="14" place="14" resultid="4475" />
                    <RANKING order="15" place="15" resultid="3505" />
                    <RANKING order="16" place="-1" resultid="4340" />
                    <RANKING order="17" place="-1" resultid="4539" />
                    <RANKING order="18" place="-1" resultid="4661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7765" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2775" />
                    <RANKING order="2" place="2" resultid="2981" />
                    <RANKING order="3" place="3" resultid="2036" />
                    <RANKING order="4" place="4" resultid="5838" />
                    <RANKING order="5" place="5" resultid="6336" />
                    <RANKING order="6" place="6" resultid="2142" />
                    <RANKING order="7" place="7" resultid="4442" />
                    <RANKING order="8" place="8" resultid="3331" />
                    <RANKING order="9" place="9" resultid="5267" />
                    <RANKING order="10" place="10" resultid="5843" />
                    <RANKING order="11" place="11" resultid="3484" />
                    <RANKING order="12" place="12" resultid="3295" />
                    <RANKING order="13" place="13" resultid="4445" />
                    <RANKING order="14" place="-1" resultid="2778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7766" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="3736" />
                    <RANKING order="3" place="3" resultid="2179" />
                    <RANKING order="4" place="4" resultid="3836" />
                    <RANKING order="5" place="5" resultid="2675" />
                    <RANKING order="6" place="6" resultid="3559" />
                    <RANKING order="7" place="7" resultid="3553" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7340" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7341" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7342" daytime="10:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7343" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7344" daytime="10:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7345" daytime="10:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7346" daytime="10:56" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7347" daytime="10:58" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7348" daytime="11:00" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="11:41" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7782" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7783" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7784" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7785" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7786" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7787" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3789" />
                    <RANKING order="2" place="2" resultid="4084" />
                    <RANKING order="3" place="3" resultid="2073" />
                    <RANKING order="4" place="-1" resultid="4091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7788" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3446" />
                    <RANKING order="2" place="2" resultid="6485" />
                    <RANKING order="3" place="3" resultid="4115" />
                    <RANKING order="4" place="4" resultid="4149" />
                    <RANKING order="5" place="5" resultid="2265" />
                    <RANKING order="6" place="6" resultid="2591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7789" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5672" />
                    <RANKING order="2" place="2" resultid="3105" />
                    <RANKING order="3" place="3" resultid="5128" />
                    <RANKING order="4" place="4" resultid="6330" />
                    <RANKING order="5" place="5" resultid="4791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7790" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3091" />
                    <RANKING order="2" place="2" resultid="3989" />
                    <RANKING order="3" place="3" resultid="2939" />
                    <RANKING order="4" place="4" resultid="2371" />
                    <RANKING order="5" place="5" resultid="3407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7791" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3156" />
                    <RANKING order="2" place="2" resultid="2082" />
                    <RANKING order="3" place="3" resultid="4323" />
                    <RANKING order="4" place="4" resultid="5491" />
                    <RANKING order="5" place="5" resultid="6212" />
                    <RANKING order="6" place="6" resultid="5890" />
                    <RANKING order="7" place="7" resultid="4374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7792" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2597" />
                    <RANKING order="2" place="2" resultid="4497" />
                    <RANKING order="3" place="3" resultid="3074" />
                    <RANKING order="4" place="4" resultid="3667" />
                    <RANKING order="5" place="5" resultid="4302" />
                    <RANKING order="6" place="6" resultid="4434" />
                    <RANKING order="7" place="7" resultid="5737" />
                    <RANKING order="8" place="8" resultid="5263" />
                    <RANKING order="9" place="9" resultid="3277" />
                    <RANKING order="10" place="-1" resultid="3958" />
                    <RANKING order="11" place="-1" resultid="6166" />
                    <RANKING order="12" place="-1" resultid="6412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7793" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3381" />
                    <RANKING order="2" place="2" resultid="2821" />
                    <RANKING order="3" place="3" resultid="4953" />
                    <RANKING order="4" place="4" resultid="4486" />
                    <RANKING order="5" place="5" resultid="4643" />
                    <RANKING order="6" place="6" resultid="2487" />
                    <RANKING order="7" place="7" resultid="2864" />
                    <RANKING order="8" place="8" resultid="2396" />
                    <RANKING order="9" place="9" resultid="3387" />
                    <RANKING order="10" place="-1" resultid="4026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7794" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5244" />
                    <RANKING order="2" place="2" resultid="3522" />
                    <RANKING order="3" place="3" resultid="4040" />
                    <RANKING order="4" place="4" resultid="3880" />
                    <RANKING order="5" place="5" resultid="6456" />
                    <RANKING order="6" place="6" resultid="5135" />
                    <RANKING order="7" place="7" resultid="4610" />
                    <RANKING order="8" place="8" resultid="5021" />
                    <RANKING order="9" place="9" resultid="6461" />
                    <RANKING order="10" place="10" resultid="3392" />
                    <RANKING order="11" place="11" resultid="4476" />
                    <RANKING order="12" place="-1" resultid="3004" />
                    <RANKING order="13" place="-1" resultid="3113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7795" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2037" />
                    <RANKING order="2" place="2" resultid="2785" />
                    <RANKING order="3" place="3" resultid="3871" />
                    <RANKING order="4" place="4" resultid="6337" />
                    <RANKING order="5" place="5" resultid="4525" />
                    <RANKING order="6" place="6" resultid="4687" />
                    <RANKING order="7" place="7" resultid="3465" />
                    <RANKING order="8" place="8" resultid="4719" />
                    <RANKING order="9" place="9" resultid="5121" />
                    <RANKING order="10" place="10" resultid="4446" />
                    <RANKING order="11" place="11" resultid="4380" />
                    <RANKING order="12" place="-1" resultid="2914" />
                    <RANKING order="13" place="-1" resultid="4465" />
                    <RANKING order="14" place="-1" resultid="6453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7796" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5984" />
                    <RANKING order="2" place="2" resultid="2621" />
                    <RANKING order="3" place="3" resultid="3556" />
                    <RANKING order="4" place="4" resultid="4018" />
                    <RANKING order="5" place="5" resultid="3837" />
                    <RANKING order="6" place="6" resultid="5299" />
                    <RANKING order="7" place="7" resultid="2676" />
                    <RANKING order="8" place="8" resultid="3539" />
                    <RANKING order="9" place="9" resultid="3562" />
                    <RANKING order="10" place="-1" resultid="4193" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7368" daytime="11:41" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7369" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7370" daytime="11:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7371" daytime="11:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7372" daytime="11:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7373" daytime="11:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7374" daytime="11:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7375" daytime="12:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7376" daytime="12:02" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1240" daytime="09:39" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7722" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7723" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7724" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7725" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7726" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7727" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5961" />
                    <RANKING order="2" place="2" resultid="4083" />
                    <RANKING order="3" place="3" resultid="2348" />
                    <RANKING order="4" place="4" resultid="3773" />
                    <RANKING order="5" place="5" resultid="2072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7728" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4148" />
                    <RANKING order="2" place="2" resultid="2264" />
                    <RANKING order="3" place="3" resultid="5292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7729" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5671" />
                    <RANKING order="2" place="2" resultid="4224" />
                    <RANKING order="3" place="3" resultid="2794" />
                    <RANKING order="4" place="4" resultid="5548" />
                    <RANKING order="5" place="5" resultid="6329" />
                    <RANKING order="6" place="6" resultid="5974" />
                    <RANKING order="7" place="-1" resultid="4076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7730" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                    <RANKING order="2" place="2" resultid="2943" />
                    <RANKING order="3" place="3" resultid="2370" />
                    <RANKING order="4" place="4" resultid="6241" />
                    <RANKING order="5" place="5" resultid="3971" />
                    <RANKING order="6" place="-1" resultid="2271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7731" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3801" />
                    <RANKING order="2" place="2" resultid="4322" />
                    <RANKING order="3" place="3" resultid="4702" />
                    <RANKING order="4" place="4" resultid="6446" />
                    <RANKING order="5" place="5" resultid="6301" />
                    <RANKING order="6" place="6" resultid="3570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7732" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5510" />
                    <RANKING order="2" place="2" resultid="3666" />
                    <RANKING order="3" place="3" resultid="4977" />
                    <RANKING order="4" place="4" resultid="4900" />
                    <RANKING order="5" place="5" resultid="5948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7733" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3710" />
                    <RANKING order="2" place="2" resultid="2656" />
                    <RANKING order="3" place="3" resultid="4593" />
                    <RANKING order="4" place="4" resultid="4025" />
                    <RANKING order="5" place="5" resultid="5610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7734" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4742" />
                    <RANKING order="2" place="2" resultid="3702" />
                    <RANKING order="3" place="3" resultid="3879" />
                    <RANKING order="4" place="4" resultid="4609" />
                    <RANKING order="5" place="5" resultid="5536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7735" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4378" />
                    <RANKING order="2" place="-1" resultid="3025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7736" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5983" />
                    <RANKING order="2" place="2" resultid="3835" />
                    <RANKING order="3" place="3" resultid="5905" />
                    <RANKING order="4" place="4" resultid="4215" />
                    <RANKING order="5" place="5" resultid="5298" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7327" daytime="09:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7328" daytime="09:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7329" daytime="09:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7330" daytime="09:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7331" daytime="10:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1368" daytime="13:16" gender="F" number="20" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7842" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7843" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4141" />
                    <RANKING order="2" place="-1" resultid="3816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7844" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7845" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3316" />
                    <RANKING order="2" place="2" resultid="2948" />
                    <RANKING order="3" place="3" resultid="5155" />
                    <RANKING order="4" place="4" resultid="6406" />
                    <RANKING order="5" place="5" resultid="4033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7846" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4546" />
                    <RANKING order="2" place="2" resultid="4761" />
                    <RANKING order="3" place="3" resultid="6264" />
                    <RANKING order="4" place="4" resultid="5061" />
                    <RANKING order="5" place="5" resultid="3319" />
                    <RANKING order="6" place="-1" resultid="4348" />
                    <RANKING order="7" place="-1" resultid="3030" />
                    <RANKING order="8" place="-1" resultid="5655" />
                    <RANKING order="9" place="-1" resultid="6476" />
                    <RANKING order="10" place="-1" resultid="5517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7847" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2789" />
                    <RANKING order="2" place="2" resultid="4455" />
                    <RANKING order="3" place="3" resultid="3596" />
                    <RANKING order="4" place="-1" resultid="3597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7848" agemax="99" agemin="80" name="0" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7399" daytime="13:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7400" daytime="13:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7401" daytime="13:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="09:17" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7707" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7708" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2243" />
                    <RANKING order="2" place="-1" resultid="2891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7709" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7710" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5686" />
                    <RANKING order="2" place="2" resultid="4649" />
                    <RANKING order="3" place="3" resultid="3941" />
                    <RANKING order="4" place="4" resultid="2506" />
                    <RANKING order="5" place="5" resultid="2702" />
                    <RANKING order="6" place="-1" resultid="5174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7711" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3783" />
                    <RANKING order="2" place="2" resultid="2455" />
                    <RANKING order="3" place="3" resultid="3947" />
                    <RANKING order="4" place="4" resultid="4066" />
                    <RANKING order="5" place="5" resultid="3933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7712" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2126" />
                    <RANKING order="2" place="2" resultid="5778" />
                    <RANKING order="3" place="3" resultid="2711" />
                    <RANKING order="4" place="4" resultid="2300" />
                    <RANKING order="5" place="5" resultid="3208" />
                    <RANKING order="6" place="6" resultid="3248" />
                    <RANKING order="7" place="-1" resultid="3650" />
                    <RANKING order="8" place="-1" resultid="5678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7713" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3213" />
                    <RANKING order="2" place="2" resultid="3765" />
                    <RANKING order="3" place="3" resultid="2838" />
                    <RANKING order="4" place="4" resultid="5695" />
                    <RANKING order="5" place="5" resultid="4157" />
                    <RANKING order="6" place="6" resultid="2750" />
                    <RANKING order="7" place="7" resultid="2758" />
                    <RANKING order="8" place="8" resultid="4844" />
                    <RANKING order="9" place="-1" resultid="4356" />
                    <RANKING order="10" place="-1" resultid="5813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7714" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3854" />
                    <RANKING order="2" place="2" resultid="2412" />
                    <RANKING order="3" place="3" resultid="4798" />
                    <RANKING order="4" place="4" resultid="5729" />
                    <RANKING order="5" place="5" resultid="2344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7715" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4922" />
                    <RANKING order="2" place="2" resultid="5992" />
                    <RANKING order="3" place="3" resultid="3081" />
                    <RANKING order="4" place="4" resultid="4580" />
                    <RANKING order="5" place="5" resultid="2800" />
                    <RANKING order="6" place="6" resultid="2463" />
                    <RANKING order="7" place="7" resultid="4275" />
                    <RANKING order="8" place="8" resultid="4297" />
                    <RANKING order="9" place="9" resultid="5083" />
                    <RANKING order="10" place="10" resultid="3964" />
                    <RANKING order="11" place="11" resultid="5140" />
                    <RANKING order="12" place="-1" resultid="3627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7716" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3742" />
                    <RANKING order="2" place="2" resultid="2668" />
                    <RANKING order="3" place="3" resultid="4386" />
                    <RANKING order="4" place="4" resultid="6345" />
                    <RANKING order="5" place="5" resultid="5882" />
                    <RANKING order="6" place="6" resultid="3634" />
                    <RANKING order="7" place="7" resultid="6194" />
                    <RANKING order="8" place="8" resultid="5076" />
                    <RANKING order="9" place="9" resultid="3756" />
                    <RANKING order="10" place="10" resultid="3615" />
                    <RANKING order="11" place="11" resultid="5704" />
                    <RANKING order="12" place="12" resultid="6108" />
                    <RANKING order="13" place="13" resultid="5195" />
                    <RANKING order="14" place="14" resultid="5828" />
                    <RANKING order="15" place="-1" resultid="5769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7717" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2994" />
                    <RANKING order="2" place="2" resultid="6044" />
                    <RANKING order="3" place="3" resultid="6372" />
                    <RANKING order="4" place="4" resultid="6138" />
                    <RANKING order="5" place="5" resultid="2900" />
                    <RANKING order="6" place="6" resultid="3053" />
                    <RANKING order="7" place="7" resultid="2055" />
                    <RANKING order="8" place="8" resultid="5014" />
                    <RANKING order="9" place="9" resultid="3043" />
                    <RANKING order="10" place="10" resultid="4694" />
                    <RANKING order="11" place="11" resultid="5039" />
                    <RANKING order="12" place="12" resultid="3620" />
                    <RANKING order="13" place="13" resultid="4831" />
                    <RANKING order="14" place="14" resultid="2255" />
                    <RANKING order="15" place="-1" resultid="2738" />
                    <RANKING order="16" place="-1" resultid="4707" />
                    <RANKING order="17" place="-1" resultid="5007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7718" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4732" />
                    <RANKING order="2" place="2" resultid="3719" />
                    <RANKING order="3" place="3" resultid="3193" />
                    <RANKING order="4" place="4" resultid="4587" />
                    <RANKING order="5" place="5" resultid="4177" />
                    <RANKING order="6" place="6" resultid="5220" />
                    <RANKING order="7" place="7" resultid="5004" />
                    <RANKING order="8" place="8" resultid="2542" />
                    <RANKING order="9" place="-1" resultid="3886" />
                    <RANKING order="10" place="-1" resultid="5236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7719" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4242" />
                    <RANKING order="2" place="2" resultid="5857" />
                    <RANKING order="3" place="3" resultid="4747" />
                    <RANKING order="4" place="4" resultid="4713" />
                    <RANKING order="5" place="5" resultid="4667" />
                    <RANKING order="6" place="6" resultid="3497" />
                    <RANKING order="7" place="7" resultid="3862" />
                    <RANKING order="8" place="8" resultid="6234" />
                    <RANKING order="9" place="-1" resultid="3266" />
                    <RANKING order="10" place="-1" resultid="4675" />
                    <RANKING order="11" place="-1" resultid="4995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7720" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5231" />
                    <RANKING order="2" place="2" resultid="2282" />
                    <RANKING order="3" place="3" resultid="6052" />
                    <RANKING order="4" place="4" resultid="5897" />
                    <RANKING order="5" place="-1" resultid="2336" />
                    <RANKING order="6" place="-1" resultid="3454" />
                    <RANKING order="7" place="-1" resultid="8161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7721" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4201" />
                    <RANKING order="2" place="2" resultid="4208" />
                    <RANKING order="3" place="3" resultid="2318" />
                    <RANKING order="4" place="-1" resultid="2135" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7315" daytime="09:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7316" daytime="09:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7317" daytime="09:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7318" daytime="09:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7319" daytime="09:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7320" daytime="09:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7321" daytime="09:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7322" daytime="09:31" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7323" daytime="09:32" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7324" daytime="09:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7325" daytime="09:35" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7326" daytime="09:37" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1336" daytime="12:36" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7812" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7813" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7814" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7815" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7816" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7817" agemax="69" agemin="65" name="I" />
                <AGEGROUP agegroupid="7818" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4824" />
                    <RANKING order="2" place="2" resultid="5293" />
                    <RANKING order="3" place="3" resultid="2310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7819" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4773" />
                    <RANKING order="2" place="2" resultid="2797" />
                    <RANKING order="3" place="3" resultid="5975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7820" agemax="54" agemin="50" name="F" />
                <AGEGROUP agegroupid="7821" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3162" />
                    <RANKING order="2" place="2" resultid="5492" />
                    <RANKING order="3" place="3" resultid="6447" />
                    <RANKING order="4" place="4" resultid="5115" />
                    <RANKING order="5" place="5" resultid="6396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7822" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3168" />
                    <RANKING order="2" place="2" resultid="4978" />
                    <RANKING order="3" place="3" resultid="4901" />
                    <RANKING order="4" place="-1" resultid="5511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7823" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4939" />
                    <RANKING order="2" place="2" resultid="3711" />
                    <RANKING order="3" place="3" resultid="5603" />
                    <RANKING order="4" place="-1" resultid="6356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7824" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6157" />
                    <RANKING order="2" place="2" resultid="5871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7825" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7826" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4194" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7391" daytime="12:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7392" daytime="12:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7393" daytime="12:47" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1207" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7692" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7693" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7694" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7695" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3778" />
                    <RANKING order="2" place="2" resultid="4097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7696" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7697" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3788" />
                    <RANKING order="2" place="2" resultid="5664" />
                    <RANKING order="3" place="3" resultid="4131" />
                    <RANKING order="4" place="4" resultid="4165" />
                    <RANKING order="5" place="5" resultid="3772" />
                    <RANKING order="6" place="-1" resultid="4090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7698" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4823" />
                    <RANKING order="2" place="2" resultid="3808" />
                    <RANKING order="3" place="3" resultid="2309" />
                    <RANKING order="4" place="4" resultid="3909" />
                    <RANKING order="5" place="5" resultid="2590" />
                    <RANKING order="6" place="6" resultid="3982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7699" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3104" />
                    <RANKING order="2" place="2" resultid="4223" />
                    <RANKING order="3" place="3" resultid="5798" />
                    <RANKING order="4" place="4" resultid="4058" />
                    <RANKING order="5" place="5" resultid="5127" />
                    <RANKING order="6" place="6" resultid="4075" />
                    <RANKING order="7" place="7" resultid="4790" />
                    <RANKING order="8" place="8" resultid="4230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7700" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3988" />
                    <RANKING order="2" place="2" resultid="5953" />
                    <RANKING order="3" place="3" resultid="6202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7701" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3155" />
                    <RANKING order="2" place="2" resultid="5804" />
                    <RANKING order="3" place="3" resultid="2354" />
                    <RANKING order="4" place="4" resultid="5503" />
                    <RANKING order="5" place="5" resultid="2081" />
                    <RANKING order="6" place="6" resultid="4373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7702" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3174" />
                    <RANKING order="2" place="2" resultid="6165" />
                    <RANKING order="3" place="3" resultid="3073" />
                    <RANKING order="4" place="4" resultid="5558" />
                    <RANKING order="5" place="5" resultid="4496" />
                    <RANKING order="6" place="6" resultid="5109" />
                    <RANKING order="7" place="7" resultid="3692" />
                    <RANKING order="8" place="8" resultid="4433" />
                    <RANKING order="9" place="9" resultid="5736" />
                    <RANKING order="10" place="10" resultid="5262" />
                    <RANKING order="11" place="11" resultid="3276" />
                    <RANKING order="12" place="12" resultid="3957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7703" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3380" />
                    <RANKING order="2" place="2" resultid="4952" />
                    <RANKING order="3" place="3" resultid="4485" />
                    <RANKING order="4" place="4" resultid="5001" />
                    <RANKING order="5" place="5" resultid="2486" />
                    <RANKING order="6" place="6" resultid="6226" />
                    <RANKING order="7" place="7" resultid="4947" />
                    <RANKING order="8" place="8" resultid="4007" />
                    <RANKING order="9" place="-1" resultid="4334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7704" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3003" />
                    <RANKING order="2" place="2" resultid="3521" />
                    <RANKING order="3" place="3" resultid="6455" />
                    <RANKING order="4" place="4" resultid="2824" />
                    <RANKING order="5" place="5" resultid="5577" />
                    <RANKING order="6" place="6" resultid="6156" />
                    <RANKING order="7" place="7" resultid="3504" />
                    <RANKING order="8" place="8" resultid="5535" />
                    <RANKING order="9" place="-1" resultid="3516" />
                    <RANKING order="10" place="-1" resultid="4339" />
                    <RANKING order="11" place="-1" resultid="5210" />
                    <RANKING order="12" place="-1" resultid="3112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7705" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3870" />
                    <RANKING order="2" place="2" resultid="2781" />
                    <RANKING order="3" place="3" resultid="4524" />
                    <RANKING order="4" place="4" resultid="4686" />
                    <RANKING order="5" place="5" resultid="4464" />
                    <RANKING order="6" place="6" resultid="4718" />
                    <RANKING order="7" place="7" resultid="5120" />
                    <RANKING order="8" place="8" resultid="3294" />
                    <RANKING order="9" place="9" resultid="2745" />
                    <RANKING order="10" place="-1" resultid="2913" />
                    <RANKING order="11" place="-1" resultid="3330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7706" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4192" />
                    <RANKING order="2" place="2" resultid="3271" />
                    <RANKING order="3" place="3" resultid="2331" />
                    <RANKING order="4" place="4" resultid="4017" />
                    <RANKING order="5" place="5" resultid="3538" />
                    <RANKING order="6" place="6" resultid="5904" />
                    <RANKING order="7" place="-1" resultid="4214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7306" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7307" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7308" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7309" daytime="09:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7310" daytime="09:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7311" daytime="09:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7312" daytime="09:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7313" daytime="09:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7314" daytime="09:15" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1391" daytime="13:29" gender="M" number="21" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7849" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3304" />
                    <RANKING order="2" place="2" resultid="3952" />
                    <RANKING order="3" place="-1" resultid="4136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7850" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3306" />
                    <RANKING order="2" place="2" resultid="4853" />
                    <RANKING order="3" place="3" resultid="5760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7851" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4756" />
                    <RANKING order="2" place="2" resultid="5656" />
                    <RANKING order="3" place="3" resultid="6874" />
                    <RANKING order="4" place="4" resultid="6267" />
                    <RANKING order="5" place="5" resultid="2326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7852" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4279" />
                    <RANKING order="2" place="2" resultid="3037" />
                    <RANKING order="3" place="3" resultid="6058" />
                    <RANKING order="4" place="4" resultid="6875" />
                    <RANKING order="5" place="5" resultid="3308" />
                    <RANKING order="6" place="6" resultid="5067" />
                    <RANKING order="7" place="7" resultid="5156" />
                    <RANKING order="8" place="8" resultid="6063" />
                    <RANKING order="9" place="9" resultid="6266" />
                    <RANKING order="10" place="10" resultid="5068" />
                    <RANKING order="11" place="11" resultid="3069" />
                    <RANKING order="12" place="12" resultid="4758" />
                    <RANKING order="13" place="13" resultid="4548" />
                    <RANKING order="14" place="14" resultid="4351" />
                    <RANKING order="15" place="-1" resultid="3441" />
                    <RANKING order="16" place="-1" resultid="4352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7853" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6265" />
                    <RANKING order="2" place="2" resultid="4757" />
                    <RANKING order="3" place="3" resultid="4905" />
                    <RANKING order="4" place="4" resultid="3033" />
                    <RANKING order="5" place="5" resultid="4762" />
                    <RANKING order="6" place="6" resultid="5069" />
                    <RANKING order="7" place="7" resultid="5070" />
                    <RANKING order="8" place="8" resultid="5273" />
                    <RANKING order="9" place="9" resultid="4456" />
                    <RANKING order="10" place="-1" resultid="6876" />
                    <RANKING order="11" place="-1" resultid="3038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7854" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5272" />
                    <RANKING order="2" place="2" resultid="3599" />
                    <RANKING order="3" place="-1" resultid="3598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7855" agemax="99" agemin="80" name="0" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7402" daytime="13:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7403" daytime="13:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7404" daytime="13:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7405" daytime="13:41" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7406" daytime="13:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:05" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7737" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7738" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7739" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7740" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4635" />
                    <RANKING order="2" place="2" resultid="2637" />
                    <RANKING order="3" place="3" resultid="2694" />
                    <RANKING order="4" place="4" resultid="2507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7741" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3097" />
                    <RANKING order="2" place="2" resultid="2201" />
                    <RANKING order="3" place="3" resultid="5166" />
                    <RANKING order="4" place="4" resultid="2421" />
                    <RANKING order="5" place="5" resultid="3948" />
                    <RANKING order="6" place="6" resultid="2729" />
                    <RANKING order="7" place="7" resultid="2685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7742" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4725" />
                    <RANKING order="2" place="2" resultid="4069" />
                    <RANKING order="3" place="3" resultid="2561" />
                    <RANKING order="4" place="-1" resultid="3651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7743" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5530" />
                    <RANKING order="2" place="2" resultid="5283" />
                    <RANKING order="3" place="3" resultid="3186" />
                    <RANKING order="4" place="4" resultid="4836" />
                    <RANKING order="5" place="5" resultid="2117" />
                    <RANKING order="6" place="6" resultid="2839" />
                    <RANKING order="7" place="-1" resultid="4604" />
                    <RANKING order="8" place="-1" resultid="3144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7744" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5651" />
                    <RANKING order="2" place="2" resultid="5594" />
                    <RANKING order="3" place="3" resultid="6031" />
                    <RANKING order="4" place="4" resultid="6099" />
                    <RANKING order="5" place="5" resultid="2568" />
                    <RANKING order="6" place="-1" resultid="2219" />
                    <RANKING order="7" place="-1" resultid="3412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7745" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3011" />
                    <RANKING order="2" place="2" resultid="2291" />
                    <RANKING order="3" place="3" resultid="4807" />
                    <RANKING order="4" place="4" resultid="3221" />
                    <RANKING order="5" place="5" resultid="2869" />
                    <RANKING order="6" place="6" resultid="2464" />
                    <RANKING order="7" place="7" resultid="4571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7746" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4261" />
                    <RANKING order="2" place="2" resultid="3660" />
                    <RANKING order="3" place="3" resultid="4364" />
                    <RANKING order="4" place="4" resultid="2812" />
                    <RANKING order="5" place="5" resultid="3611" />
                    <RANKING order="6" place="6" resultid="4002" />
                    <RANKING order="7" place="7" resultid="3994" />
                    <RANKING order="8" place="8" resultid="5829" />
                    <RANKING order="9" place="-1" resultid="2249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7747" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2045" />
                    <RANKING order="2" place="2" resultid="3201" />
                    <RANKING order="3" place="3" resultid="3234" />
                    <RANKING order="4" place="4" resultid="2879" />
                    <RANKING order="5" place="5" resultid="5096" />
                    <RANKING order="6" place="6" resultid="5921" />
                    <RANKING order="7" place="7" resultid="6187" />
                    <RANKING order="8" place="8" resultid="4552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7748" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6016" />
                    <RANKING order="2" place="2" resultid="6092" />
                    <RANKING order="3" place="3" resultid="5045" />
                    <RANKING order="4" place="4" resultid="6219" />
                    <RANKING order="5" place="5" resultid="3416" />
                    <RANKING order="6" place="6" resultid="5586" />
                    <RANKING order="7" place="7" resultid="4967" />
                    <RANKING order="8" place="8" resultid="5033" />
                    <RANKING order="9" place="-1" resultid="2447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7749" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4284" />
                    <RANKING order="2" place="2" resultid="5484" />
                    <RANKING order="3" place="3" resultid="2159" />
                    <RANKING order="4" place="4" resultid="2017" />
                    <RANKING order="5" place="-1" resultid="4437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7750" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5147" />
                    <RANKING order="2" place="2" resultid="5848" />
                    <RANKING order="3" place="3" resultid="5898" />
                    <RANKING order="4" place="-1" resultid="3455" />
                    <RANKING order="5" place="-1" resultid="3566" />
                    <RANKING order="6" place="-1" resultid="4631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7751" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3844" />
                    <RANKING order="2" place="2" resultid="5742" />
                    <RANKING order="3" place="3" resultid="2155" />
                    <RANKING order="4" place="4" resultid="3976" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7332" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7333" daytime="10:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7334" daytime="10:17" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7335" daytime="10:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7336" daytime="10:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7337" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7338" daytime="10:34" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7339" daytime="10:38" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1320" daytime="12:04" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7797" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7798" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7799" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4102" />
                    <RANKING order="2" place="2" resultid="4565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7800" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5687" />
                    <RANKING order="2" place="2" resultid="2638" />
                    <RANKING order="3" place="3" resultid="2695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7801" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2202" />
                    <RANKING order="2" place="2" resultid="3796" />
                    <RANKING order="3" place="3" resultid="3127" />
                    <RANKING order="4" place="4" resultid="2686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7802" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5104" />
                    <RANKING order="2" place="2" resultid="4726" />
                    <RANKING order="3" place="-1" resultid="2091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7803" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5284" />
                    <RANKING order="2" place="2" resultid="5531" />
                    <RANKING order="3" place="3" resultid="3187" />
                    <RANKING order="4" place="4" resultid="2475" />
                    <RANKING order="5" place="5" resultid="5696" />
                    <RANKING order="6" place="6" resultid="4605" />
                    <RANKING order="7" place="7" resultid="2605" />
                    <RANKING order="8" place="8" resultid="2751" />
                    <RANKING order="9" place="9" resultid="4655" />
                    <RANKING order="10" place="10" resultid="2759" />
                    <RANKING order="11" place="-1" resultid="6502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7804" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2413" />
                    <RANKING order="2" place="2" resultid="3855" />
                    <RANKING order="3" place="3" resultid="4618" />
                    <RANKING order="4" place="4" resultid="2432" />
                    <RANKING order="5" place="5" resultid="4799" />
                    <RANKING order="6" place="6" resultid="5748" />
                    <RANKING order="7" place="7" resultid="2569" />
                    <RANKING order="8" place="8" resultid="6100" />
                    <RANKING order="9" place="9" resultid="3120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7805" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5620" />
                    <RANKING order="2" place="2" resultid="6306" />
                    <RANKING order="3" place="3" resultid="4581" />
                    <RANKING order="4" place="4" resultid="6479" />
                    <RANKING order="5" place="5" resultid="4923" />
                    <RANKING order="6" place="6" resultid="3082" />
                    <RANKING order="7" place="7" resultid="2388" />
                    <RANKING order="8" place="8" resultid="5820" />
                    <RANKING order="9" place="9" resultid="4276" />
                    <RANKING order="10" place="10" resultid="4808" />
                    <RANKING order="11" place="11" resultid="2721" />
                    <RANKING order="12" place="12" resultid="5141" />
                    <RANKING order="13" place="13" resultid="4290" />
                    <RANKING order="14" place="14" resultid="4572" />
                    <RANKING order="15" place="15" resultid="2233" />
                    <RANKING order="16" place="16" resultid="3965" />
                    <RANKING order="17" place="-1" resultid="2278" />
                    <RANKING order="18" place="-1" resultid="3181" />
                    <RANKING order="19" place="-1" resultid="6471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7806" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4262" />
                    <RANKING order="2" place="2" resultid="2362" />
                    <RANKING order="3" place="3" resultid="2669" />
                    <RANKING order="4" place="4" resultid="3743" />
                    <RANKING order="5" place="5" resultid="4365" />
                    <RANKING order="6" place="6" resultid="3685" />
                    <RANKING order="7" place="7" resultid="5883" />
                    <RANKING order="8" place="8" resultid="3399" />
                    <RANKING order="9" place="9" resultid="5077" />
                    <RANKING order="10" place="10" resultid="6346" />
                    <RANKING order="11" place="11" resultid="2813" />
                    <RANKING order="12" place="12" resultid="4529" />
                    <RANKING order="13" place="13" resultid="4003" />
                    <RANKING order="14" place="-1" resultid="4307" />
                    <RANKING order="15" place="-1" resultid="4427" />
                    <RANKING order="16" place="-1" resultid="5771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7807" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3202" />
                    <RANKING order="2" place="2" resultid="6373" />
                    <RANKING order="3" place="3" resultid="2901" />
                    <RANKING order="4" place="4" resultid="4961" />
                    <RANKING order="5" place="5" resultid="3054" />
                    <RANKING order="6" place="6" resultid="5716" />
                    <RANKING order="7" place="7" resultid="3021" />
                    <RANKING order="8" place="8" resultid="2880" />
                    <RANKING order="9" place="9" resultid="2014" />
                    <RANKING order="10" place="10" resultid="5015" />
                    <RANKING order="11" place="11" resultid="5628" />
                    <RANKING order="12" place="12" resultid="2056" />
                    <RANKING order="13" place="13" resultid="4316" />
                    <RANKING order="14" place="14" resultid="6386" />
                    <RANKING order="15" place="15" resultid="3254" />
                    <RANKING order="16" place="16" resultid="5026" />
                    <RANKING order="17" place="17" resultid="4553" />
                    <RANKING order="18" place="18" resultid="5040" />
                    <RANKING order="19" place="19" resultid="3528" />
                    <RANKING order="20" place="20" resultid="5256" />
                    <RANKING order="21" place="21" resultid="4832" />
                    <RANKING order="22" place="22" resultid="2256" />
                    <RANKING order="23" place="-1" resultid="6381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7808" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4733" />
                    <RANKING order="2" place="2" resultid="6427" />
                    <RANKING order="3" place="3" resultid="3720" />
                    <RANKING order="4" place="4" resultid="5046" />
                    <RANKING order="5" place="5" resultid="6093" />
                    <RANKING order="6" place="6" resultid="4935" />
                    <RANKING order="7" place="7" resultid="5206" />
                    <RANKING order="8" place="8" resultid="3417" />
                    <RANKING order="9" place="9" resultid="5587" />
                    <RANKING order="10" place="10" resultid="5216" />
                    <RANKING order="11" place="11" resultid="4968" />
                    <RANKING order="12" place="12" resultid="4942" />
                    <RANKING order="13" place="13" resultid="5034" />
                    <RANKING order="14" place="14" resultid="4505" />
                    <RANKING order="15" place="-1" resultid="6865" />
                    <RANKING order="16" place="-1" resultid="3887" />
                    <RANKING order="17" place="-1" resultid="4452" />
                    <RANKING order="18" place="-1" resultid="4589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7809" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4285" />
                    <RANKING order="2" place="2" resultid="3227" />
                    <RANKING order="3" place="3" resultid="2856" />
                    <RANKING order="4" place="4" resultid="4398" />
                    <RANKING order="5" place="5" resultid="4243" />
                    <RANKING order="6" place="6" resultid="5250" />
                    <RANKING order="7" place="7" resultid="2953" />
                    <RANKING order="8" place="8" resultid="5915" />
                    <RANKING order="9" place="9" resultid="2847" />
                    <RANKING order="10" place="10" resultid="2018" />
                    <RANKING order="11" place="-1" resultid="2213" />
                    <RANKING order="12" place="-1" resultid="3436" />
                    <RANKING order="13" place="-1" resultid="3498" />
                    <RANKING order="14" place="-1" resultid="4892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7810" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6174" />
                    <RANKING order="2" place="2" resultid="3729" />
                    <RANKING order="3" place="3" resultid="5226" />
                    <RANKING order="4" place="4" resultid="2283" />
                    <RANKING order="5" place="5" resultid="5849" />
                    <RANKING order="6" place="6" resultid="2407" />
                    <RANKING order="7" place="7" resultid="6441" />
                    <RANKING order="8" place="-1" resultid="2189" />
                    <RANKING order="9" place="-1" resultid="2337" />
                    <RANKING order="10" place="-1" resultid="2519" />
                    <RANKING order="11" place="-1" resultid="3456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7811" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4202" />
                    <RANKING order="2" place="2" resultid="4187" />
                    <RANKING order="3" place="3" resultid="3846" />
                    <RANKING order="4" place="4" resultid="2629" />
                    <RANKING order="5" place="5" resultid="2612" />
                    <RANKING order="6" place="6" resultid="3977" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7377" daytime="12:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7378" daytime="12:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7379" daytime="12:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7380" daytime="12:13" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7381" daytime="12:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7382" daytime="12:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7383" daytime="12:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7384" daytime="12:22" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7385" daytime="12:24" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7386" daytime="12:26" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7387" daytime="12:28" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7388" daytime="12:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7389" daytime="12:32" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7390" daytime="12:33" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1352" daytime="12:52" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7827" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7828" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7829" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7830" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7831" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4782" />
                    <RANKING order="2" place="2" resultid="2422" />
                    <RANKING order="3" place="3" resultid="2730" />
                    <RANKING order="4" place="4" resultid="3934" />
                    <RANKING order="5" place="-1" resultid="5167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7832" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2712" />
                    <RANKING order="2" place="2" resultid="5779" />
                    <RANKING order="3" place="3" resultid="2764" />
                    <RANKING order="4" place="4" resultid="4109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7833" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5553" />
                    <RANKING order="2" place="2" resultid="2118" />
                    <RANKING order="3" place="3" resultid="4837" />
                    <RANKING order="4" place="4" resultid="5864" />
                    <RANKING order="5" place="5" resultid="3242" />
                    <RANKING order="6" place="6" resultid="3150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7834" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5595" />
                    <RANKING order="2" place="2" resultid="6036" />
                    <RANKING order="3" place="3" resultid="3280" />
                    <RANKING order="4" place="-1" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7835" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2389" />
                    <RANKING order="2" place="2" resultid="2805" />
                    <RANKING order="3" place="3" resultid="5523" />
                    <RANKING order="4" place="4" resultid="6249" />
                    <RANKING order="5" place="5" resultid="2870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7836" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6148" />
                    <RANKING order="2" place="2" resultid="4249" />
                    <RANKING order="3" place="3" resultid="3676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7837" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2046" />
                    <RANKING order="2" place="2" resultid="6382" />
                    <RANKING order="3" place="3" resultid="6008" />
                    <RANKING order="4" place="4" resultid="2881" />
                    <RANKING order="5" place="5" resultid="4930" />
                    <RANKING order="6" place="6" resultid="3235" />
                    <RANKING order="7" place="7" resultid="5629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7838" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6220" />
                    <RANKING order="2" place="2" resultid="6025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7839" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="5485" />
                    <RANKING order="3" place="3" resultid="2160" />
                    <RANKING order="4" place="4" resultid="2585" />
                    <RANKING order="5" place="5" resultid="4438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7840" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5792" />
                    <RANKING order="2" place="2" resultid="6175" />
                    <RANKING order="3" place="3" resultid="3510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7841" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6361" />
                    <RANKING order="2" place="-1" resultid="2136" />
                    <RANKING order="3" place="-1" resultid="3824" />
                    <RANKING order="4" place="-1" resultid="4209" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7394" daytime="12:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7395" daytime="12:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7396" daytime="13:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7397" daytime="13:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7398" daytime="13:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-11-16" daytime="16:00" endtime="21:29" name="Zimowe Mistrzostwa Polskiw Pływaniu Masters BLOK III" number="3" warmupfrom="15:00" warmupuntil="15:50">
          <EVENTS>
            <EVENT eventid="1417" daytime="16:20" gender="M" number="23" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7885" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7886" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2245" />
                    <RANKING order="2" place="-1" resultid="2893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7887" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4103" />
                    <RANKING order="2" place="2" resultid="4566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7888" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4637" />
                    <RANKING order="2" place="2" resultid="2639" />
                    <RANKING order="3" place="3" resultid="2508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7889" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                    <RANKING order="2" place="2" resultid="5168" />
                    <RANKING order="3" place="3" resultid="3949" />
                    <RANKING order="4" place="4" resultid="2687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7890" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4727" />
                    <RANKING order="2" place="2" resultid="4070" />
                    <RANKING order="3" place="3" resultid="2562" />
                    <RANKING order="4" place="4" resultid="5935" />
                    <RANKING order="5" place="5" resultid="3249" />
                    <RANKING order="6" place="-1" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7891" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5532" />
                    <RANKING order="2" place="2" resultid="3188" />
                    <RANKING order="3" place="3" resultid="2476" />
                    <RANKING order="4" place="4" resultid="2119" />
                    <RANKING order="5" place="5" resultid="4606" />
                    <RANKING order="6" place="6" resultid="4838" />
                    <RANKING order="7" place="7" resultid="5814" />
                    <RANKING order="8" place="8" resultid="4846" />
                    <RANKING order="9" place="-1" resultid="3145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7892" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3413" />
                    <RANKING order="2" place="2" resultid="5652" />
                    <RANKING order="3" place="3" resultid="6032" />
                    <RANKING order="4" place="4" resultid="5596" />
                    <RANKING order="5" place="5" resultid="2570" />
                    <RANKING order="6" place="6" resultid="6101" />
                    <RANKING order="7" place="7" resultid="3290" />
                    <RANKING order="8" place="-1" resultid="4359" />
                    <RANKING order="9" place="-1" resultid="4619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7893" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3012" />
                    <RANKING order="2" place="2" resultid="2293" />
                    <RANKING order="3" place="3" resultid="5821" />
                    <RANKING order="4" place="4" resultid="3222" />
                    <RANKING order="5" place="5" resultid="5878" />
                    <RANKING order="6" place="6" resultid="6124" />
                    <RANKING order="7" place="7" resultid="4809" />
                    <RANKING order="8" place="8" resultid="4291" />
                    <RANKING order="9" place="9" resultid="4573" />
                    <RANKING order="10" place="10" resultid="5142" />
                    <RANKING order="11" place="11" resultid="3966" />
                    <RANKING order="12" place="12" resultid="2234" />
                    <RANKING order="13" place="-1" resultid="2167" />
                    <RANKING order="14" place="-1" resultid="6307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7894" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4263" />
                    <RANKING order="2" place="2" resultid="3661" />
                    <RANKING order="3" place="3" resultid="3686" />
                    <RANKING order="4" place="4" resultid="4366" />
                    <RANKING order="5" place="5" resultid="2811" />
                    <RANKING order="6" place="6" resultid="3612" />
                    <RANKING order="7" place="7" resultid="3133" />
                    <RANKING order="8" place="8" resultid="4004" />
                    <RANKING order="9" place="9" resultid="4308" />
                    <RANKING order="10" place="10" resultid="3996" />
                    <RANKING order="11" place="11" resultid="5830" />
                    <RANKING order="12" place="-1" resultid="2250" />
                    <RANKING order="13" place="-1" resultid="4428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7895" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3203" />
                    <RANKING order="2" place="2" resultid="4696" />
                    <RANKING order="3" place="3" resultid="3055" />
                    <RANKING order="4" place="4" resultid="2902" />
                    <RANKING order="5" place="5" resultid="5098" />
                    <RANKING order="6" place="6" resultid="6189" />
                    <RANKING order="7" place="7" resultid="5922" />
                    <RANKING order="8" place="8" resultid="6387" />
                    <RANKING order="9" place="9" resultid="4554" />
                    <RANKING order="10" place="10" resultid="3050" />
                    <RANKING order="11" place="11" resultid="2492" />
                    <RANKING order="12" place="12" resultid="2740" />
                    <RANKING order="13" place="-1" resultid="1997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7896" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6018" />
                    <RANKING order="2" place="2" resultid="5047" />
                    <RANKING order="3" place="3" resultid="6094" />
                    <RANKING order="4" place="4" resultid="4936" />
                    <RANKING order="5" place="5" resultid="5055" />
                    <RANKING order="6" place="6" resultid="4888" />
                    <RANKING order="7" place="7" resultid="3418" />
                    <RANKING order="8" place="8" resultid="6221" />
                    <RANKING order="9" place="9" resultid="5588" />
                    <RANKING order="10" place="10" resultid="4969" />
                    <RANKING order="11" place="11" resultid="4453" />
                    <RANKING order="12" place="12" resultid="5052" />
                    <RANKING order="13" place="13" resultid="5035" />
                    <RANKING order="14" place="14" resultid="2449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7897" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4286" />
                    <RANKING order="2" place="2" resultid="3228" />
                    <RANKING order="3" place="3" resultid="5998" />
                    <RANKING order="4" place="4" resultid="2161" />
                    <RANKING order="5" place="5" resultid="3864" />
                    <RANKING order="6" place="6" resultid="5916" />
                    <RANKING order="7" place="7" resultid="3427" />
                    <RANKING order="8" place="8" resultid="2019" />
                    <RANKING order="9" place="-1" resultid="3437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7898" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2960" />
                    <RANKING order="2" place="2" resultid="5899" />
                    <RANKING order="3" place="-1" resultid="2338" />
                    <RANKING order="4" place="-1" resultid="3457" />
                    <RANKING order="5" place="-1" resultid="3567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7899" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4203" />
                    <RANKING order="2" place="2" resultid="4188" />
                    <RANKING order="3" place="3" resultid="3847" />
                    <RANKING order="4" place="4" resultid="2630" />
                    <RANKING order="5" place="5" resultid="5743" />
                    <RANKING order="6" place="6" resultid="2156" />
                    <RANKING order="7" place="7" resultid="2661" />
                    <RANKING order="8" place="8" resultid="3978" />
                    <RANKING order="9" place="9" resultid="3564" />
                    <RANKING order="10" place="-1" resultid="2320" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7414" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7415" daytime="16:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7416" daytime="16:27" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7417" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7418" daytime="16:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7419" daytime="16:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7420" daytime="16:37" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7421" daytime="16:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7422" daytime="16:42" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7423" daytime="16:44" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7424" daytime="16:46" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7425" daytime="16:48" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1497" daytime="18:15" gender="F" number="28" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7960" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7961" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7962" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7963" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7964" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7965" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5667" />
                    <RANKING order="2" place="2" resultid="5964" />
                    <RANKING order="3" place="3" resultid="2351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7966" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3088" />
                    <RANKING order="2" place="2" resultid="2472" />
                    <RANKING order="3" place="3" resultid="3811" />
                    <RANKING order="4" place="4" resultid="3912" />
                    <RANKING order="5" place="5" resultid="2267" />
                    <RANKING order="6" place="6" resultid="5294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7967" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5800" />
                    <RANKING order="2" place="2" resultid="4774" />
                    <RANKING order="3" place="3" resultid="4061" />
                    <RANKING order="4" place="4" resultid="4232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7968" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2556" />
                    <RANKING order="2" place="2" resultid="6243" />
                    <RANKING order="3" place="3" resultid="4271" />
                    <RANKING order="4" place="4" resultid="5956" />
                    <RANKING order="5" place="5" resultid="6205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7969" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3803" />
                    <RANKING order="2" place="2" resultid="5505" />
                    <RANKING order="3" place="3" resultid="5091" />
                    <RANKING order="4" place="4" resultid="3920" />
                    <RANKING order="5" place="5" resultid="6214" />
                    <RANKING order="6" place="6" resultid="5892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7970" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2483" />
                    <RANKING order="2" place="2" resultid="3695" />
                    <RANKING order="3" place="3" resultid="5739" />
                    <RANKING order="4" place="-1" resultid="4499" />
                    <RANKING order="5" place="-1" resultid="5513" />
                    <RANKING order="6" place="-1" resultid="6168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7971" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4488" />
                    <RANKING order="2" place="2" resultid="3712" />
                    <RANKING order="3" place="3" resultid="4645" />
                    <RANKING order="4" place="4" resultid="6392" />
                    <RANKING order="5" place="5" resultid="2866" />
                    <RANKING order="6" place="6" resultid="4028" />
                    <RANKING order="7" place="7" resultid="2398" />
                    <RANKING order="8" place="8" resultid="5613" />
                    <RANKING order="9" place="-1" resultid="5605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7972" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4042" />
                    <RANKING order="2" place="2" resultid="4745" />
                    <RANKING order="3" place="3" resultid="3705" />
                    <RANKING order="4" place="4" resultid="2829" />
                    <RANKING order="5" place="5" resultid="5136" />
                    <RANKING order="6" place="6" resultid="3471" />
                    <RANKING order="7" place="7" resultid="5580" />
                    <RANKING order="8" place="8" resultid="2648" />
                    <RANKING order="9" place="9" resultid="4663" />
                    <RANKING order="10" place="10" resultid="5873" />
                    <RANKING order="11" place="11" resultid="6463" />
                    <RANKING order="12" place="-1" resultid="4342" />
                    <RANKING order="13" place="-1" resultid="4541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7973" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2982" />
                    <RANKING order="2" place="2" resultid="2038" />
                    <RANKING order="3" place="3" resultid="6132" />
                    <RANKING order="4" place="4" resultid="2143" />
                    <RANKING order="5" place="5" resultid="5845" />
                    <RANKING order="6" place="6" resultid="3485" />
                    <RANKING order="7" place="7" resultid="3297" />
                    <RANKING order="8" place="8" resultid="4448" />
                    <RANKING order="9" place="-1" resultid="3333" />
                    <RANKING order="10" place="-1" resultid="4443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7974" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4196" />
                    <RANKING order="2" place="2" resultid="3737" />
                    <RANKING order="3" place="3" resultid="3840" />
                    <RANKING order="4" place="4" resultid="3560" />
                    <RANKING order="5" place="-1" resultid="3554" />
                    <RANKING order="6" place="-1" resultid="4216" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7468" daytime="18:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7469" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7470" daytime="18:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7471" daytime="18:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7472" daytime="18:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7473" daytime="18:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7474" daytime="18:39" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1481" daytime="17:50" gender="M" number="27" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7945" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7946" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7947" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4104" />
                    <RANKING order="2" place="2" resultid="4567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7948" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5689" />
                    <RANKING order="2" place="2" resultid="3943" />
                    <RANKING order="3" place="3" resultid="2509" />
                    <RANKING order="4" place="4" resultid="2704" />
                    <RANKING order="5" place="-1" resultid="5176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7949" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3099" />
                    <RANKING order="2" place="2" resultid="3784" />
                    <RANKING order="3" place="3" resultid="2456" />
                    <RANKING order="4" place="4" resultid="2423" />
                    <RANKING order="5" place="-1" resultid="3950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7950" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4600" />
                    <RANKING order="2" place="2" resultid="2127" />
                    <RANKING order="3" place="3" resultid="2713" />
                    <RANKING order="4" place="4" resultid="5780" />
                    <RANKING order="5" place="5" resultid="2302" />
                    <RANKING order="6" place="6" resultid="3250" />
                    <RANKING order="7" place="-1" resultid="3209" />
                    <RANKING order="8" place="-1" resultid="3653" />
                    <RANKING order="9" place="-1" resultid="5679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7951" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3215" />
                    <RANKING order="2" place="2" resultid="3768" />
                    <RANKING order="3" place="3" resultid="5697" />
                    <RANKING order="4" place="4" resultid="4159" />
                    <RANKING order="5" place="5" resultid="2752" />
                    <RANKING order="6" place="-1" resultid="4357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7952" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3857" />
                    <RANKING order="2" place="2" resultid="2414" />
                    <RANKING order="3" place="3" resultid="2434" />
                    <RANKING order="4" place="4" resultid="4801" />
                    <RANKING order="5" place="5" resultid="2345" />
                    <RANKING order="6" place="-1" resultid="2571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7953" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4924" />
                    <RANKING order="2" place="2" resultid="4583" />
                    <RANKING order="3" place="3" resultid="5993" />
                    <RANKING order="4" place="4" resultid="2801" />
                    <RANKING order="5" place="5" resultid="5524" />
                    <RANKING order="6" place="6" resultid="2465" />
                    <RANKING order="7" place="7" resultid="4299" />
                    <RANKING order="8" place="8" resultid="5085" />
                    <RANKING order="9" place="9" resultid="3967" />
                    <RANKING order="10" place="-1" resultid="2279" />
                    <RANKING order="11" place="-1" resultid="4277" />
                    <RANKING order="12" place="-1" resultid="5622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7954" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3745" />
                    <RANKING order="2" place="2" resultid="2670" />
                    <RANKING order="3" place="3" resultid="4388" />
                    <RANKING order="4" place="4" resultid="5078" />
                    <RANKING order="5" place="5" resultid="3400" />
                    <RANKING order="6" place="6" resultid="5885" />
                    <RANKING order="7" place="7" resultid="6196" />
                    <RANKING order="8" place="8" resultid="3617" />
                    <RANKING order="9" place="9" resultid="3677" />
                    <RANKING order="10" place="10" resultid="5831" />
                    <RANKING order="11" place="-1" resultid="5198" />
                    <RANKING order="12" place="-1" resultid="5772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7955" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2996" />
                    <RANKING order="2" place="2" resultid="6047" />
                    <RANKING order="3" place="3" resultid="3044" />
                    <RANKING order="4" place="4" resultid="2058" />
                    <RANKING order="5" place="5" resultid="4833" />
                    <RANKING order="6" place="6" resultid="2258" />
                    <RANKING order="7" place="-1" resultid="2741" />
                    <RANKING order="8" place="-1" resultid="3056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7956" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3722" />
                    <RANKING order="2" place="2" resultid="4735" />
                    <RANKING order="3" place="3" resultid="3195" />
                    <RANKING order="4" place="4" resultid="3888" />
                    <RANKING order="5" place="5" resultid="4179" />
                    <RANKING order="6" place="6" resultid="2544" />
                    <RANKING order="7" place="7" resultid="5222" />
                    <RANKING order="8" place="-1" resultid="4590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7957" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2969" />
                    <RANKING order="2" place="2" resultid="5858" />
                    <RANKING order="3" place="3" resultid="4244" />
                    <RANKING order="4" place="4" resultid="3499" />
                    <RANKING order="5" place="5" resultid="4714" />
                    <RANKING order="6" place="6" resultid="4670" />
                    <RANKING order="7" place="7" resultid="3865" />
                    <RANKING order="8" place="-1" resultid="4439" />
                    <RANKING order="9" place="-1" resultid="5486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7958" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5233" />
                    <RANKING order="2" place="2" resultid="2284" />
                    <RANKING order="3" place="3" resultid="5900" />
                    <RANKING order="4" place="-1" resultid="2339" />
                    <RANKING order="5" place="-1" resultid="3458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7959" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4210" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7459" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7460" daytime="17:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7461" daytime="17:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7462" daytime="18:01" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7463" daytime="18:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7464" daytime="18:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7465" daytime="18:09" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7466" daytime="18:11" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7467" daytime="18:13" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1577" daytime="20:29" gender="M" number="33" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8005" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8006" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="8007" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8008" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2640" />
                    <RANKING order="2" place="2" resultid="2697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8009" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2204" />
                    <RANKING order="2" place="2" resultid="5169" />
                    <RANKING order="3" place="3" resultid="2424" />
                    <RANKING order="4" place="4" resultid="2732" />
                    <RANKING order="5" place="5" resultid="3936" />
                    <RANKING order="6" place="-1" resultid="4784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8010" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4728" />
                    <RANKING order="2" place="2" resultid="2714" />
                    <RANKING order="3" place="3" resultid="5781" />
                    <RANKING order="4" place="-1" resultid="2765" />
                    <RANKING order="5" place="-1" resultid="4110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8011" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5286" />
                    <RANKING order="2" place="2" resultid="5698" />
                    <RANKING order="3" place="3" resultid="2120" />
                    <RANKING order="4" place="4" resultid="3189" />
                    <RANKING order="5" place="5" resultid="2606" />
                    <RANKING order="6" place="6" resultid="3244" />
                    <RANKING order="7" place="-1" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8012" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5749" />
                    <RANKING order="2" place="2" resultid="5597" />
                    <RANKING order="3" place="3" resultid="6102" />
                    <RANKING order="4" place="4" resultid="6038" />
                    <RANKING order="5" place="5" resultid="2886" />
                    <RANKING order="6" place="-1" resultid="2221" />
                    <RANKING order="7" place="-1" resultid="3281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8013" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2804" />
                    <RANKING order="2" place="2" resultid="2391" />
                    <RANKING order="3" place="3" resultid="6250" />
                    <RANKING order="4" place="4" resultid="2723" />
                    <RANKING order="5" place="5" resultid="2466" />
                    <RANKING order="6" place="6" resultid="2235" />
                    <RANKING order="7" place="-1" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8014" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6150" />
                    <RANKING order="2" place="2" resultid="3662" />
                    <RANKING order="3" place="3" resultid="2671" />
                    <RANKING order="4" place="4" resultid="4368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8015" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2048" />
                    <RANKING order="2" place="2" resultid="3236" />
                    <RANKING order="3" place="3" resultid="6141" />
                    <RANKING order="4" place="4" resultid="2882" />
                    <RANKING order="5" place="5" resultid="5923" />
                    <RANKING order="6" place="6" resultid="5631" />
                    <RANKING order="7" place="7" resultid="3529" />
                    <RANKING order="8" place="-1" resultid="2112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8016" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3889" />
                    <RANKING order="2" place="2" resultid="5589" />
                    <RANKING order="3" place="3" resultid="4971" />
                    <RANKING order="4" place="-1" resultid="6222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8017" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4400" />
                    <RANKING order="2" place="2" resultid="2586" />
                    <RANKING order="3" place="-1" resultid="3500" />
                    <RANKING order="4" place="-1" resultid="4440" />
                    <RANKING order="5" place="-1" resultid="5487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8018" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5794" />
                    <RANKING order="2" place="2" resultid="6177" />
                    <RANKING order="3" place="3" resultid="3511" />
                    <RANKING order="4" place="4" resultid="2285" />
                    <RANKING order="5" place="-1" resultid="3459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8019" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4211" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8152" daytime="20:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8153" daytime="20:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8154" daytime="20:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8155" daytime="21:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8156" daytime="21:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8157" daytime="21:21" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8158" daytime="21:28" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1545" daytime="19:46" gender="M" number="31" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7863" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3305" />
                    <RANKING order="2" place="2" resultid="4135" />
                    <RANKING order="3" place="3" resultid="3953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7864" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3307" />
                    <RANKING order="2" place="2" resultid="4852" />
                    <RANKING order="3" place="3" resultid="5763" />
                    <RANKING order="4" place="4" resultid="2327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7865" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4759" />
                    <RANKING order="2" place="2" resultid="6873" />
                    <RANKING order="3" place="3" resultid="6271" />
                    <RANKING order="4" place="4" resultid="3320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7866" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6408" />
                    <RANKING order="2" place="2" resultid="6059" />
                    <RANKING order="3" place="3" resultid="4280" />
                    <RANKING order="4" place="4" resultid="5065" />
                    <RANKING order="5" place="5" resultid="3309" />
                    <RANKING order="6" place="6" resultid="6270" />
                    <RANKING order="7" place="7" resultid="5064" />
                    <RANKING order="8" place="8" resultid="3440" />
                    <RANKING order="9" place="9" resultid="3638" />
                    <RANKING order="10" place="10" resultid="3070" />
                    <RANKING order="11" place="11" resultid="4549" />
                    <RANKING order="12" place="12" resultid="4458" />
                    <RANKING order="13" place="13" resultid="5271" />
                    <RANKING order="14" place="-1" resultid="5658" />
                    <RANKING order="15" place="-1" resultid="3039" />
                    <RANKING order="16" place="-1" resultid="4354" />
                    <RANKING order="17" place="-1" resultid="5158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7867" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3031" />
                    <RANKING order="2" place="2" resultid="4760" />
                    <RANKING order="3" place="3" resultid="6269" />
                    <RANKING order="4" place="4" resultid="5270" />
                    <RANKING order="5" place="5" resultid="4763" />
                    <RANKING order="6" place="6" resultid="4906" />
                    <RANKING order="7" place="7" resultid="3032" />
                    <RANKING order="8" place="8" resultid="6062" />
                    <RANKING order="9" place="9" resultid="4353" />
                    <RANKING order="10" place="10" resultid="5063" />
                    <RANKING order="11" place="11" resultid="2874" />
                    <RANKING order="12" place="-1" resultid="6405" />
                    <RANKING order="13" place="-1" resultid="3605" />
                    <RANKING order="14" place="-1" resultid="5066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7868" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2215" />
                    <RANKING order="2" place="2" resultid="3604" />
                    <RANKING order="3" place="-1" resultid="3603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7869" agemax="99" agemin="80" name="0" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7492" daytime="19:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7493" daytime="19:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7494" daytime="19:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7495" daytime="19:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7496" daytime="20:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1433" daytime="16:50" gender="F" number="24" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7900" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7901" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7902" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7903" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7904" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7905" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3790" />
                    <RANKING order="2" place="2" resultid="5666" />
                    <RANKING order="3" place="3" resultid="4086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7906" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3087" />
                    <RANKING order="2" place="2" resultid="6487" />
                    <RANKING order="3" place="3" resultid="4825" />
                    <RANKING order="4" place="4" resultid="4117" />
                    <RANKING order="5" place="-1" resultid="2311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7907" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3106" />
                    <RANKING order="2" place="2" resultid="5674" />
                    <RANKING order="3" place="3" resultid="2795" />
                    <RANKING order="4" place="4" resultid="6332" />
                    <RANKING order="5" place="5" resultid="4793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7908" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2940" />
                    <RANKING order="2" place="2" resultid="3990" />
                    <RANKING order="3" place="3" resultid="2373" />
                    <RANKING order="4" place="4" resultid="3408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7909" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3163" />
                    <RANKING order="2" place="2" resultid="5493" />
                    <RANKING order="3" place="3" resultid="4766" />
                    <RANKING order="4" place="4" resultid="6213" />
                    <RANKING order="5" place="5" resultid="6397" />
                    <RANKING order="6" place="6" resultid="4375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7910" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2599" />
                    <RANKING order="2" place="2" resultid="4988" />
                    <RANKING order="3" place="3" resultid="4498" />
                    <RANKING order="4" place="4" resultid="3169" />
                    <RANKING order="5" place="5" resultid="5512" />
                    <RANKING order="6" place="6" resultid="5560" />
                    <RANKING order="7" place="7" resultid="3694" />
                    <RANKING order="8" place="8" resultid="2935" />
                    <RANKING order="9" place="9" resultid="5738" />
                    <RANKING order="10" place="10" resultid="4979" />
                    <RANKING order="11" place="11" resultid="5264" />
                    <RANKING order="12" place="12" resultid="5643" />
                    <RANKING order="13" place="13" resultid="3960" />
                    <RANKING order="14" place="-1" resultid="6413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7911" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3382" />
                    <RANKING order="2" place="2" resultid="2442" />
                    <RANKING order="3" place="3" resultid="2817" />
                    <RANKING order="4" place="4" resultid="4644" />
                    <RANKING order="5" place="5" resultid="5604" />
                    <RANKING order="6" place="6" resultid="6228" />
                    <RANKING order="7" place="7" resultid="2865" />
                    <RANKING order="8" place="8" resultid="3388" />
                    <RANKING order="9" place="-1" resultid="4954" />
                    <RANKING order="10" place="-1" resultid="4008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7912" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5810" />
                    <RANKING order="2" place="2" resultid="5245" />
                    <RANKING order="3" place="3" resultid="3750" />
                    <RANKING order="4" place="4" resultid="2647" />
                    <RANKING order="5" place="5" resultid="6158" />
                    <RANKING order="6" place="6" resultid="4611" />
                    <RANKING order="7" place="7" resultid="3393" />
                    <RANKING order="8" place="8" resultid="4662" />
                    <RANKING order="9" place="9" resultid="6462" />
                    <RANKING order="10" place="10" resultid="5872" />
                    <RANKING order="11" place="-1" resultid="2991" />
                    <RANKING order="12" place="-1" resultid="5211" />
                    <RANKING order="13" place="-1" resultid="3115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7913" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6338" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="2782" />
                    <RANKING order="4" place="4" resultid="2779" />
                    <RANKING order="5" place="5" resultid="6131" />
                    <RANKING order="6" place="6" resultid="4414" />
                    <RANKING order="7" place="7" resultid="2550" />
                    <RANKING order="8" place="8" resultid="4688" />
                    <RANKING order="9" place="9" resultid="3872" />
                    <RANKING order="10" place="10" resultid="5844" />
                    <RANKING order="11" place="11" resultid="4720" />
                    <RANKING order="12" place="12" resultid="5496" />
                    <RANKING order="13" place="-1" resultid="2916" />
                    <RANKING order="14" place="-1" resultid="3332" />
                    <RANKING order="15" place="-1" resultid="4466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7914" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2622" />
                    <RANKING order="2" place="2" resultid="2180" />
                    <RANKING order="3" place="3" resultid="5967" />
                    <RANKING order="4" place="4" resultid="3557" />
                    <RANKING order="5" place="5" resultid="5907" />
                    <RANKING order="6" place="6" resultid="3839" />
                    <RANKING order="7" place="-1" resultid="5301" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7426" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7427" daytime="16:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7428" daytime="16:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7429" daytime="16:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7430" daytime="16:57" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7431" daytime="16:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7432" daytime="17:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7433" daytime="17:01" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7434" daytime="17:02" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1561" daytime="20:03" gender="F" number="32" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7990" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7991" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7992" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7993" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7994" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7995" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7996" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3448" />
                    <RANKING order="2" place="2" resultid="4826" />
                    <RANKING order="3" place="3" resultid="4151" />
                    <RANKING order="4" place="4" resultid="5295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7997" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4775" />
                    <RANKING order="2" place="2" resultid="5130" />
                    <RANKING order="3" place="3" resultid="5977" />
                    <RANKING order="4" place="4" resultid="4078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7998" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7999" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3158" />
                    <RANKING order="2" place="2" resultid="5506" />
                    <RANKING order="3" place="3" resultid="5494" />
                    <RANKING order="4" place="4" resultid="4325" />
                    <RANKING order="5" place="5" resultid="6448" />
                    <RANKING order="6" place="6" resultid="4767" />
                    <RANKING order="7" place="7" resultid="5116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8000" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3170" />
                    <RANKING order="2" place="2" resultid="3669" />
                    <RANKING order="3" place="3" resultid="4980" />
                    <RANKING order="4" place="-1" resultid="4903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8001" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3713" />
                    <RANKING order="2" place="2" resultid="6357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8002" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3006" />
                    <RANKING order="2" place="2" resultid="6159" />
                    <RANKING order="3" place="3" resultid="4612" />
                    <RANKING order="4" place="-1" resultid="3882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8003" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8004" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5986" />
                    <RANKING order="2" place="2" resultid="4217" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8149" daytime="20:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8150" daytime="20:13" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8151" daytime="20:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1465" daytime="17:30" gender="F" number="26" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7930" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7931" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7932" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7933" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7934" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7935" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3791" />
                    <RANKING order="2" place="2" resultid="4132" />
                    <RANKING order="3" place="3" resultid="4167" />
                    <RANKING order="4" place="4" resultid="2075" />
                    <RANKING order="5" place="-1" resultid="4093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7936" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3447" />
                    <RANKING order="2" place="2" resultid="3810" />
                    <RANKING order="3" place="3" resultid="2312" />
                    <RANKING order="4" place="4" resultid="3911" />
                    <RANKING order="5" place="5" resultid="3984" />
                    <RANKING order="6" place="6" resultid="2593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7937" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3107" />
                    <RANKING order="2" place="2" resultid="4226" />
                    <RANKING order="3" place="3" resultid="5129" />
                    <RANKING order="4" place="4" resultid="4060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7938" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3991" />
                    <RANKING order="2" place="2" resultid="2944" />
                    <RANKING order="3" place="3" resultid="5955" />
                    <RANKING order="4" place="4" resultid="2273" />
                    <RANKING order="5" place="5" resultid="6204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7939" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                    <RANKING order="2" place="2" resultid="2355" />
                    <RANKING order="3" place="3" resultid="5806" />
                    <RANKING order="4" place="4" resultid="2084" />
                    <RANKING order="5" place="5" resultid="3919" />
                    <RANKING order="6" place="6" resultid="5891" />
                    <RANKING order="7" place="-1" resultid="3572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7940" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3176" />
                    <RANKING order="2" place="2" resultid="3075" />
                    <RANKING order="3" place="3" resultid="5561" />
                    <RANKING order="4" place="4" resultid="6167" />
                    <RANKING order="5" place="5" resultid="5111" />
                    <RANKING order="6" place="6" resultid="4303" />
                    <RANKING order="7" place="7" resultid="4435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7941" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3383" />
                    <RANKING order="2" place="2" resultid="4487" />
                    <RANKING order="3" place="3" resultid="4955" />
                    <RANKING order="4" place="4" resultid="5002" />
                    <RANKING order="5" place="5" resultid="2397" />
                    <RANKING order="6" place="6" resultid="4009" />
                    <RANKING order="7" place="7" resultid="4336" />
                    <RANKING order="8" place="-1" resultid="2488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7942" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3005" />
                    <RANKING order="2" place="2" resultid="8229" />
                    <RANKING order="3" place="3" resultid="6457" />
                    <RANKING order="4" place="4" resultid="5579" />
                    <RANKING order="5" place="5" resultid="2825" />
                    <RANKING order="6" place="-1" resultid="4341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7943" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3873" />
                    <RANKING order="2" place="2" resultid="4689" />
                    <RANKING order="3" place="3" resultid="5839" />
                    <RANKING order="4" place="4" resultid="2783" />
                    <RANKING order="5" place="5" resultid="4721" />
                    <RANKING order="6" place="6" resultid="5497" />
                    <RANKING order="7" place="7" resultid="3027" />
                    <RANKING order="8" place="8" resultid="5122" />
                    <RANKING order="9" place="9" resultid="2746" />
                    <RANKING order="10" place="-1" resultid="3296" />
                    <RANKING order="11" place="-1" resultid="4450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7944" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4195" />
                    <RANKING order="2" place="2" resultid="3272" />
                    <RANKING order="3" place="3" resultid="2332" />
                    <RANKING order="4" place="4" resultid="4019" />
                    <RANKING order="5" place="5" resultid="2623" />
                    <RANKING order="6" place="6" resultid="5968" />
                    <RANKING order="7" place="7" resultid="2678" />
                    <RANKING order="8" place="8" resultid="3540" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7452" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7453" daytime="17:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7454" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7455" daytime="17:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7456" daytime="17:43" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7457" daytime="17:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7458" daytime="17:48" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1400" daytime="16:00" gender="F" number="22" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7870" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7871" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7872" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7873" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="7874" agemax="74" agemin="70" name="J" />
                <AGEGROUP agegroupid="7875" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5963" />
                    <RANKING order="2" place="2" resultid="4085" />
                    <RANKING order="3" place="3" resultid="2350" />
                    <RANKING order="4" place="4" resultid="3774" />
                    <RANKING order="5" place="5" resultid="2074" />
                    <RANKING order="6" place="-1" resultid="4092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7876" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6486" />
                    <RANKING order="2" place="2" resultid="4116" />
                    <RANKING order="3" place="3" resultid="4150" />
                    <RANKING order="4" place="4" resultid="2266" />
                    <RANKING order="5" place="5" resultid="3983" />
                    <RANKING order="6" place="6" resultid="2592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7877" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5673" />
                    <RANKING order="2" place="2" resultid="2793" />
                    <RANKING order="3" place="3" resultid="4225" />
                    <RANKING order="4" place="4" resultid="6331" />
                    <RANKING order="5" place="5" resultid="5549" />
                    <RANKING order="6" place="6" resultid="4077" />
                    <RANKING order="7" place="7" resultid="4792" />
                    <RANKING order="8" place="-1" resultid="5976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7878" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3092" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="4270" />
                    <RANKING order="4" place="4" resultid="2272" />
                    <RANKING order="5" place="5" resultid="3973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7879" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3802" />
                    <RANKING order="2" place="2" resultid="4324" />
                    <RANKING order="3" place="3" resultid="4703" />
                    <RANKING order="4" place="4" resultid="2083" />
                    <RANKING order="5" place="5" resultid="3571" />
                    <RANKING order="6" place="-1" resultid="5090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7880" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2598" />
                    <RANKING order="2" place="2" resultid="3175" />
                    <RANKING order="3" place="3" resultid="3668" />
                    <RANKING order="4" place="4" resultid="4902" />
                    <RANKING order="5" place="5" resultid="3278" />
                    <RANKING order="6" place="6" resultid="3959" />
                    <RANKING order="7" place="7" resultid="3302" />
                    <RANKING order="8" place="8" resultid="5949" />
                    <RANKING order="9" place="-1" resultid="2934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7881" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2820" />
                    <RANKING order="2" place="2" resultid="4418" />
                    <RANKING order="3" place="3" resultid="4594" />
                    <RANKING order="4" place="4" resultid="4027" />
                    <RANKING order="5" place="5" resultid="5612" />
                    <RANKING order="6" place="-1" resultid="5648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7882" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3704" />
                    <RANKING order="2" place="2" resultid="4744" />
                    <RANKING order="3" place="3" resultid="4041" />
                    <RANKING order="4" place="4" resultid="3881" />
                    <RANKING order="5" place="5" resultid="5537" />
                    <RANKING order="6" place="-1" resultid="4540" />
                    <RANKING order="7" place="-1" resultid="3114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7883" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2549" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="3" resultid="5268" />
                    <RANKING order="4" place="4" resultid="4379" />
                    <RANKING order="5" place="5" resultid="4447" />
                    <RANKING order="6" place="-1" resultid="2915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7884" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5985" />
                    <RANKING order="2" place="2" resultid="3838" />
                    <RANKING order="3" place="3" resultid="2225" />
                    <RANKING order="4" place="4" resultid="5906" />
                    <RANKING order="5" place="5" resultid="5300" />
                    <RANKING order="6" place="6" resultid="2677" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7407" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7408" daytime="16:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7409" daytime="16:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7410" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7411" daytime="16:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7412" daytime="16:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7413" daytime="16:17" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1449" daytime="17:04" gender="M" number="25" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7915" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7916" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="7917" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7918" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5688" />
                    <RANKING order="2" place="2" resultid="4638" />
                    <RANKING order="3" place="3" resultid="4172" />
                    <RANKING order="4" place="-1" resultid="2696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7919" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3797" />
                    <RANKING order="2" place="2" resultid="2203" />
                    <RANKING order="3" place="3" resultid="3128" />
                    <RANKING order="4" place="4" resultid="2731" />
                    <RANKING order="5" place="5" resultid="2688" />
                    <RANKING order="6" place="-1" resultid="3815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7920" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5105" />
                    <RANKING order="2" place="2" resultid="3927" />
                    <RANKING order="3" place="3" resultid="2563" />
                    <RANKING order="4" place="4" resultid="2105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7921" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5554" />
                    <RANKING order="2" place="2" resultid="5285" />
                    <RANKING order="3" place="3" resultid="3767" />
                    <RANKING order="4" place="4" resultid="2477" />
                    <RANKING order="5" place="5" resultid="4839" />
                    <RANKING order="6" place="6" resultid="4656" />
                    <RANKING order="7" place="7" resultid="2760" />
                    <RANKING order="8" place="-1" resultid="6503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7922" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3856" />
                    <RANKING order="2" place="2" resultid="2433" />
                    <RANKING order="3" place="3" resultid="4800" />
                    <RANKING order="4" place="4" resultid="5731" />
                    <RANKING order="5" place="5" resultid="6037" />
                    <RANKING order="6" place="6" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7923" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6308" />
                    <RANKING order="2" place="2" resultid="5621" />
                    <RANKING order="3" place="3" resultid="4582" />
                    <RANKING order="4" place="4" resultid="4913" />
                    <RANKING order="5" place="5" resultid="3083" />
                    <RANKING order="6" place="6" resultid="2390" />
                    <RANKING order="7" place="7" resultid="3182" />
                    <RANKING order="8" place="8" resultid="4520" />
                    <RANKING order="9" place="9" resultid="6125" />
                    <RANKING order="10" place="10" resultid="2722" />
                    <RANKING order="11" place="11" resultid="4810" />
                    <RANKING order="12" place="12" resultid="2526" />
                    <RANKING order="13" place="-1" resultid="2871" />
                    <RANKING order="14" place="-1" resultid="6472" />
                    <RANKING order="15" place="-1" resultid="6490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7924" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4250" />
                    <RANKING order="2" place="2" resultid="2363" />
                    <RANKING order="3" place="3" resultid="6347" />
                    <RANKING order="4" place="4" resultid="3744" />
                    <RANKING order="5" place="5" resultid="4256" />
                    <RANKING order="6" place="6" resultid="4367" />
                    <RANKING order="7" place="7" resultid="3623" />
                    <RANKING order="8" place="8" resultid="3635" />
                    <RANKING order="9" place="9" resultid="3326" />
                    <RANKING order="10" place="10" resultid="3758" />
                    <RANKING order="11" place="11" resultid="5884" />
                    <RANKING order="12" place="12" resultid="2531" />
                    <RANKING order="13" place="13" resultid="4530" />
                    <RANKING order="14" place="14" resultid="5706" />
                    <RANKING order="15" place="15" resultid="6110" />
                    <RANKING order="16" place="16" resultid="5202" />
                    <RANKING order="17" place="17" resultid="5197" />
                    <RANKING order="18" place="-1" resultid="2251" />
                    <RANKING order="19" place="-1" resultid="5929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7925" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2995" />
                    <RANKING order="2" place="2" resultid="6383" />
                    <RANKING order="3" place="3" resultid="4931" />
                    <RANKING order="4" place="4" resultid="6374" />
                    <RANKING order="5" place="5" resultid="2903" />
                    <RANKING order="6" place="6" resultid="6046" />
                    <RANKING order="7" place="7" resultid="4962" />
                    <RANKING order="8" place="8" resultid="2011" />
                    <RANKING order="9" place="9" resultid="3022" />
                    <RANKING order="10" place="10" resultid="4697" />
                    <RANKING order="11" place="11" resultid="4626" />
                    <RANKING order="12" place="12" resultid="4709" />
                    <RANKING order="13" place="13" resultid="5717" />
                    <RANKING order="14" place="14" resultid="5009" />
                    <RANKING order="15" place="15" resultid="5016" />
                    <RANKING order="16" place="16" resultid="3422" />
                    <RANKING order="17" place="17" resultid="2057" />
                    <RANKING order="18" place="18" resultid="4317" />
                    <RANKING order="19" place="19" resultid="5027" />
                    <RANKING order="20" place="19" resultid="5630" />
                    <RANKING order="21" place="21" resultid="5041" />
                    <RANKING order="22" place="22" resultid="2069" />
                    <RANKING order="23" place="23" resultid="5257" />
                    <RANKING order="24" place="24" resultid="3142" />
                    <RANKING order="25" place="25" resultid="2257" />
                    <RANKING order="26" place="-1" resultid="2031" />
                    <RANKING order="27" place="-1" resultid="6009" />
                    <RANKING order="28" place="-1" resultid="6342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7926" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6428" />
                    <RANKING order="2" place="2" resultid="4734" />
                    <RANKING order="3" place="3" resultid="6019" />
                    <RANKING order="4" place="4" resultid="3721" />
                    <RANKING order="5" place="5" resultid="3194" />
                    <RANKING order="6" place="6" resultid="5048" />
                    <RANKING order="7" place="7" resultid="4178" />
                    <RANKING order="8" place="8" resultid="2380" />
                    <RANKING order="9" place="9" resultid="5207" />
                    <RANKING order="10" place="10" resultid="4991" />
                    <RANKING order="11" place="11" resultid="3590" />
                    <RANKING order="12" place="12" resultid="3431" />
                    <RANKING order="13" place="13" resultid="5217" />
                    <RANKING order="14" place="14" resultid="4943" />
                    <RANKING order="15" place="15" resultid="4506" />
                    <RANKING order="16" place="16" resultid="5238" />
                    <RANKING order="17" place="-1" resultid="2026" />
                    <RANKING order="18" place="-1" resultid="2450" />
                    <RANKING order="19" place="-1" resultid="2966" />
                    <RANKING order="20" place="-1" resultid="4683" />
                    <RANKING order="21" place="-1" resultid="6183" />
                    <RANKING order="22" place="-1" resultid="6866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7927" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4893" />
                    <RANKING order="2" place="2" resultid="2857" />
                    <RANKING order="3" place="3" resultid="2957" />
                    <RANKING order="4" place="4" resultid="3229" />
                    <RANKING order="5" place="5" resultid="3491" />
                    <RANKING order="6" place="6" resultid="2968" />
                    <RANKING order="7" place="7" resultid="2977" />
                    <RANKING order="8" place="7" resultid="4749" />
                    <RANKING order="9" place="9" resultid="2954" />
                    <RANKING order="10" place="10" resultid="4669" />
                    <RANKING order="11" place="11" resultid="5251" />
                    <RANKING order="12" place="12" resultid="6434" />
                    <RANKING order="13" place="13" resultid="4997" />
                    <RANKING order="14" place="14" resultid="2162" />
                    <RANKING order="15" place="15" resultid="6236" />
                    <RANKING order="16" place="16" resultid="2988" />
                    <RANKING order="17" place="17" resultid="4312" />
                    <RANKING order="18" place="18" resultid="2848" />
                    <RANKING order="19" place="19" resultid="2020" />
                    <RANKING order="20" place="-1" resultid="4677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7928" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4897" />
                    <RANKING order="2" place="2" resultid="3730" />
                    <RANKING order="3" place="3" resultid="5232" />
                    <RANKING order="4" place="4" resultid="6257" />
                    <RANKING order="5" place="5" resultid="5149" />
                    <RANKING order="6" place="6" resultid="2581" />
                    <RANKING order="7" place="7" resultid="5227" />
                    <RANKING order="8" place="8" resultid="2909" />
                    <RANKING order="9" place="9" resultid="2961" />
                    <RANKING order="10" place="10" resultid="2403" />
                    <RANKING order="11" place="11" resultid="6054" />
                    <RANKING order="12" place="12" resultid="3017" />
                    <RANKING order="13" place="13" resultid="4918" />
                    <RANKING order="14" place="14" resultid="5850" />
                    <RANKING order="15" place="15" resultid="6442" />
                    <RANKING order="16" place="16" resultid="3475" />
                    <RANKING order="17" place="17" resultid="3579" />
                    <RANKING order="18" place="18" resultid="2209" />
                    <RANKING order="19" place="-1" resultid="2190" />
                    <RANKING order="20" place="-1" resultid="4633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7929" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4204" />
                    <RANKING order="2" place="2" resultid="5190" />
                    <RANKING order="3" place="3" resultid="6362" />
                    <RANKING order="4" place="4" resultid="2137" />
                    <RANKING order="5" place="5" resultid="2613" />
                    <RANKING order="6" place="6" resultid="3825" />
                    <RANKING order="7" place="7" resultid="4513" />
                    <RANKING order="8" place="8" resultid="2662" />
                    <RANKING order="9" place="9" resultid="3895" />
                    <RANKING order="10" place="10" resultid="3479" />
                    <RANKING order="11" place="11" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7435" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7436" daytime="17:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7437" daytime="17:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7438" daytime="17:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7439" daytime="17:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7440" daytime="17:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7441" daytime="17:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7442" daytime="17:17" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7443" daytime="17:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7444" daytime="17:19" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7445" daytime="17:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7446" daytime="17:22" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7447" daytime="17:23" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7448" daytime="17:24" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7449" daytime="17:25" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7450" daytime="17:27" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7451" daytime="17:28" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1529" daytime="19:34" gender="F" number="30" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7856" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7857" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3818" />
                    <RANKING order="2" place="2" resultid="4140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7858" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7859" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3317" />
                    <RANKING order="2" place="2" resultid="5157" />
                    <RANKING order="3" place="3" resultid="2947" />
                    <RANKING order="4" place="-1" resultid="6407" />
                    <RANKING order="5" place="-1" resultid="4034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7860" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4751" />
                    <RANKING order="2" place="2" resultid="6268" />
                    <RANKING order="3" place="3" resultid="4547" />
                    <RANKING order="4" place="4" resultid="5062" />
                    <RANKING order="5" place="5" resultid="4457" />
                    <RANKING order="6" place="6" resultid="4349" />
                    <RANKING order="7" place="-1" resultid="3318" />
                    <RANKING order="8" place="-1" resultid="5657" />
                    <RANKING order="9" place="-1" resultid="6477" />
                    <RANKING order="10" place="-1" resultid="3601" />
                    <RANKING order="11" place="-1" resultid="5516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7861" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2788" />
                    <RANKING order="2" place="2" resultid="3600" />
                    <RANKING order="3" place="-1" resultid="3035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7862" agemax="99" agemin="80" name="0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3602" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7489" daytime="19:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7490" daytime="19:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7491" daytime="19:42" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1513" daytime="18:43" gender="M" number="29" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7975" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="7976" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7977" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="7978" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4173" />
                    <RANKING order="2" place="2" resultid="4817" />
                    <RANKING order="3" place="3" resultid="2705" />
                    <RANKING order="4" place="-1" resultid="5177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7979" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4783" />
                    <RANKING order="2" place="2" resultid="2099" />
                    <RANKING order="3" place="3" resultid="3935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7980" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3928" />
                    <RANKING order="2" place="2" resultid="3138" />
                    <RANKING order="3" place="3" resultid="2106" />
                    <RANKING order="4" place="4" resultid="2303" />
                    <RANKING order="5" place="-1" resultid="2092" />
                    <RANKING order="6" place="-1" resultid="5680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7981" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3261" />
                    <RANKING order="2" place="2" resultid="6504" />
                    <RANKING order="3" place="3" resultid="2840" />
                    <RANKING order="4" place="4" resultid="5865" />
                    <RANKING order="5" place="5" resultid="4160" />
                    <RANKING order="6" place="6" resultid="4657" />
                    <RANKING order="7" place="7" resultid="3243" />
                    <RANKING order="8" place="8" resultid="3151" />
                    <RANKING order="9" place="9" resultid="4847" />
                    <RANKING order="10" place="-1" resultid="3216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7982" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4391" />
                    <RANKING order="2" place="2" resultid="5184" />
                    <RANKING order="3" place="3" resultid="6002" />
                    <RANKING order="4" place="4" resultid="5732" />
                    <RANKING order="5" place="5" resultid="6118" />
                    <RANKING order="6" place="-1" resultid="3122" />
                    <RANKING order="7" place="-1" resultid="4620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7983" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5638" />
                    <RANKING order="2" place="2" resultid="4914" />
                    <RANKING order="3" place="3" resultid="5755" />
                    <RANKING order="4" place="4" resultid="5994" />
                    <RANKING order="5" place="5" resultid="5822" />
                    <RANKING order="6" place="6" resultid="4574" />
                    <RANKING order="7" place="7" resultid="4292" />
                    <RANKING order="8" place="-1" resultid="2003" />
                    <RANKING order="9" place="-1" resultid="2294" />
                    <RANKING order="10" place="-1" resultid="5525" />
                    <RANKING order="11" place="-1" resultid="6473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7984" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4560" />
                    <RANKING order="2" place="2" resultid="2364" />
                    <RANKING order="3" place="3" resultid="6149" />
                    <RANKING order="4" place="4" resultid="4264" />
                    <RANKING order="5" place="5" resultid="3687" />
                    <RANKING order="6" place="6" resultid="3401" />
                    <RANKING order="7" place="7" resultid="6197" />
                    <RANKING order="8" place="8" resultid="3759" />
                    <RANKING order="9" place="9" resultid="3678" />
                    <RANKING order="10" place="10" resultid="5707" />
                    <RANKING order="11" place="11" resultid="6111" />
                    <RANKING order="12" place="12" resultid="2808" />
                    <RANKING order="13" place="13" resultid="2532" />
                    <RANKING order="14" place="14" resultid="4531" />
                    <RANKING order="15" place="15" resultid="5724" />
                    <RANKING order="16" place="16" resultid="3060" />
                    <RANKING order="17" place="17" resultid="4429" />
                    <RANKING order="18" place="18" resultid="5930" />
                    <RANKING order="19" place="19" resultid="3997" />
                    <RANKING order="20" place="-1" resultid="5773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7985" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2047" />
                    <RANKING order="2" place="2" resultid="6010" />
                    <RANKING order="3" place="3" resultid="3204" />
                    <RANKING order="4" place="4" resultid="4627" />
                    <RANKING order="5" place="5" resultid="6140" />
                    <RANKING order="6" place="6" resultid="4932" />
                    <RANKING order="7" place="7" resultid="5718" />
                    <RANKING order="8" place="8" resultid="4710" />
                    <RANKING order="9" place="9" resultid="5010" />
                    <RANKING order="10" place="10" resultid="5099" />
                    <RANKING order="11" place="11" resultid="4883" />
                    <RANKING order="12" place="12" resultid="4555" />
                    <RANKING order="13" place="13" resultid="3255" />
                    <RANKING order="14" place="14" resultid="3621" />
                    <RANKING order="15" place="15" resultid="2070" />
                    <RANKING order="16" place="16" resultid="4910" />
                    <RANKING order="17" place="17" resultid="5258" />
                    <RANKING order="18" place="18" resultid="4535" />
                    <RANKING order="19" place="-1" resultid="3048" />
                    <RANKING order="20" place="-1" resultid="3423" />
                    <RANKING order="21" place="-1" resultid="5028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7986" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4423" />
                    <RANKING order="2" place="2" resultid="4591" />
                    <RANKING order="3" place="3" resultid="6095" />
                    <RANKING order="4" place="4" resultid="6026" />
                    <RANKING order="5" place="5" resultid="6184" />
                    <RANKING order="6" place="6" resultid="2381" />
                    <RANKING order="7" place="7" resultid="5789" />
                    <RANKING order="8" place="8" resultid="5223" />
                    <RANKING order="9" place="9" resultid="2545" />
                    <RANKING order="10" place="10" resultid="5239" />
                    <RANKING order="11" place="11" resultid="4507" />
                    <RANKING order="12" place="12" resultid="3550" />
                    <RANKING order="13" place="13" resultid="6867" />
                    <RANKING order="14" place="-1" resultid="4331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7987" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2132" />
                    <RANKING order="2" place="2" resultid="2978" />
                    <RANKING order="3" place="3" resultid="4399" />
                    <RANKING order="4" place="4" resultid="3492" />
                    <RANKING order="5" place="5" resultid="2858" />
                    <RANKING order="6" place="6" resultid="4750" />
                    <RANKING order="7" place="7" resultid="6435" />
                    <RANKING order="8" place="8" resultid="4678" />
                    <RANKING order="9" place="9" resultid="2152" />
                    <RANKING order="10" place="10" resultid="5917" />
                    <RANKING order="11" place="11" resultid="3268" />
                    <RANKING order="12" place="12" resultid="2849" />
                    <RANKING order="13" place="-1" resultid="6368" />
                    <RANKING order="14" place="-1" resultid="3438" />
                    <RANKING order="15" place="-1" resultid="3544" />
                    <RANKING order="16" place="-1" resultid="4894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7988" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8231" />
                    <RANKING order="2" place="2" resultid="5793" />
                    <RANKING order="3" place="3" resultid="3731" />
                    <RANKING order="4" place="4" resultid="6176" />
                    <RANKING order="5" place="5" resultid="6352" />
                    <RANKING order="6" place="6" resultid="6258" />
                    <RANKING order="7" place="7" resultid="2177" />
                    <RANKING order="8" place="8" resultid="6055" />
                    <RANKING order="9" place="9" resultid="5851" />
                    <RANKING order="10" place="10" resultid="4919" />
                    <RANKING order="11" place="-1" resultid="2185" />
                    <RANKING order="12" place="-1" resultid="2520" />
                    <RANKING order="13" place="-1" resultid="3583" />
                    <RANKING order="14" place="-1" resultid="5150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7989" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5191" />
                    <RANKING order="2" place="2" resultid="4189" />
                    <RANKING order="3" place="3" resultid="3826" />
                    <RANKING order="4" place="4" resultid="2614" />
                    <RANKING order="5" place="5" resultid="2138" />
                    <RANKING order="6" place="6" resultid="4514" />
                    <RANKING order="7" place="7" resultid="3979" />
                    <RANKING order="8" place="-1" resultid="2321" />
                    <RANKING order="9" place="-1" resultid="3848" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7475" daytime="18:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7476" daytime="18:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7477" daytime="18:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7478" daytime="18:59" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7479" daytime="19:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7480" daytime="19:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7481" daytime="19:09" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7482" daytime="19:13" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7483" daytime="19:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7484" daytime="19:19" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7485" daytime="19:22" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7486" daytime="19:25" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7487" daytime="19:28" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7488" daytime="19:31" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-11-17" daytime="09:00" endtime="13:57" name="Zimowe Mistrzostwa Polskiw Pływaniu Masters BLOK IV" number="4" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1673" daytime="10:49" gender="F" number="38" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8080" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8081" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="8082" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8083" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8084" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8085" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5965" />
                    <RANKING order="2" place="2" resultid="4094" />
                    <RANKING order="3" place="3" resultid="3775" />
                    <RANKING order="4" place="4" resultid="2352" />
                    <RANKING order="5" place="5" resultid="2077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8086" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6488" />
                    <RANKING order="2" place="2" resultid="4828" />
                    <RANKING order="3" place="3" resultid="4119" />
                    <RANKING order="4" place="4" resultid="4153" />
                    <RANKING order="5" place="5" resultid="2268" />
                    <RANKING order="6" place="6" resultid="3985" />
                    <RANKING order="7" place="7" resultid="2594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8087" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                    <RANKING order="2" place="2" resultid="6333" />
                    <RANKING order="3" place="3" resultid="5550" />
                    <RANKING order="4" place="4" resultid="5979" />
                    <RANKING order="5" place="5" resultid="5132" />
                    <RANKING order="6" place="6" resultid="4080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8088" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3093" />
                    <RANKING order="2" place="2" resultid="2375" />
                    <RANKING order="3" place="3" resultid="4272" />
                    <RANKING order="4" place="4" resultid="2275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8089" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3165" />
                    <RANKING order="2" place="2" resultid="4326" />
                    <RANKING order="3" place="3" resultid="3804" />
                    <RANKING order="4" place="4" resultid="4704" />
                    <RANKING order="5" place="5" resultid="2085" />
                    <RANKING order="6" place="6" resultid="4376" />
                    <RANKING order="7" place="7" resultid="5117" />
                    <RANKING order="8" place="-1" resultid="5092" />
                    <RANKING order="9" place="-1" resultid="6216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8090" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2600" />
                    <RANKING order="2" place="2" resultid="3178" />
                    <RANKING order="3" place="3" resultid="3303" />
                    <RANKING order="4" place="4" resultid="3671" />
                    <RANKING order="5" place="5" resultid="2936" />
                    <RANKING order="6" place="6" resultid="4501" />
                    <RANKING order="7" place="7" resultid="5515" />
                    <RANKING order="8" place="8" resultid="3696" />
                    <RANKING order="9" place="9" resultid="5265" />
                    <RANKING order="10" place="10" resultid="5644" />
                    <RANKING order="11" place="11" resultid="3961" />
                    <RANKING order="12" place="12" resultid="5950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8091" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2819" />
                    <RANKING order="2" place="2" resultid="3714" />
                    <RANKING order="3" place="3" resultid="4419" />
                    <RANKING order="4" place="4" resultid="4957" />
                    <RANKING order="5" place="5" resultid="4949" />
                    <RANKING order="6" place="6" resultid="4595" />
                    <RANKING order="7" place="7" resultid="5614" />
                    <RANKING order="8" place="8" resultid="3389" />
                    <RANKING order="9" place="-1" resultid="4029" />
                    <RANKING order="10" place="-1" resultid="5649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8092" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3706" />
                    <RANKING order="2" place="2" resultid="4043" />
                    <RANKING order="3" place="3" resultid="5246" />
                    <RANKING order="4" place="4" resultid="3523" />
                    <RANKING order="5" place="5" resultid="3752" />
                    <RANKING order="6" place="6" resultid="3394" />
                    <RANKING order="7" place="7" resultid="6465" />
                    <RANKING order="8" place="8" resultid="4477" />
                    <RANKING order="9" place="-1" resultid="3008" />
                    <RANKING order="10" place="-1" resultid="3519" />
                    <RANKING order="11" place="-1" resultid="3883" />
                    <RANKING order="12" place="-1" resultid="4542" />
                    <RANKING order="13" place="-1" resultid="5212" />
                    <RANKING order="14" place="-1" resultid="5538" />
                    <RANKING order="15" place="-1" resultid="3116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8093" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                    <RANKING order="2" place="2" resultid="2040" />
                    <RANKING order="3" place="3" resultid="3467" />
                    <RANKING order="4" place="4" resultid="5123" />
                    <RANKING order="5" place="5" resultid="4381" />
                    <RANKING order="6" place="6" resultid="3298" />
                    <RANKING order="7" place="-1" resultid="2918" />
                    <RANKING order="8" place="-1" resultid="5269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8094" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5987" />
                    <RANKING order="2" place="2" resultid="2181" />
                    <RANKING order="3" place="3" resultid="2625" />
                    <RANKING order="4" place="4" resultid="2226" />
                    <RANKING order="5" place="5" resultid="3841" />
                    <RANKING order="6" place="6" resultid="4021" />
                    <RANKING order="7" place="7" resultid="2679" />
                    <RANKING order="8" place="-1" resultid="5302" />
                    <RANKING order="9" place="-1" resultid="5909" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7537" daytime="10:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7538" daytime="10:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7539" daytime="10:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7540" daytime="10:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7541" daytime="10:57" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7542" daytime="10:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7543" daytime="11:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7544" daytime="11:01" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7545" daytime="11:02" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1641" daytime="09:39" gender="F" number="36" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8050" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8051" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8052" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8053" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="8054" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8055" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3792" />
                    <RANKING order="2" place="2" resultid="4168" />
                    <RANKING order="3" place="3" resultid="4133" />
                    <RANKING order="4" place="4" resultid="2076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8056" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3449" />
                    <RANKING order="2" place="2" resultid="3812" />
                    <RANKING order="3" place="3" resultid="3913" />
                    <RANKING order="4" place="4" resultid="5296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8057" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4227" />
                    <RANKING order="2" place="2" resultid="3109" />
                    <RANKING order="3" place="3" resultid="5131" />
                    <RANKING order="4" place="4" resultid="4062" />
                    <RANKING order="5" place="5" resultid="5978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8058" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2557" />
                    <RANKING order="2" place="2" resultid="6245" />
                    <RANKING order="3" place="3" resultid="5957" />
                    <RANKING order="4" place="4" resultid="2274" />
                    <RANKING order="5" place="5" resultid="6206" />
                    <RANKING order="6" place="-1" resultid="2945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8059" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3159" />
                    <RANKING order="2" place="2" resultid="2356" />
                    <RANKING order="3" place="3" resultid="3921" />
                    <RANKING order="4" place="4" resultid="5893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8060" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3177" />
                    <RANKING order="2" place="2" resultid="5562" />
                    <RANKING order="3" place="3" resultid="3076" />
                    <RANKING order="4" place="4" resultid="5112" />
                    <RANKING order="5" place="5" resultid="4304" />
                    <RANKING order="6" place="6" resultid="6169" />
                    <RANKING order="7" place="7" resultid="4981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8061" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4489" />
                    <RANKING order="2" place="2" resultid="6231" />
                    <RANKING order="3" place="3" resultid="2399" />
                    <RANKING order="4" place="4" resultid="4010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8062" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3007" />
                    <RANKING order="2" place="2" resultid="5581" />
                    <RANKING order="3" place="3" resultid="2826" />
                    <RANKING order="4" place="4" resultid="4613" />
                    <RANKING order="5" place="-1" resultid="3518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8063" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3874" />
                    <RANKING order="2" place="2" resultid="4690" />
                    <RANKING order="3" place="3" resultid="4722" />
                    <RANKING order="4" place="4" resultid="5499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8064" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4198" />
                    <RANKING order="2" place="2" resultid="2333" />
                    <RANKING order="3" place="3" resultid="4020" />
                    <RANKING order="4" place="-1" resultid="3273" />
                    <RANKING order="5" place="-1" resultid="4218" />
                    <RANKING order="6" place="-1" resultid="5908" />
                    <RANKING order="7" place="-1" resultid="5970" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7523" daytime="09:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7524" daytime="09:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7525" daytime="09:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7526" daytime="09:59" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7527" daytime="10:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7528" daytime="10:08" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1689" daytime="11:04" gender="M" number="39" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8095" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8096" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2247" />
                    <RANKING order="2" place="-1" resultid="2896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8097" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4106" />
                    <RANKING order="2" place="-1" resultid="4569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8098" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4640" />
                    <RANKING order="2" place="2" resultid="5691" />
                    <RANKING order="3" place="3" resultid="2642" />
                    <RANKING order="4" place="4" resultid="2699" />
                    <RANKING order="5" place="5" resultid="2511" />
                    <RANKING order="6" place="6" resultid="4818" />
                    <RANKING order="7" place="7" resultid="2707" />
                    <RANKING order="8" place="-1" resultid="5179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8099" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3101" />
                    <RANKING order="2" place="2" resultid="2206" />
                    <RANKING order="3" place="3" resultid="3798" />
                    <RANKING order="4" place="4" resultid="3951" />
                    <RANKING order="5" place="5" resultid="2690" />
                    <RANKING order="6" place="6" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8100" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4729" />
                    <RANKING order="2" place="2" resultid="4071" />
                    <RANKING order="3" place="3" resultid="2564" />
                    <RANKING order="4" place="4" resultid="2767" />
                    <RANKING order="5" place="5" resultid="4112" />
                    <RANKING order="6" place="6" resultid="5936" />
                    <RANKING order="7" place="7" resultid="3251" />
                    <RANKING order="8" place="-1" resultid="3655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8101" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5533" />
                    <RANKING order="2" place="2" resultid="2478" />
                    <RANKING order="3" place="3" resultid="3191" />
                    <RANKING order="4" place="4" resultid="2122" />
                    <RANKING order="5" place="5" resultid="4607" />
                    <RANKING order="6" place="6" resultid="4841" />
                    <RANKING order="7" place="7" resultid="4849" />
                    <RANKING order="8" place="-1" resultid="5815" />
                    <RANKING order="9" place="-1" resultid="3146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8102" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2415" />
                    <RANKING order="2" place="2" resultid="3414" />
                    <RANKING order="3" place="3" resultid="2436" />
                    <RANKING order="4" place="4" resultid="5653" />
                    <RANKING order="5" place="5" resultid="4803" />
                    <RANKING order="6" place="6" resultid="6033" />
                    <RANKING order="7" place="7" resultid="2573" />
                    <RANKING order="8" place="8" resultid="3291" />
                    <RANKING order="9" place="9" resultid="3123" />
                    <RANKING order="10" place="-1" resultid="4360" />
                    <RANKING order="11" place="-1" resultid="4621" />
                    <RANKING order="12" place="-1" resultid="5186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8103" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3013" />
                    <RANKING order="2" place="2" resultid="6310" />
                    <RANKING order="3" place="3" resultid="2295" />
                    <RANKING order="4" place="4" resultid="3223" />
                    <RANKING order="5" place="5" resultid="3085" />
                    <RANKING order="6" place="6" resultid="5879" />
                    <RANKING order="7" place="7" resultid="4811" />
                    <RANKING order="8" place="8" resultid="6127" />
                    <RANKING order="9" place="9" resultid="6251" />
                    <RANKING order="10" place="10" resultid="4521" />
                    <RANKING order="11" place="11" resultid="2873" />
                    <RANKING order="12" place="12" resultid="4293" />
                    <RANKING order="13" place="13" resultid="2725" />
                    <RANKING order="14" place="14" resultid="4575" />
                    <RANKING order="15" place="15" resultid="3969" />
                    <RANKING order="16" place="16" resultid="5143" />
                    <RANKING order="17" place="17" resultid="2236" />
                    <RANKING order="18" place="-1" resultid="2168" />
                    <RANKING order="19" place="-1" resultid="5823" />
                    <RANKING order="20" place="-1" resultid="6475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8104" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4265" />
                    <RANKING order="2" place="2" resultid="3663" />
                    <RANKING order="3" place="3" resultid="4257" />
                    <RANKING order="4" place="4" resultid="6348" />
                    <RANKING order="5" place="5" resultid="3689" />
                    <RANKING order="6" place="6" resultid="4370" />
                    <RANKING order="7" place="7" resultid="2810" />
                    <RANKING order="8" place="8" resultid="4533" />
                    <RANKING order="9" place="9" resultid="4005" />
                    <RANKING order="10" place="10" resultid="3134" />
                    <RANKING order="11" place="11" resultid="3998" />
                    <RANKING order="12" place="-1" resultid="2252" />
                    <RANKING order="13" place="-1" resultid="4430" />
                    <RANKING order="14" place="-1" resultid="5708" />
                    <RANKING order="15" place="-1" resultid="5833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8105" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4699" />
                    <RANKING order="2" place="2" resultid="3206" />
                    <RANKING order="3" place="3" resultid="6375" />
                    <RANKING order="4" place="4" resultid="6049" />
                    <RANKING order="5" place="5" resultid="2904" />
                    <RANKING order="6" place="6" resultid="6190" />
                    <RANKING order="7" place="7" resultid="5100" />
                    <RANKING order="8" place="8" resultid="4963" />
                    <RANKING order="9" place="9" resultid="4318" />
                    <RANKING order="10" place="10" resultid="5925" />
                    <RANKING order="11" place="11" resultid="2013" />
                    <RANKING order="12" place="12" resultid="6388" />
                    <RANKING order="13" place="13" resultid="5017" />
                    <RANKING order="14" place="14" resultid="3045" />
                    <RANKING order="15" place="15" resultid="2060" />
                    <RANKING order="16" place="16" resultid="5633" />
                    <RANKING order="17" place="17" resultid="3256" />
                    <RANKING order="18" place="18" resultid="5042" />
                    <RANKING order="19" place="19" resultid="4985" />
                    <RANKING order="20" place="20" resultid="3051" />
                    <RANKING order="21" place="21" resultid="5259" />
                    <RANKING order="22" place="22" resultid="2493" />
                    <RANKING order="23" place="23" resultid="4834" />
                    <RANKING order="24" place="24" resultid="2260" />
                    <RANKING order="25" place="-1" resultid="1998" />
                    <RANKING order="26" place="-1" resultid="2742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8106" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6020" />
                    <RANKING order="2" place="2" resultid="6430" />
                    <RANKING order="3" place="3" resultid="4737" />
                    <RANKING order="4" place="4" resultid="3481" />
                    <RANKING order="5" place="5" resultid="5049" />
                    <RANKING order="6" place="6" resultid="6096" />
                    <RANKING order="7" place="7" resultid="4937" />
                    <RANKING order="8" place="8" resultid="5056" />
                    <RANKING order="9" place="9" resultid="4992" />
                    <RANKING order="10" place="10" resultid="3419" />
                    <RANKING order="11" place="11" resultid="4973" />
                    <RANKING order="12" place="12" resultid="5053" />
                    <RANKING order="13" place="13" resultid="5036" />
                    <RANKING order="14" place="-1" resultid="2382" />
                    <RANKING order="15" place="-1" resultid="2452" />
                    <RANKING order="16" place="-1" resultid="4508" />
                    <RANKING order="17" place="-1" resultid="4889" />
                    <RANKING order="18" place="-1" resultid="5591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8107" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4287" />
                    <RANKING order="2" place="2" resultid="3231" />
                    <RANKING order="3" place="3" resultid="5999" />
                    <RANKING order="4" place="4" resultid="4245" />
                    <RANKING order="5" place="5" resultid="4679" />
                    <RANKING order="6" place="6" resultid="2164" />
                    <RANKING order="7" place="-1" resultid="2021" />
                    <RANKING order="8" place="-1" resultid="2214" />
                    <RANKING order="9" place="-1" resultid="3439" />
                    <RANKING order="10" place="-1" resultid="4471" />
                    <RANKING order="11" place="-1" resultid="6237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8108" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2910" />
                    <RANKING order="2" place="2" resultid="2962" />
                    <RANKING order="3" place="3" resultid="2408" />
                    <RANKING order="4" place="4" resultid="6443" />
                    <RANKING order="5" place="5" resultid="4480" />
                    <RANKING order="6" place="-1" resultid="2191" />
                    <RANKING order="7" place="-1" resultid="2341" />
                    <RANKING order="8" place="-1" resultid="3461" />
                    <RANKING order="9" place="-1" resultid="3568" />
                    <RANKING order="10" place="-1" resultid="5902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8109" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4206" />
                    <RANKING order="2" place="2" resultid="4190" />
                    <RANKING order="3" place="3" resultid="3849" />
                    <RANKING order="4" place="4" resultid="2157" />
                    <RANKING order="5" place="5" resultid="2631" />
                    <RANKING order="6" place="6" resultid="2664" />
                    <RANKING order="7" place="7" resultid="2140" />
                    <RANKING order="8" place="8" resultid="3980" />
                    <RANKING order="9" place="-1" resultid="2323" />
                    <RANKING order="10" place="-1" resultid="3831" />
                    <RANKING order="11" place="-1" resultid="5744" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7546" daytime="11:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7547" daytime="11:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7548" daytime="11:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7549" daytime="11:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7550" daytime="11:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7551" daytime="11:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7552" daytime="11:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7553" daytime="11:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7554" daytime="11:17" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7555" daytime="11:19" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7556" daytime="11:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7557" daytime="11:21" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7558" daytime="11:23" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7559" daytime="11:24" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7560" daytime="11:25" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7561" daytime="11:27" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1625" daytime="09:13" gender="M" number="35" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8035" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8036" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="8037" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8038" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4639" />
                    <RANKING order="2" place="2" resultid="2641" />
                    <RANKING order="3" place="3" resultid="2698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8039" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2205" />
                    <RANKING order="2" place="2" resultid="3129" />
                    <RANKING order="3" place="3" resultid="4785" />
                    <RANKING order="4" place="4" resultid="5170" />
                    <RANKING order="5" place="5" resultid="2425" />
                    <RANKING order="6" place="6" resultid="2733" />
                    <RANKING order="7" place="7" resultid="3937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8040" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5106" />
                    <RANKING order="2" place="2" resultid="3929" />
                    <RANKING order="3" place="3" resultid="2715" />
                    <RANKING order="4" place="4" resultid="2766" />
                    <RANKING order="5" place="-1" resultid="4111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8041" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5555" />
                    <RANKING order="2" place="2" resultid="3190" />
                    <RANKING order="3" place="3" resultid="2121" />
                    <RANKING order="4" place="4" resultid="5866" />
                    <RANKING order="5" place="5" resultid="4840" />
                    <RANKING order="6" place="6" resultid="2761" />
                    <RANKING order="7" place="7" resultid="3245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8042" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2435" />
                    <RANKING order="2" place="2" resultid="4802" />
                    <RANKING order="3" place="3" resultid="5185" />
                    <RANKING order="4" place="4" resultid="5598" />
                    <RANKING order="5" place="5" resultid="2572" />
                    <RANKING order="6" place="6" resultid="6103" />
                    <RANKING order="7" place="7" resultid="6039" />
                    <RANKING order="8" place="-1" resultid="2222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8043" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5623" />
                    <RANKING order="2" place="2" resultid="6309" />
                    <RANKING order="3" place="3" resultid="4584" />
                    <RANKING order="4" place="4" resultid="4915" />
                    <RANKING order="5" place="5" resultid="3084" />
                    <RANKING order="6" place="6" resultid="2392" />
                    <RANKING order="7" place="7" resultid="6126" />
                    <RANKING order="8" place="8" resultid="2872" />
                    <RANKING order="9" place="9" resultid="2724" />
                    <RANKING order="10" place="-1" resultid="2005" />
                    <RANKING order="11" place="-1" resultid="2527" />
                    <RANKING order="12" place="-1" resultid="6474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8044" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2365" />
                    <RANKING order="2" place="2" resultid="6151" />
                    <RANKING order="3" place="3" resultid="4251" />
                    <RANKING order="4" place="4" resultid="4369" />
                    <RANKING order="5" place="5" resultid="3688" />
                    <RANKING order="6" place="6" resultid="3760" />
                    <RANKING order="7" place="7" resultid="4532" />
                    <RANKING order="8" place="8" resultid="2533" />
                    <RANKING order="9" place="-1" resultid="3624" />
                    <RANKING order="10" place="-1" resultid="5931" />
                    <RANKING order="11" place="-1" resultid="6112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8045" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2997" />
                    <RANKING order="2" place="2" resultid="6384" />
                    <RANKING order="3" place="3" resultid="4933" />
                    <RANKING order="4" place="4" resultid="2049" />
                    <RANKING order="5" place="5" resultid="6011" />
                    <RANKING order="6" place="6" resultid="2012" />
                    <RANKING order="7" place="7" resultid="2883" />
                    <RANKING order="8" place="8" resultid="3000" />
                    <RANKING order="9" place="9" resultid="4698" />
                    <RANKING order="10" place="10" resultid="5632" />
                    <RANKING order="11" place="11" resultid="4556" />
                    <RANKING order="12" place="12" resultid="2259" />
                    <RANKING order="13" place="-1" resultid="3205" />
                    <RANKING order="14" place="-1" resultid="3424" />
                    <RANKING order="15" place="-1" resultid="5029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8046" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6429" />
                    <RANKING order="2" place="2" resultid="3723" />
                    <RANKING order="3" place="3" resultid="4736" />
                    <RANKING order="4" place="4" resultid="3196" />
                    <RANKING order="5" place="5" resultid="4180" />
                    <RANKING order="6" place="6" resultid="3432" />
                    <RANKING order="7" place="7" resultid="6027" />
                    <RANKING order="8" place="8" resultid="4944" />
                    <RANKING order="9" place="-1" resultid="2451" />
                    <RANKING order="10" place="-1" resultid="5590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8047" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3230" />
                    <RANKING order="2" place="2" resultid="2133" />
                    <RANKING order="3" place="3" resultid="2970" />
                    <RANKING order="4" place="4" resultid="2859" />
                    <RANKING order="5" place="5" resultid="3493" />
                    <RANKING order="6" place="6" resultid="4671" />
                    <RANKING order="7" place="7" resultid="2163" />
                    <RANKING order="8" place="8" resultid="6436" />
                    <RANKING order="9" place="9" resultid="2850" />
                    <RANKING order="10" place="-1" resultid="5488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8048" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3732" />
                    <RANKING order="2" place="2" resultid="6178" />
                    <RANKING order="3" place="3" resultid="5234" />
                    <RANKING order="4" place="4" resultid="2582" />
                    <RANKING order="5" place="5" resultid="5151" />
                    <RANKING order="6" place="6" resultid="5228" />
                    <RANKING order="7" place="7" resultid="3512" />
                    <RANKING order="8" place="8" resultid="6056" />
                    <RANKING order="9" place="-1" resultid="2186" />
                    <RANKING order="10" place="-1" resultid="4898" />
                    <RANKING order="11" place="-1" resultid="5945" />
                    <RANKING order="12" place="-1" resultid="6259" />
                    <RANKING order="13" place="-1" resultid="8162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8049" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4205" />
                    <RANKING order="2" place="2" resultid="6363" />
                    <RANKING order="3" place="3" resultid="2139" />
                    <RANKING order="4" place="4" resultid="2615" />
                    <RANKING order="5" place="5" resultid="4515" />
                    <RANKING order="6" place="6" resultid="3896" />
                    <RANKING order="7" place="7" resultid="2663" />
                    <RANKING order="8" place="-1" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7512" daytime="09:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7513" daytime="09:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7514" daytime="09:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7515" daytime="09:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7516" daytime="09:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7517" daytime="09:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7518" daytime="09:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7519" daytime="09:31" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7520" daytime="09:33" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7521" daytime="09:35" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7522" daytime="09:37" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1657" daytime="10:12" gender="M" number="37" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8065" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8066" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8067" agemax="84" agemin="80" name="L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4105" />
                    <RANKING order="2" place="-1" resultid="4568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8068" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5690" />
                    <RANKING order="2" place="2" resultid="3944" />
                    <RANKING order="3" place="3" resultid="2510" />
                    <RANKING order="4" place="4" resultid="2706" />
                    <RANKING order="5" place="-1" resultid="5178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8069" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3100" />
                    <RANKING order="2" place="2" resultid="2457" />
                    <RANKING order="3" place="3" resultid="3785" />
                    <RANKING order="4" place="4" resultid="2426" />
                    <RANKING order="5" place="5" resultid="2689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8070" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4601" />
                    <RANKING order="2" place="2" resultid="2716" />
                    <RANKING order="3" place="3" resultid="5782" />
                    <RANKING order="4" place="4" resultid="2304" />
                    <RANKING order="5" place="-1" resultid="3654" />
                    <RANKING order="6" place="-1" resultid="5681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8071" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5287" />
                    <RANKING order="2" place="2" resultid="3217" />
                    <RANKING order="3" place="3" resultid="5699" />
                    <RANKING order="4" place="4" resultid="2841" />
                    <RANKING order="5" place="5" resultid="3769" />
                    <RANKING order="6" place="6" resultid="4161" />
                    <RANKING order="7" place="7" resultid="2754" />
                    <RANKING order="8" place="8" resultid="3246" />
                    <RANKING order="9" place="9" resultid="4848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8072" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3858" />
                    <RANKING order="2" place="2" resultid="2346" />
                    <RANKING order="3" place="3" resultid="6119" />
                    <RANKING order="4" place="4" resultid="6040" />
                    <RANKING order="5" place="5" resultid="3282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8073" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4925" />
                    <RANKING order="2" place="2" resultid="4585" />
                    <RANKING order="3" place="3" resultid="5995" />
                    <RANKING order="4" place="4" resultid="2802" />
                    <RANKING order="5" place="5" resultid="5526" />
                    <RANKING order="6" place="6" resultid="2467" />
                    <RANKING order="7" place="7" resultid="5086" />
                    <RANKING order="8" place="8" resultid="3968" />
                    <RANKING order="9" place="-1" resultid="4278" />
                    <RANKING order="10" place="-1" resultid="5624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8074" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3746" />
                    <RANKING order="2" place="2" resultid="2366" />
                    <RANKING order="3" place="3" resultid="2672" />
                    <RANKING order="4" place="4" resultid="4389" />
                    <RANKING order="5" place="5" resultid="5079" />
                    <RANKING order="6" place="6" resultid="6198" />
                    <RANKING order="7" place="7" resultid="3679" />
                    <RANKING order="8" place="-1" resultid="3402" />
                    <RANKING order="9" place="-1" resultid="5774" />
                    <RANKING order="10" place="-1" resultid="5832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8075" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6048" />
                    <RANKING order="2" place="2" resultid="6142" />
                    <RANKING order="3" place="3" resultid="3001" />
                    <RANKING order="4" place="4" resultid="2059" />
                    <RANKING order="5" place="5" resultid="5924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8076" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3724" />
                    <RANKING order="2" place="2" resultid="3197" />
                    <RANKING order="3" place="3" resultid="3890" />
                    <RANKING order="4" place="4" resultid="2546" />
                    <RANKING order="5" place="5" resultid="4972" />
                    <RANKING order="6" place="-1" resultid="5240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8077" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5859" />
                    <RANKING order="2" place="2" resultid="3501" />
                    <RANKING order="3" place="3" resultid="5252" />
                    <RANKING order="4" place="4" resultid="4401" />
                    <RANKING order="5" place="5" resultid="4715" />
                    <RANKING order="6" place="6" resultid="3866" />
                    <RANKING order="7" place="-1" resultid="4672" />
                    <RANKING order="8" place="-1" resultid="5489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8078" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6179" />
                    <RANKING order="2" place="2" resultid="2286" />
                    <RANKING order="3" place="3" resultid="6353" />
                    <RANKING order="4" place="-1" resultid="2340" />
                    <RANKING order="5" place="-1" resultid="3460" />
                    <RANKING order="6" place="-1" resultid="5901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8079" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2322" />
                    <RANKING order="2" place="2" resultid="4212" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7529" daytime="10:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7530" daytime="10:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7531" daytime="10:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7532" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7533" daytime="10:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7534" daytime="10:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7535" daytime="10:41" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7536" daytime="10:45" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1737" daytime="12:39" gender="M" number="42" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8125" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8126" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="8127" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8128" agemax="79" agemin="75" name="K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4174" />
                    <RANKING order="2" place="2" resultid="4819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8129" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4786" />
                    <RANKING order="2" place="2" resultid="2100" />
                    <RANKING order="3" place="3" resultid="2734" />
                    <RANKING order="4" place="-1" resultid="3938" />
                    <RANKING order="5" place="-1" resultid="5171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8130" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5783" />
                    <RANKING order="2" place="2" resultid="3930" />
                    <RANKING order="3" place="3" resultid="3139" />
                    <RANKING order="4" place="4" resultid="2107" />
                    <RANKING order="5" place="-1" resultid="2093" />
                    <RANKING order="6" place="-1" resultid="2305" />
                    <RANKING order="7" place="-1" resultid="5682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8131" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5288" />
                    <RANKING order="2" place="2" resultid="3262" />
                    <RANKING order="3" place="3" resultid="6505" />
                    <RANKING order="4" place="4" resultid="2842" />
                    <RANKING order="5" place="5" resultid="5867" />
                    <RANKING order="6" place="6" resultid="4162" />
                    <RANKING order="7" place="7" resultid="4658" />
                    <RANKING order="8" place="8" resultid="3152" />
                    <RANKING order="9" place="-1" resultid="2479" />
                    <RANKING order="10" place="-1" resultid="3218" />
                    <RANKING order="11" place="-1" resultid="5700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8132" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4392" />
                    <RANKING order="2" place="2" resultid="6003" />
                    <RANKING order="3" place="3" resultid="5733" />
                    <RANKING order="4" place="4" resultid="5750" />
                    <RANKING order="5" place="5" resultid="6120" />
                    <RANKING order="6" place="6" resultid="2416" />
                    <RANKING order="7" place="7" resultid="6104" />
                    <RANKING order="8" place="8" resultid="2887" />
                    <RANKING order="9" place="-1" resultid="2223" />
                    <RANKING order="10" place="-1" resultid="4622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8133" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5639" />
                    <RANKING order="2" place="2" resultid="4916" />
                    <RANKING order="3" place="3" resultid="5996" />
                    <RANKING order="4" place="4" resultid="5527" />
                    <RANKING order="5" place="5" resultid="2393" />
                    <RANKING order="6" place="6" resultid="4812" />
                    <RANKING order="7" place="7" resultid="6252" />
                    <RANKING order="8" place="8" resultid="2237" />
                    <RANKING order="9" place="9" resultid="4576" />
                    <RANKING order="10" place="-1" resultid="2006" />
                    <RANKING order="11" place="-1" resultid="2296" />
                    <RANKING order="12" place="-1" resultid="2468" />
                    <RANKING order="13" place="-1" resultid="5824" />
                    <RANKING order="14" place="-1" resultid="6491" />
                    <RANKING order="15" place="-1" resultid="4294" />
                    <RANKING order="16" place="-1" resultid="5756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8134" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6152" />
                    <RANKING order="2" place="2" resultid="4561" />
                    <RANKING order="3" place="3" resultid="3403" />
                    <RANKING order="4" place="4" resultid="4258" />
                    <RANKING order="5" place="5" resultid="6199" />
                    <RANKING order="6" place="6" resultid="3761" />
                    <RANKING order="7" place="7" resultid="3680" />
                    <RANKING order="8" place="8" resultid="6113" />
                    <RANKING order="9" place="9" resultid="5709" />
                    <RANKING order="10" place="10" resultid="3061" />
                    <RANKING order="11" place="-1" resultid="2253" />
                    <RANKING order="12" place="-1" resultid="4266" />
                    <RANKING order="13" place="-1" resultid="5080" />
                    <RANKING order="14" place="-1" resultid="5725" />
                    <RANKING order="15" place="-1" resultid="3999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8135" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2050" />
                    <RANKING order="2" place="2" resultid="6143" />
                    <RANKING order="3" place="3" resultid="4628" />
                    <RANKING order="4" place="4" resultid="5719" />
                    <RANKING order="5" place="5" resultid="6012" />
                    <RANKING order="6" place="6" resultid="3237" />
                    <RANKING order="7" place="7" resultid="5011" />
                    <RANKING order="8" place="8" resultid="4884" />
                    <RANKING order="9" place="9" resultid="4536" />
                    <RANKING order="10" place="-1" resultid="2113" />
                    <RANKING order="11" place="-1" resultid="5030" />
                    <RANKING order="12" place="-1" resultid="5101" />
                    <RANKING order="13" place="-1" resultid="4711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8136" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6021" />
                    <RANKING order="2" place="2" resultid="6028" />
                    <RANKING order="3" place="3" resultid="2547" />
                    <RANKING order="4" place="4" resultid="4181" />
                    <RANKING order="5" place="5" resultid="4509" />
                    <RANKING order="6" place="6" resultid="3551" />
                    <RANKING order="7" place="-1" resultid="3891" />
                    <RANKING order="8" place="-1" resultid="5790" />
                    <RANKING order="9" place="-1" resultid="4332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8137" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4402" />
                    <RANKING order="2" place="2" resultid="2860" />
                    <RANKING order="3" place="3" resultid="3502" />
                    <RANKING order="4" place="4" resultid="4680" />
                    <RANKING order="5" place="5" resultid="6437" />
                    <RANKING order="6" place="6" resultid="6369" />
                    <RANKING order="7" place="7" resultid="2587" />
                    <RANKING order="8" place="8" resultid="3269" />
                    <RANKING order="9" place="9" resultid="2851" />
                    <RANKING order="10" place="-1" resultid="2022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8138" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3733" />
                    <RANKING order="2" place="2" resultid="5152" />
                    <RANKING order="3" place="3" resultid="5852" />
                    <RANKING order="4" place="4" resultid="6260" />
                    <RANKING order="5" place="5" resultid="6057" />
                    <RANKING order="6" place="6" resultid="3513" />
                    <RANKING order="7" place="7" resultid="4481" />
                    <RANKING order="8" place="-1" resultid="2287" />
                    <RANKING order="9" place="-1" resultid="2521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8139" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2616" />
                    <RANKING order="2" place="2" resultid="3828" />
                    <RANKING order="3" place="3" resultid="2632" />
                    <RANKING order="4" place="4" resultid="4516" />
                    <RANKING order="5" place="-1" resultid="2324" />
                    <RANKING order="6" place="-1" resultid="5745" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7573" daytime="12:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7574" daytime="12:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7575" daytime="12:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7576" daytime="12:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7577" daytime="13:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7578" daytime="13:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7579" daytime="13:13" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7580" daytime="13:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7581" daytime="13:27" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7582" daytime="13:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7583" daytime="13:42" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7584" daytime="13:52" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1721" daytime="11:44" gender="F" number="41" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8110" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8111" agemax="89" agemin="85" name="M">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8112" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8113" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="8114" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4128" />
                    <RANKING order="2" place="2" resultid="4740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8115" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5669" />
                    <RANKING order="2" place="2" resultid="3287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8116" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3450" />
                    <RANKING order="2" place="2" resultid="2314" />
                    <RANKING order="3" place="3" resultid="5297" />
                    <RANKING order="4" place="4" resultid="3914" />
                    <RANKING order="5" place="5" resultid="2269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8117" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5675" />
                    <RANKING order="2" place="2" resultid="5801" />
                    <RANKING order="3" place="3" resultid="4777" />
                    <RANKING order="4" place="4" resultid="4795" />
                    <RANKING order="5" place="-1" resultid="4063" />
                    <RANKING order="6" place="-1" resultid="4233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8118" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2558" />
                    <RANKING order="2" place="2" resultid="6246" />
                    <RANKING order="3" place="3" resultid="4273" />
                    <RANKING order="4" place="4" resultid="5958" />
                    <RANKING order="5" place="5" resultid="3409" />
                    <RANKING order="6" place="6" resultid="6207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8119" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3805" />
                    <RANKING order="2" place="2" resultid="4327" />
                    <RANKING order="3" place="3" resultid="5093" />
                    <RANKING order="4" place="4" resultid="6450" />
                    <RANKING order="5" place="5" resultid="3922" />
                    <RANKING order="6" place="6" resultid="5894" />
                    <RANKING order="7" place="-1" resultid="6399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8120" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2484" />
                    <RANKING order="2" place="2" resultid="5563" />
                    <RANKING order="3" place="3" resultid="6170" />
                    <RANKING order="4" place="4" resultid="4982" />
                    <RANKING order="5" place="5" resultid="4493" />
                    <RANKING order="6" place="-1" resultid="5740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8121" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3715" />
                    <RANKING order="2" place="2" resultid="4646" />
                    <RANKING order="3" place="3" resultid="4490" />
                    <RANKING order="4" place="4" resultid="2400" />
                    <RANKING order="5" place="-1" resultid="5607" />
                    <RANKING order="6" place="-1" resultid="5615" />
                    <RANKING order="7" place="-1" resultid="6358" />
                    <RANKING order="8" place="-1" resultid="6393" />
                    <RANKING order="9" place="-1" resultid="4030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8122" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4044" />
                    <RANKING order="2" place="2" resultid="2830" />
                    <RANKING order="3" place="3" resultid="5137" />
                    <RANKING order="4" place="4" resultid="5582" />
                    <RANKING order="5" place="5" resultid="6161" />
                    <RANKING order="6" place="6" resultid="4665" />
                    <RANKING order="7" place="7" resultid="5875" />
                    <RANKING order="8" place="8" resultid="4478" />
                    <RANKING order="9" place="-1" resultid="4543" />
                    <RANKING order="10" place="-1" resultid="3884" />
                    <RANKING order="11" place="-1" resultid="4343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8123" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2983" />
                    <RANKING order="2" place="2" resultid="6134" />
                    <RANKING order="3" place="3" resultid="2041" />
                    <RANKING order="4" place="4" resultid="5840" />
                    <RANKING order="5" place="5" resultid="2144" />
                    <RANKING order="6" place="6" resultid="4382" />
                    <RANKING order="7" place="-1" resultid="3299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8124" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5988" />
                    <RANKING order="2" place="2" resultid="4219" />
                    <RANKING order="3" place="3" resultid="2680" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7566" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7567" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7568" daytime="11:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7569" daytime="12:03" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7570" daytime="12:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7571" daytime="12:19" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7572" daytime="12:28" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1705" daytime="11:28" gender="X" number="40" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8140" agemax="-1" agemin="280" name="F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3817" />
                    <RANKING order="2" place="2" resultid="4134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8141" agemax="279" agemin="240" name="E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="5710" />
                    <RANKING order="3" place="3" resultid="4138" />
                    <RANKING order="4" place="-1" resultid="4183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8142" agemax="239" agemin="200" name="D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4851" />
                    <RANKING order="2" place="2" resultid="5161" />
                    <RANKING order="3" place="3" resultid="6274" />
                    <RANKING order="4" place="4" resultid="3315" />
                    <RANKING order="5" place="5" resultid="6060" />
                    <RANKING order="6" place="6" resultid="4755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8143" agemax="199" agemin="160" name="C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3313" />
                    <RANKING order="2" place="2" resultid="6273" />
                    <RANKING order="3" place="3" resultid="2833" />
                    <RANKING order="4" place="4" resultid="3698" />
                    <RANKING order="5" place="5" resultid="4545" />
                    <RANKING order="6" place="6" resultid="6879" />
                    <RANKING order="7" place="7" resultid="5659" />
                    <RANKING order="8" place="8" resultid="4032" />
                    <RANKING order="9" place="9" resultid="5160" />
                    <RANKING order="10" place="-1" resultid="2328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8144" agemax="159" agemin="120" name="B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3036" />
                    <RANKING order="2" place="2" resultid="4753" />
                    <RANKING order="3" place="3" resultid="5278" />
                    <RANKING order="4" place="4" resultid="4754" />
                    <RANKING order="5" place="5" resultid="5060" />
                    <RANKING order="6" place="6" resultid="6878" />
                    <RANKING order="7" place="7" resultid="5071" />
                    <RANKING order="8" place="-1" resultid="5159" />
                    <RANKING order="9" place="-1" resultid="6478" />
                    <RANKING order="10" place="-1" resultid="3029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8145" agemax="119" agemin="100" name="A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6272" />
                    <RANKING order="2" place="2" resultid="3606" />
                    <RANKING order="3" place="-1" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8146" agemax="99" agemin="80" name="0" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3608" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7562" daytime="11:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7563" daytime="11:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7564" daytime="11:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7565" daytime="11:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1608" daytime="09:00" gender="F" number="34" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8020" agemax="94" agemin="90" name="N" />
                <AGEGROUP agegroupid="8021" agemax="89" agemin="85" name="M" />
                <AGEGROUP agegroupid="8022" agemax="84" agemin="80" name="L" />
                <AGEGROUP agegroupid="8023" agemax="79" agemin="75" name="K" />
                <AGEGROUP agegroupid="8024" agemax="74" agemin="70" name="J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8025" agemax="69" agemin="65" name="I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4087" />
                    <RANKING order="2" place="2" resultid="5668" />
                    <RANKING order="3" place="-1" resultid="3286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8026" agemax="64" agemin="60" name="H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3089" />
                    <RANKING order="2" place="2" resultid="4827" />
                    <RANKING order="3" place="3" resultid="4118" />
                    <RANKING order="4" place="4" resultid="4152" />
                    <RANKING order="5" place="-1" resultid="2313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8027" agemax="59" agemin="55" name="G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2796" />
                    <RANKING order="2" place="2" resultid="4776" />
                    <RANKING order="3" place="3" resultid="4794" />
                    <RANKING order="4" place="-1" resultid="3108" />
                    <RANKING order="5" place="-1" resultid="4079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8028" agemax="54" agemin="50" name="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2941" />
                    <RANKING order="2" place="2" resultid="2374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8029" agemax="49" agemin="45" name="E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3164" />
                    <RANKING order="2" place="2" resultid="6449" />
                    <RANKING order="3" place="3" resultid="4768" />
                    <RANKING order="4" place="4" resultid="6215" />
                    <RANKING order="5" place="5" resultid="6398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8030" agemax="44" agemin="40" name="D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3171" />
                    <RANKING order="2" place="2" resultid="4500" />
                    <RANKING order="3" place="3" resultid="5514" />
                    <RANKING order="4" place="4" resultid="3670" />
                    <RANKING order="5" place="-1" resultid="4904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8031" agemax="39" agemin="35" name="C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3384" />
                    <RANKING order="2" place="2" resultid="4940" />
                    <RANKING order="3" place="3" resultid="4956" />
                    <RANKING order="4" place="4" resultid="2818" />
                    <RANKING order="5" place="5" resultid="2867" />
                    <RANKING order="6" place="-1" resultid="5606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8032" agemax="34" agemin="30" name="B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6160" />
                    <RANKING order="2" place="2" resultid="3751" />
                    <RANKING order="3" place="3" resultid="2649" />
                    <RANKING order="4" place="4" resultid="6464" />
                    <RANKING order="5" place="5" resultid="5874" />
                    <RANKING order="6" place="-1" resultid="4664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8033" agemax="29" agemin="25" name="A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6133" />
                    <RANKING order="2" place="2" resultid="2787" />
                    <RANKING order="3" place="3" resultid="5498" />
                    <RANKING order="4" place="-1" resultid="2917" />
                    <RANKING order="5" place="-1" resultid="4467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8034" agemax="24" agemin="20" name="0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4197" />
                    <RANKING order="2" place="2" resultid="2624" />
                    <RANKING order="3" place="3" resultid="5969" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7507" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7508" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7509" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7510" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7511" daytime="09:11" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="3WADG" nation="POL" region="11" clubid="2930" name="3Waters  ASW Dąbrowa Grn.">
          <CONTACT email="borkowskasonia@interia.pl" name="Sonia Borkowska" phone="501273493" />
          <ATHLETES>
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="2931">
              <RESULTS>
                <RESULT eventid="1059" points="360" reactiontime="+75" swimtime="00:00:32.22" resultid="2932" heatid="7240" lane="3" entrytime="00:00:33.20" />
                <RESULT eventid="1272" points="305" reactiontime="+80" swimtime="00:01:14.65" resultid="2933" heatid="7344" lane="2" entrytime="00:01:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="2934" heatid="7410" lane="3" entrytime="00:01:42.00" />
                <RESULT eventid="1433" points="263" reactiontime="+73" swimtime="00:00:38.04" resultid="2935" heatid="7429" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1673" points="309" reactiontime="+69" swimtime="00:00:42.23" resultid="2936" heatid="7542" lane="7" entrytime="00:00:42.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-09-09" firstname="Anna" gender="F" lastname="Chmiel" nation="POL" athleteid="2946" />
            <ATHLETE birthdate="1966-03-15" firstname="Krystyna" gender="F" lastname="Noskiewicz - Czarnecka" nation="POL" athleteid="2937">
              <RESULTS>
                <RESULT eventid="1092" points="300" reactiontime="+95" swimtime="00:03:01.86" resultid="2938" heatid="7272" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:29.53" />
                    <SPLIT distance="150" swimtime="00:02:21.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="312" reactiontime="+85" swimtime="00:01:23.25" resultid="2939" heatid="7374" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="323" reactiontime="+74" swimtime="00:00:35.53" resultid="2940" heatid="7431" lane="3" entrytime="00:00:35.20" />
                <RESULT eventid="1608" points="249" reactiontime="+79" swimtime="00:01:26.71" resultid="2941" heatid="7509" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-20" firstname="Agnieszka" gender="F" lastname="Więk-Bernat" nation="POL" athleteid="2942">
              <RESULTS>
                <RESULT eventid="1240" points="296" reactiontime="+99" swimtime="00:03:21.91" resultid="2943" heatid="7330" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="211" reactiontime="+99" swimtime="00:01:32.41" resultid="2944" heatid="7455" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="2945" heatid="7527" lane="1" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="323" reactiontime="+92" swimtime="00:02:16.83" resultid="2947" heatid="7490" lane="6" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:06.82" />
                    <SPLIT distance="150" swimtime="00:01:44.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2946" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="2931" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2942" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="2937" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="293" reactiontime="+89" swimtime="00:02:34.05" resultid="2948" heatid="7400" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:01:57.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2942" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2931" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2937" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2946" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4MTZO" nation="POL" region="11" clubid="5847" name="4 Masters Team Żory">
          <ATHLETES>
            <ATHLETE birthdate="1993-04-01" firstname="Adrian" gender="M" lastname="Majdziński" nation="POL" athleteid="5846">
              <RESULTS>
                <RESULT eventid="1256" points="461" reactiontime="+76" swimtime="00:02:35.49" resultid="5848" heatid="7337" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="432" reactiontime="+78" swimtime="00:01:06.44" resultid="5849" heatid="7382" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="441" reactiontime="+74" swimtime="00:00:28.57" resultid="5850" heatid="7445" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1513" points="464" reactiontime="+76" swimtime="00:02:08.33" resultid="5851" heatid="7485" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:02.10" />
                    <SPLIT distance="150" swimtime="00:01:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="450" reactiontime="+74" swimtime="00:04:36.92" resultid="5852" heatid="7575" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:03.49" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:02:13.27" />
                    <SPLIT distance="250" swimtime="00:02:49.18" />
                    <SPLIT distance="300" swimtime="00:03:25.21" />
                    <SPLIT distance="350" swimtime="00:04:01.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5TWAR" nation="POL" region="14" clubid="4854" name="5 Styl Warszawa">
          <CONTACT name="Rodziewicz" />
          <ATHLETES>
            <ATHLETE birthdate="1977-01-01" firstname="Kamila" gender="F" lastname="Castoral" nation="POL" athleteid="4899">
              <RESULTS>
                <RESULT eventid="1240" points="176" reactiontime="+86" swimtime="00:03:59.78" resultid="4900" heatid="7329" lane="0" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                    <SPLIT distance="100" swimtime="00:01:53.86" />
                    <SPLIT distance="150" swimtime="00:02:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="48" swimtime="00:05:28.00" resultid="4901" heatid="7391" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.28" />
                    <SPLIT distance="100" swimtime="00:02:34.07" />
                    <SPLIT distance="150" swimtime="00:04:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="176" swimtime="00:01:51.25" resultid="4902" heatid="7409" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" status="DNF" swimtime="00:00:00.00" resultid="4903" heatid="8149" lane="5" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.25" />
                    <SPLIT distance="100" swimtime="00:02:32.42" />
                    <SPLIT distance="150" swimtime="00:03:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="4904" heatid="7508" lane="0" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-07" firstname="Marcin" gender="M" lastname="Cieślak" nation="POL" athleteid="4895">
              <RESULTS>
                <RESULT eventid="1288" points="807" reactiontime="+70" swimtime="00:00:48.26" resultid="4896" heatid="7367" lane="5" entrytime="00:00:47.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="792" reactiontime="+65" swimtime="00:00:23.50" resultid="4897" heatid="7451" lane="4" entrytime="00:00:22.80" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="4898" heatid="7522" lane="4" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-02" firstname="Tomasz" gender="M" lastname="Iwańczyk" nation="POL" athleteid="4885">
              <RESULTS>
                <RESULT eventid="1076" points="262" reactiontime="+86" swimtime="00:00:31.64" resultid="4886" heatid="7253" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1288" points="258" reactiontime="+92" swimtime="00:01:10.56" resultid="4887" heatid="7356" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="330" reactiontime="+75" swimtime="00:01:20.45" resultid="4888" heatid="7421" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4889" heatid="7552" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-09" firstname="Paweł" gender="M" lastname="Korzeniowski" nation="POL" athleteid="4890">
              <RESULTS>
                <RESULT eventid="1288" points="786" reactiontime="+69" swimtime="00:00:48.69" resultid="4891" heatid="7367" lane="4" entrytime="00:00:47.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="4892" heatid="7390" lane="4" entrytime="00:00:54.20" />
                <RESULT eventid="1449" points="780" reactiontime="+73" swimtime="00:00:23.62" resultid="4893" heatid="7451" lane="5" entrytime="00:00:23.50" />
                <RESULT eventid="1513" status="WDR" swimtime="00:00:00.00" resultid="4894" heatid="7488" lane="4" entrytime="00:01:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-16" firstname="Adrian" gender="M" lastname="Kulisz" nation="POL" athleteid="4880">
              <RESULTS>
                <RESULT eventid="1076" points="302" reactiontime="+95" swimtime="00:00:30.19" resultid="4881" heatid="7255" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1288" points="300" reactiontime="+81" swimtime="00:01:07.09" resultid="4882" heatid="7356" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="291" reactiontime="+76" swimtime="00:02:29.86" resultid="4883" heatid="7480" lane="5" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:50.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="230" reactiontime="+84" swimtime="00:05:45.94" resultid="4884" heatid="7580" lane="4" entrytime="00:05:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:15.86" />
                    <SPLIT distance="200" swimtime="00:02:40.16" />
                    <SPLIT distance="300" swimtime="00:04:09.30" />
                    <SPLIT distance="350" swimtime="00:04:55.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="495" reactiontime="+69" swimtime="00:01:54.31" resultid="4905" heatid="7403" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                    <SPLIT distance="150" swimtime="00:01:24.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4895" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4885" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="4890" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="4880" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="472" reactiontime="+69" swimtime="00:01:44.99" resultid="4906" heatid="7493" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.24" />
                    <SPLIT distance="100" swimtime="00:00:44.26" />
                    <SPLIT distance="150" swimtime="00:01:15.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4895" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4890" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="4885" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4880" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AASRY" nation="POL" region="11" clubid="2681" name="Ak. Aktywn. Seniora Rydułtowy">
          <CONTACT name="MARIAN OTLIK" phone="692112775" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="2691">
              <RESULTS>
                <RESULT eventid="1076" points="55" swimtime="00:00:53.01" resultid="2692" heatid="7247" lane="4" entrytime="00:00:52.00" />
                <RESULT comment="zmana stylu" eventid="1108" status="DSQ" swimtime="00:05:14.62" resultid="2693" heatid="7277" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.41" />
                    <SPLIT distance="100" swimtime="00:02:31.37" />
                    <SPLIT distance="150" swimtime="00:03:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="55" swimtime="00:05:15.12" resultid="2694" heatid="7333" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.10" />
                    <SPLIT distance="100" swimtime="00:02:36.69" />
                    <SPLIT distance="150" swimtime="00:03:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="45" swimtime="00:02:20.65" resultid="2695" heatid="7377" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2696" heatid="7435" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="1577" points="43" swimtime="00:11:10.55" resultid="2697" heatid="8154" lane="9" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.20" />
                    <SPLIT distance="100" swimtime="00:03:04.39" />
                    <SPLIT distance="150" swimtime="00:04:27.03" />
                    <SPLIT distance="200" swimtime="00:05:50.58" />
                    <SPLIT distance="250" swimtime="00:07:16.11" />
                    <SPLIT distance="300" swimtime="00:08:37.99" />
                    <SPLIT distance="350" swimtime="00:09:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="24" swimtime="00:02:45.00" resultid="2698" heatid="7513" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="70" swimtime="00:01:01.19" resultid="2699" heatid="7547" lane="3" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="2708">
              <RESULTS>
                <RESULT eventid="1108" points="155" reactiontime="+85" swimtime="00:03:23.99" resultid="2709" heatid="7279" lane="6" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                    <SPLIT distance="150" swimtime="00:02:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="181" reactiontime="+85" swimtime="00:24:58.61" resultid="2710" heatid="7304" lane="7" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:31.27" />
                    <SPLIT distance="150" swimtime="00:02:19.91" />
                    <SPLIT distance="200" swimtime="00:03:09.36" />
                    <SPLIT distance="250" swimtime="00:03:59.07" />
                    <SPLIT distance="300" swimtime="00:04:49.39" />
                    <SPLIT distance="350" swimtime="00:05:39.76" />
                    <SPLIT distance="400" swimtime="00:06:29.53" />
                    <SPLIT distance="450" swimtime="00:07:20.22" />
                    <SPLIT distance="500" swimtime="00:08:10.83" />
                    <SPLIT distance="550" swimtime="00:09:01.62" />
                    <SPLIT distance="600" swimtime="00:09:52.40" />
                    <SPLIT distance="650" swimtime="00:10:42.84" />
                    <SPLIT distance="700" swimtime="00:11:33.54" />
                    <SPLIT distance="750" swimtime="00:12:24.39" />
                    <SPLIT distance="800" swimtime="00:13:15.21" />
                    <SPLIT distance="850" swimtime="00:14:06.02" />
                    <SPLIT distance="900" swimtime="00:14:57.05" />
                    <SPLIT distance="950" swimtime="00:15:47.37" />
                    <SPLIT distance="1000" swimtime="00:16:38.45" />
                    <SPLIT distance="1050" swimtime="00:17:29.20" />
                    <SPLIT distance="1100" swimtime="00:18:19.72" />
                    <SPLIT distance="1150" swimtime="00:19:10.29" />
                    <SPLIT distance="1200" swimtime="00:20:00.86" />
                    <SPLIT distance="1250" swimtime="00:20:51.76" />
                    <SPLIT distance="1300" swimtime="00:21:42.18" />
                    <SPLIT distance="1350" swimtime="00:22:32.96" />
                    <SPLIT distance="1400" swimtime="00:23:23.47" />
                    <SPLIT distance="1450" swimtime="00:24:11.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="154" reactiontime="+82" swimtime="00:00:41.41" resultid="2711" heatid="7320" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1352" points="92" reactiontime="+92" swimtime="00:03:59.68" resultid="2712" heatid="7395" lane="2" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                    <SPLIT distance="100" swimtime="00:01:53.35" />
                    <SPLIT distance="150" swimtime="00:02:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="152" reactiontime="+97" swimtime="00:01:31.40" resultid="2713" heatid="7462" lane="6" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="137" reactiontime="+73" swimtime="00:07:35.79" resultid="2714" heatid="8155" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                    <SPLIT distance="100" swimtime="00:01:52.45" />
                    <SPLIT distance="150" swimtime="00:02:49.58" />
                    <SPLIT distance="200" swimtime="00:03:46.46" />
                    <SPLIT distance="250" swimtime="00:04:53.88" />
                    <SPLIT distance="300" swimtime="00:05:58.87" />
                    <SPLIT distance="350" swimtime="00:06:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="122" reactiontime="+79" swimtime="00:01:36.88" resultid="2715" heatid="7515" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="136" reactiontime="+79" swimtime="00:03:25.04" resultid="2716" heatid="7531" lane="5" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="2717">
              <RESULTS>
                <RESULT eventid="1076" points="304" reactiontime="+67" swimtime="00:00:30.12" resultid="2718" heatid="7252" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1108" points="205" reactiontime="+81" swimtime="00:03:05.69" resultid="2719" heatid="7279" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:29.73" />
                    <SPLIT distance="150" swimtime="00:02:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="259" reactiontime="+70" swimtime="00:01:10.47" resultid="2720" heatid="7354" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="198" reactiontime="+76" swimtime="00:01:26.10" resultid="2721" heatid="7379" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="225" reactiontime="+71" swimtime="00:00:35.75" resultid="2722" heatid="7439" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1577" points="160" reactiontime="+77" swimtime="00:07:13.38" resultid="2723" heatid="8155" lane="7" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:34.30" />
                    <SPLIT distance="150" swimtime="00:02:35.88" />
                    <SPLIT distance="200" swimtime="00:03:38.35" />
                    <SPLIT distance="250" swimtime="00:04:36.92" />
                    <SPLIT distance="300" swimtime="00:05:39.94" />
                    <SPLIT distance="350" swimtime="00:06:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="149" swimtime="00:01:30.52" resultid="2724" heatid="7514" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="175" reactiontime="+72" swimtime="00:00:45.11" resultid="2725" heatid="7548" lane="6" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="2682">
              <RESULTS>
                <RESULT eventid="1076" points="59" reactiontime="+95" swimtime="00:00:51.76" resultid="2683" heatid="7248" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1108" points="53" swimtime="00:04:50.49" resultid="2684" heatid="7277" lane="2" entrytime="00:04:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.85" />
                    <SPLIT distance="100" swimtime="00:02:16.37" />
                    <SPLIT distance="150" swimtime="00:03:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="53" swimtime="00:05:18.95" resultid="2685" heatid="7332" lane="5" entrytime="00:05:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.12" />
                    <SPLIT distance="100" swimtime="00:02:26.63" />
                    <SPLIT distance="150" swimtime="00:03:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="52" swimtime="00:02:13.86" resultid="2686" heatid="7377" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="58" reactiontime="+44" swimtime="00:02:23.27" resultid="2687" heatid="7415" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="32" swimtime="00:01:07.95" resultid="2688" heatid="7436" lane="2" entrytime="00:01:07.00" />
                <RESULT eventid="1657" points="44" reactiontime="+97" swimtime="00:04:57.74" resultid="2689" heatid="7530" lane="0" entrytime="00:04:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.63" />
                    <SPLIT distance="100" swimtime="00:02:22.64" />
                    <SPLIT distance="150" swimtime="00:03:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="63" reactiontime="+93" swimtime="00:01:03.24" resultid="2690" heatid="7547" lane="8" entrytime="00:01:01.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="2700">
              <RESULTS>
                <RESULT eventid="1076" points="20" swimtime="00:01:14.51" resultid="2701" heatid="7247" lane="7" />
                <RESULT eventid="1224" points="14" swimtime="00:01:31.66" resultid="2702" heatid="7316" lane="1" />
                <RESULT eventid="1288" points="20" reactiontime="+98" swimtime="00:02:44.56" resultid="2703" heatid="7350" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="14" swimtime="00:03:21.17" resultid="2704" heatid="7459" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="22" reactiontime="+85" swimtime="00:05:52.85" resultid="2705" heatid="7475" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.04" />
                    <SPLIT distance="100" swimtime="00:02:44.15" />
                    <SPLIT distance="150" swimtime="00:04:18.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="15" reactiontime="+93" swimtime="00:07:04.03" resultid="2706" heatid="7529" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.83" />
                    <SPLIT distance="100" swimtime="00:03:26.43" />
                    <SPLIT distance="150" swimtime="00:05:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="10" swimtime="00:01:56.95" resultid="2707" heatid="7546" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AFSSL" nation="POL" region="01" clubid="5854" name="Aqua Fit Środa Śl.">
          <ATHLETES>
            <ATHLETE birthdate="1985-07-05" firstname="Sebastian" gender="M" lastname="Figarski" nation="POL" athleteid="5853">
              <RESULTS>
                <RESULT eventid="1156" points="458" reactiontime="+95" swimtime="00:09:35.05" resultid="5855" heatid="7294" lane="9" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:42.00" />
                    <SPLIT distance="200" swimtime="00:02:17.72" />
                    <SPLIT distance="250" swimtime="00:02:53.77" />
                    <SPLIT distance="300" swimtime="00:03:30.65" />
                    <SPLIT distance="350" swimtime="00:04:07.83" />
                    <SPLIT distance="400" swimtime="00:04:44.89" />
                    <SPLIT distance="450" swimtime="00:05:21.62" />
                    <SPLIT distance="500" swimtime="00:05:58.19" />
                    <SPLIT distance="550" swimtime="00:06:34.87" />
                    <SPLIT distance="600" swimtime="00:07:11.46" />
                    <SPLIT distance="650" swimtime="00:07:48.20" />
                    <SPLIT distance="700" swimtime="00:08:24.85" />
                    <SPLIT distance="750" swimtime="00:09:00.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="418" reactiontime="+69" swimtime="00:00:29.71" resultid="5857" heatid="7325" lane="9" entrytime="00:00:31.20" />
                <RESULT eventid="1481" points="471" reactiontime="+72" swimtime="00:01:02.81" resultid="5858" heatid="7467" lane="9" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="424" reactiontime="+70" swimtime="00:02:20.57" resultid="5859" heatid="7536" lane="8" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQOLS" nation="POL" region="13" clubid="6088" name="Aquasfera Masters Olsztyn">
          <CONTACT name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="6162">
              <RESULTS>
                <RESULT eventid="1059" points="313" reactiontime="+81" swimtime="00:00:33.75" resultid="6163" heatid="7239" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1140" points="211" reactiontime="+86" swimtime="00:13:24.11" resultid="6164" heatid="7292" lane="3" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:15.66" />
                    <SPLIT distance="200" swimtime="00:03:08.38" />
                    <SPLIT distance="250" swimtime="00:04:03.56" />
                    <SPLIT distance="300" swimtime="00:04:53.77" />
                    <SPLIT distance="350" swimtime="00:05:45.24" />
                    <SPLIT distance="500" swimtime="00:08:21.30" />
                    <SPLIT distance="600" swimtime="00:10:04.95" />
                    <SPLIT distance="650" swimtime="00:10:56.04" />
                    <SPLIT distance="700" swimtime="00:11:47.05" />
                    <SPLIT distance="750" swimtime="00:12:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="338" reactiontime="+80" swimtime="00:00:36.85" resultid="6165" heatid="7311" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="6166" heatid="7368" lane="2" />
                <RESULT eventid="1465" points="276" reactiontime="+78" swimtime="00:01:24.48" resultid="6167" heatid="7456" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="6168" heatid="7468" lane="0" />
                <RESULT eventid="1641" points="199" reactiontime="+94" swimtime="00:03:24.03" resultid="6169" heatid="7524" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.95" />
                    <SPLIT distance="150" swimtime="00:02:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="215" reactiontime="+79" swimtime="00:06:30.06" resultid="6170" heatid="7569" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:01:31.37" />
                    <SPLIT distance="150" swimtime="00:02:19.92" />
                    <SPLIT distance="250" swimtime="00:04:00.86" />
                    <SPLIT distance="300" swimtime="00:04:51.53" />
                    <SPLIT distance="350" swimtime="00:05:41.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-14" firstname="Paweł" gender="M" lastname="Dąbrowski" nation="POL" athleteid="6191">
              <RESULTS>
                <RESULT eventid="1076" points="330" reactiontime="+78" swimtime="00:00:29.30" resultid="6192" heatid="7258" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1156" points="273" reactiontime="+86" swimtime="00:11:23.11" resultid="6193" heatid="7296" lane="7" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                    <SPLIT distance="200" swimtime="00:02:39.43" />
                    <SPLIT distance="250" swimtime="00:03:21.67" />
                    <SPLIT distance="300" swimtime="00:04:04.31" />
                    <SPLIT distance="350" swimtime="00:04:47.50" />
                    <SPLIT distance="400" swimtime="00:05:30.98" />
                    <SPLIT distance="450" swimtime="00:06:14.33" />
                    <SPLIT distance="500" swimtime="00:06:57.92" />
                    <SPLIT distance="550" swimtime="00:07:42.19" />
                    <SPLIT distance="600" swimtime="00:08:26.21" />
                    <SPLIT distance="650" swimtime="00:09:10.68" />
                    <SPLIT distance="700" swimtime="00:09:55.18" />
                    <SPLIT distance="750" swimtime="00:10:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="258" reactiontime="+73" swimtime="00:00:34.89" resultid="6194" heatid="7322" lane="9" entrytime="00:00:35.50" />
                <RESULT eventid="1288" points="327" reactiontime="+79" swimtime="00:01:05.21" resultid="6195" heatid="7357" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="263" reactiontime="+74" swimtime="00:01:16.29" resultid="6196" heatid="7459" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="312" reactiontime="+85" swimtime="00:02:26.36" resultid="6197" heatid="7481" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="244" reactiontime="+83" swimtime="00:02:48.92" resultid="6198" heatid="7533" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:06.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="290" reactiontime="+75" swimtime="00:05:20.44" resultid="6199" heatid="7578" lane="3" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:55.16" />
                    <SPLIT distance="200" swimtime="00:02:36.28" />
                    <SPLIT distance="250" swimtime="00:03:17.53" />
                    <SPLIT distance="300" swimtime="00:03:59.38" />
                    <SPLIT distance="350" swimtime="00:04:41.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="6238">
              <RESULTS>
                <RESULT eventid="1092" points="232" reactiontime="+92" swimtime="00:03:18.16" resultid="6239" heatid="7272" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:37.56" />
                    <SPLIT distance="150" swimtime="00:02:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="292" reactiontime="+93" swimtime="00:23:04.82" resultid="6240" heatid="7300" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:10.36" />
                    <SPLIT distance="200" swimtime="00:02:55.90" />
                    <SPLIT distance="250" swimtime="00:03:41.89" />
                    <SPLIT distance="300" swimtime="00:04:28.21" />
                    <SPLIT distance="350" swimtime="00:05:14.87" />
                    <SPLIT distance="400" swimtime="00:06:01.34" />
                    <SPLIT distance="450" swimtime="00:06:47.84" />
                    <SPLIT distance="500" swimtime="00:07:34.25" />
                    <SPLIT distance="550" swimtime="00:08:20.87" />
                    <SPLIT distance="600" swimtime="00:09:07.13" />
                    <SPLIT distance="650" swimtime="00:09:53.70" />
                    <SPLIT distance="700" swimtime="00:10:40.31" />
                    <SPLIT distance="750" swimtime="00:11:26.52" />
                    <SPLIT distance="800" swimtime="00:12:13.11" />
                    <SPLIT distance="850" swimtime="00:12:59.75" />
                    <SPLIT distance="900" swimtime="00:13:46.11" />
                    <SPLIT distance="950" swimtime="00:14:32.99" />
                    <SPLIT distance="1000" swimtime="00:15:19.55" />
                    <SPLIT distance="1050" swimtime="00:16:06.69" />
                    <SPLIT distance="1100" swimtime="00:16:53.08" />
                    <SPLIT distance="1150" swimtime="00:17:39.75" />
                    <SPLIT distance="1200" swimtime="00:18:26.01" />
                    <SPLIT distance="1250" swimtime="00:19:12.43" />
                    <SPLIT distance="1300" swimtime="00:19:59.08" />
                    <SPLIT distance="1350" swimtime="00:20:45.79" />
                    <SPLIT distance="1400" swimtime="00:21:32.41" />
                    <SPLIT distance="1450" swimtime="00:22:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="221" reactiontime="+93" swimtime="00:03:42.43" resultid="6241" heatid="7330" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                    <SPLIT distance="100" swimtime="00:01:48.57" />
                    <SPLIT distance="150" swimtime="00:02:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="278" reactiontime="+89" swimtime="00:01:16.98" resultid="6242" heatid="7343" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="295" reactiontime="+91" swimtime="00:02:45.79" resultid="6243" heatid="7469" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:21.72" />
                    <SPLIT distance="150" swimtime="00:02:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="232" reactiontime="+98" swimtime="00:07:01.14" resultid="6244" heatid="8150" lane="6" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.93" />
                    <SPLIT distance="100" swimtime="00:01:51.57" />
                    <SPLIT distance="150" swimtime="00:02:45.21" />
                    <SPLIT distance="200" swimtime="00:03:37.93" />
                    <SPLIT distance="250" swimtime="00:04:35.36" />
                    <SPLIT distance="300" swimtime="00:05:31.81" />
                    <SPLIT distance="350" swimtime="00:06:17.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="202" reactiontime="+97" swimtime="00:03:23.00" resultid="6245" heatid="7525" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:41.05" />
                    <SPLIT distance="150" swimtime="00:02:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="285" reactiontime="+90" swimtime="00:05:55.45" resultid="6246" heatid="7568" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="150" swimtime="00:02:10.59" />
                    <SPLIT distance="200" swimtime="00:02:56.36" />
                    <SPLIT distance="250" swimtime="00:03:41.59" />
                    <SPLIT distance="300" swimtime="00:04:26.72" />
                    <SPLIT distance="350" swimtime="00:05:12.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-10-02" firstname="Grzegorz" gender="M" lastname="Grabowski" nation="POL" athleteid="6232">
              <RESULTS>
                <RESULT eventid="1076" points="437" reactiontime="+74" swimtime="00:00:26.69" resultid="6233" heatid="7264" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1224" points="256" reactiontime="+66" swimtime="00:00:34.99" resultid="6234" heatid="7323" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1288" points="415" reactiontime="+64" swimtime="00:01:00.24" resultid="6235" heatid="7356" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="370" reactiontime="+70" swimtime="00:00:30.27" resultid="6236" heatid="7444" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="6237" heatid="7558" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="6144">
              <RESULTS>
                <RESULT eventid="1076" points="493" reactiontime="+69" swimtime="00:00:25.63" resultid="6145" heatid="7263" lane="4" entrytime="00:00:27.20" />
                <RESULT comment="Rekord Polski Masters kategoria E" eventid="1188" points="486" reactiontime="+79" swimtime="00:17:57.93" resultid="6146" heatid="7302" lane="6" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:44.52" />
                    <SPLIT distance="200" swimtime="00:02:20.63" />
                    <SPLIT distance="250" swimtime="00:02:56.78" />
                    <SPLIT distance="300" swimtime="00:03:32.85" />
                    <SPLIT distance="350" swimtime="00:04:08.98" />
                    <SPLIT distance="400" swimtime="00:04:45.55" />
                    <SPLIT distance="450" swimtime="00:05:21.82" />
                    <SPLIT distance="500" swimtime="00:05:57.98" />
                    <SPLIT distance="550" swimtime="00:06:34.09" />
                    <SPLIT distance="600" swimtime="00:07:10.01" />
                    <SPLIT distance="650" swimtime="00:07:46.45" />
                    <SPLIT distance="700" swimtime="00:08:23.00" />
                    <SPLIT distance="750" swimtime="00:08:59.14" />
                    <SPLIT distance="800" swimtime="00:09:35.67" />
                    <SPLIT distance="850" swimtime="00:10:11.96" />
                    <SPLIT distance="900" swimtime="00:10:48.20" />
                    <SPLIT distance="950" swimtime="00:11:24.23" />
                    <SPLIT distance="1000" swimtime="00:12:00.24" />
                    <SPLIT distance="1050" swimtime="00:12:36.35" />
                    <SPLIT distance="1100" swimtime="00:13:12.12" />
                    <SPLIT distance="1150" swimtime="00:13:48.08" />
                    <SPLIT distance="1200" swimtime="00:14:24.17" />
                    <SPLIT distance="1250" swimtime="00:15:00.13" />
                    <SPLIT distance="1300" swimtime="00:15:36.09" />
                    <SPLIT distance="1350" swimtime="00:16:12.37" />
                    <SPLIT distance="1400" swimtime="00:16:48.42" />
                    <SPLIT distance="1450" swimtime="00:17:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="499" reactiontime="+72" swimtime="00:00:56.65" resultid="6147" heatid="7365" lane="2" entrytime="00:00:57.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="422" reactiontime="+79" swimtime="00:02:24.22" resultid="6148" heatid="7397" lane="2" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="150" swimtime="00:01:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="522" reactiontime="+72" swimtime="00:02:03.40" resultid="6149" heatid="7487" lane="3" entrytime="00:02:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:00:59.91" />
                    <SPLIT distance="150" swimtime="00:01:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="442" reactiontime="+74" swimtime="00:05:09.01" resultid="6150" heatid="8158" lane="7" entrytime="00:05:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                    <SPLIT distance="200" swimtime="00:02:33.21" />
                    <SPLIT distance="250" swimtime="00:03:17.32" />
                    <SPLIT distance="300" swimtime="00:04:01.16" />
                    <SPLIT distance="350" swimtime="00:04:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="461" reactiontime="+70" swimtime="00:01:02.20" resultid="6151" heatid="7520" lane="9" entrytime="00:01:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria E" eventid="1737" points="498" reactiontime="+74" swimtime="00:04:27.64" resultid="6152" heatid="7573" lane="2" entrytime="00:04:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:04.00" />
                    <SPLIT distance="150" swimtime="00:01:38.06" />
                    <SPLIT distance="200" swimtime="00:02:12.52" />
                    <SPLIT distance="250" swimtime="00:02:47.31" />
                    <SPLIT distance="300" swimtime="00:03:21.81" />
                    <SPLIT distance="350" swimtime="00:03:55.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="6217">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="6218" heatid="7281" lane="5" entrytime="00:02:45.00" />
                <RESULT eventid="1256" points="298" reactiontime="+79" swimtime="00:02:59.74" resultid="6219" heatid="7338" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="283" reactiontime="+78" swimtime="00:02:44.85" resultid="6220" heatid="7397" lane="5" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:57.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="325" reactiontime="+77" swimtime="00:01:20.86" resultid="6221" heatid="7423" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="6222" heatid="8157" lane="7" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="6135">
              <RESULTS>
                <RESULT eventid="1076" points="438" reactiontime="+63" swimtime="00:00:26.67" resultid="6136" heatid="7262" lane="5" entrytime="00:00:27.80" />
                <RESULT eventid="1188" points="426" reactiontime="+68" swimtime="00:18:46.49" resultid="6137" heatid="7302" lane="5" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:47.39" />
                    <SPLIT distance="200" swimtime="00:02:24.81" />
                    <SPLIT distance="250" swimtime="00:03:02.46" />
                    <SPLIT distance="300" swimtime="00:03:40.15" />
                    <SPLIT distance="350" swimtime="00:04:17.88" />
                    <SPLIT distance="400" swimtime="00:04:56.07" />
                    <SPLIT distance="450" swimtime="00:05:34.38" />
                    <SPLIT distance="500" swimtime="00:06:12.33" />
                    <SPLIT distance="550" swimtime="00:06:50.34" />
                    <SPLIT distance="600" swimtime="00:07:28.10" />
                    <SPLIT distance="650" swimtime="00:08:06.11" />
                    <SPLIT distance="700" swimtime="00:08:44.20" />
                    <SPLIT distance="750" swimtime="00:09:21.96" />
                    <SPLIT distance="800" swimtime="00:09:59.93" />
                    <SPLIT distance="850" swimtime="00:10:37.59" />
                    <SPLIT distance="900" swimtime="00:11:15.39" />
                    <SPLIT distance="950" swimtime="00:11:53.19" />
                    <SPLIT distance="1000" swimtime="00:12:31.21" />
                    <SPLIT distance="1050" swimtime="00:13:08.96" />
                    <SPLIT distance="1100" swimtime="00:13:46.79" />
                    <SPLIT distance="1150" swimtime="00:14:24.75" />
                    <SPLIT distance="1200" swimtime="00:15:02.30" />
                    <SPLIT distance="1250" swimtime="00:15:40.01" />
                    <SPLIT distance="1300" swimtime="00:16:17.73" />
                    <SPLIT distance="1350" swimtime="00:16:55.88" />
                    <SPLIT distance="1400" swimtime="00:17:33.82" />
                    <SPLIT distance="1450" swimtime="00:18:11.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="337" reactiontime="+66" swimtime="00:00:31.92" resultid="6138" heatid="7324" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1288" points="422" reactiontime="+64" swimtime="00:00:59.87" resultid="6139" heatid="7362" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="425" reactiontime="+64" swimtime="00:02:12.09" resultid="6140" heatid="7485" lane="5" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:03.52" />
                    <SPLIT distance="150" swimtime="00:01:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="359" reactiontime="+63" swimtime="00:05:31.25" resultid="6141" heatid="8158" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:02.68" />
                    <SPLIT distance="200" swimtime="00:02:45.62" />
                    <SPLIT distance="250" swimtime="00:03:33.28" />
                    <SPLIT distance="300" swimtime="00:04:20.62" />
                    <SPLIT distance="350" swimtime="00:04:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="307" reactiontime="+63" swimtime="00:02:36.45" resultid="6142" heatid="7534" lane="8" entrytime="00:02:41.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                    <SPLIT distance="150" swimtime="00:01:57.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="429" reactiontime="+65" swimtime="00:04:41.40" resultid="6143" heatid="7575" lane="4" entrytime="00:04:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:43.21" />
                    <SPLIT distance="200" swimtime="00:02:19.24" />
                    <SPLIT distance="250" swimtime="00:02:55.34" />
                    <SPLIT distance="300" swimtime="00:03:32.06" />
                    <SPLIT distance="350" swimtime="00:04:08.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-14" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="6089">
              <RESULTS>
                <RESULT eventid="1076" points="442" reactiontime="+74" swimtime="00:00:26.59" resultid="6090" heatid="7263" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1108" points="399" reactiontime="+73" swimtime="00:02:28.90" resultid="6091" heatid="7283" lane="2" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="434" reactiontime="+67" swimtime="00:02:38.65" resultid="6092" heatid="7338" lane="4" entrytime="00:02:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="397" reactiontime="+68" swimtime="00:01:08.37" resultid="6093" heatid="7386" lane="0" entrytime="00:01:11.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="460" reactiontime="+56" swimtime="00:01:12.00" resultid="6094" heatid="7423" lane="4" entrytime="00:01:17.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="364" reactiontime="+72" swimtime="00:02:19.08" resultid="6095" heatid="7481" lane="0" entrytime="00:02:35.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:45.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="468" reactiontime="+63" swimtime="00:00:32.52" resultid="6096" heatid="7557" lane="6" entrytime="00:00:35.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="6097">
              <RESULTS>
                <RESULT eventid="1156" points="242" reactiontime="+99" swimtime="00:11:51.29" resultid="6098" heatid="7297" lane="2" entrytime="00:12:06.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:22.58" />
                    <SPLIT distance="150" swimtime="00:02:08.01" />
                    <SPLIT distance="200" swimtime="00:02:52.61" />
                    <SPLIT distance="250" swimtime="00:03:37.41" />
                    <SPLIT distance="300" swimtime="00:04:22.43" />
                    <SPLIT distance="350" swimtime="00:05:07.33" />
                    <SPLIT distance="400" swimtime="00:05:52.59" />
                    <SPLIT distance="450" swimtime="00:06:38.19" />
                    <SPLIT distance="500" swimtime="00:07:23.22" />
                    <SPLIT distance="550" swimtime="00:08:09.09" />
                    <SPLIT distance="600" swimtime="00:08:54.98" />
                    <SPLIT distance="650" swimtime="00:09:40.74" />
                    <SPLIT distance="700" swimtime="00:10:25.74" />
                    <SPLIT distance="750" swimtime="00:11:10.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="235" reactiontime="+99" swimtime="00:03:14.70" resultid="6099" heatid="7335" lane="2" entrytime="00:03:24.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="100" swimtime="00:01:36.50" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="221" swimtime="00:01:23.05" resultid="6100" heatid="7381" lane="0" entrytime="00:01:25.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="225" swimtime="00:01:31.31" resultid="6101" heatid="7417" lane="6" entrytime="00:01:43.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="222" reactiontime="+99" swimtime="00:06:28.43" resultid="6102" heatid="8156" lane="9" entrytime="00:06:59.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:35.02" />
                    <SPLIT distance="150" swimtime="00:02:30.21" />
                    <SPLIT distance="200" swimtime="00:03:23.11" />
                    <SPLIT distance="250" swimtime="00:04:14.81" />
                    <SPLIT distance="300" swimtime="00:05:06.75" />
                    <SPLIT distance="350" swimtime="00:05:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="149" swimtime="00:01:30.50" resultid="6103" heatid="7515" lane="0" entrytime="00:01:34.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="221" reactiontime="+97" swimtime="00:05:50.61" resultid="6104" heatid="7580" lane="1" entrytime="00:06:01.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:07.29" />
                    <SPLIT distance="200" swimtime="00:02:51.65" />
                    <SPLIT distance="250" swimtime="00:03:36.09" />
                    <SPLIT distance="300" swimtime="00:04:20.13" />
                    <SPLIT distance="350" swimtime="00:05:03.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="6223">
              <RESULTS>
                <RESULT eventid="1059" points="362" reactiontime="+93" swimtime="00:00:32.17" resultid="6224" heatid="7241" lane="3" entrytime="00:00:32.10" />
                <RESULT eventid="1207" points="282" reactiontime="+79" swimtime="00:00:39.11" resultid="6226" heatid="7311" lane="9" entrytime="00:00:39.90" />
                <RESULT eventid="1272" points="342" reactiontime="+86" swimtime="00:01:11.83" resultid="6227" heatid="7345" lane="6" entrytime="00:01:12.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="292" reactiontime="+83" swimtime="00:00:36.74" resultid="6228" heatid="7431" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1641" points="258" reactiontime="+82" swimtime="00:03:07.16" resultid="6231" heatid="7526" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:30.21" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-19" firstname="Oriana" gender="F" lastname="Lewandowska" nation="POL" athleteid="6128">
              <RESULTS>
                <RESULT eventid="1140" points="607" reactiontime="+86" swimtime="00:09:25.86" resultid="6129" heatid="7290" lane="4" entrytime="00:09:40.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                    <SPLIT distance="200" swimtime="00:02:20.41" />
                    <SPLIT distance="250" swimtime="00:02:56.26" />
                    <SPLIT distance="300" swimtime="00:03:32.00" />
                    <SPLIT distance="350" swimtime="00:04:07.79" />
                    <SPLIT distance="400" swimtime="00:04:43.72" />
                    <SPLIT distance="450" swimtime="00:05:19.35" />
                    <SPLIT distance="500" swimtime="00:05:54.98" />
                    <SPLIT distance="550" swimtime="00:06:30.91" />
                    <SPLIT distance="600" swimtime="00:07:06.36" />
                    <SPLIT distance="650" swimtime="00:07:42.06" />
                    <SPLIT distance="700" swimtime="00:08:17.66" />
                    <SPLIT distance="750" swimtime="00:08:52.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="638" reactiontime="+89" swimtime="00:02:18.91" resultid="6130" heatid="7393" lane="4" entrytime="00:02:20.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="507" reactiontime="+87" swimtime="00:00:30.57" resultid="6131" heatid="7434" lane="0" entrytime="00:00:30.20" />
                <RESULT eventid="1497" points="565" reactiontime="+81" swimtime="00:02:13.56" resultid="6132" heatid="7474" lane="2" entrytime="00:02:15.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:05.75" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="567" reactiontime="+79" swimtime="00:01:05.95" resultid="6133" heatid="7511" lane="3" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="563" reactiontime="+84" swimtime="00:04:43.20" resultid="6134" heatid="7566" lane="3" entrytime="00:04:48.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:45.48" />
                    <SPLIT distance="200" swimtime="00:02:21.65" />
                    <SPLIT distance="250" swimtime="00:02:57.89" />
                    <SPLIT distance="300" swimtime="00:03:33.88" />
                    <SPLIT distance="350" swimtime="00:04:09.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="6105">
              <RESULTS>
                <RESULT eventid="1076" points="245" reactiontime="+87" swimtime="00:00:32.37" resultid="6106" heatid="7254" lane="7" entrytime="00:00:33.21" />
                <RESULT eventid="1156" points="284" reactiontime="+89" swimtime="00:11:14.24" resultid="6107" heatid="7296" lane="1" entrytime="00:11:24.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                    <SPLIT distance="200" swimtime="00:02:40.76" />
                    <SPLIT distance="250" swimtime="00:03:22.51" />
                    <SPLIT distance="300" swimtime="00:04:04.85" />
                    <SPLIT distance="350" swimtime="00:04:46.99" />
                    <SPLIT distance="400" swimtime="00:05:30.10" />
                    <SPLIT distance="450" swimtime="00:06:13.27" />
                    <SPLIT distance="500" swimtime="00:06:56.52" />
                    <SPLIT distance="550" swimtime="00:07:39.73" />
                    <SPLIT distance="600" swimtime="00:08:23.11" />
                    <SPLIT distance="650" swimtime="00:09:06.14" />
                    <SPLIT distance="700" swimtime="00:09:49.21" />
                    <SPLIT distance="750" swimtime="00:10:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="172" reactiontime="+68" swimtime="00:00:39.92" resultid="6108" heatid="7319" lane="5" entrytime="00:00:41.36" />
                <RESULT eventid="1288" points="249" reactiontime="+75" swimtime="00:01:11.38" resultid="6109" heatid="7355" lane="8" entrytime="00:01:13.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="186" reactiontime="+85" swimtime="00:00:38.05" resultid="6110" heatid="7439" lane="8" entrytime="00:00:38.05" />
                <RESULT eventid="1513" points="267" reactiontime="+84" swimtime="00:02:34.23" resultid="6111" heatid="7481" lane="8" entrytime="00:02:35.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="6112" heatid="7514" lane="5" entrytime="00:01:42.68" />
                <RESULT eventid="1737" points="274" reactiontime="+77" swimtime="00:05:26.59" resultid="6113" heatid="7578" lane="2" entrytime="00:05:28.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:57.07" />
                    <SPLIT distance="200" swimtime="00:02:38.32" />
                    <SPLIT distance="250" swimtime="00:03:20.14" />
                    <SPLIT distance="300" swimtime="00:04:02.43" />
                    <SPLIT distance="350" swimtime="00:04:44.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-18" firstname="Bogdan" gender="M" lastname="Milewski" nation="POL" athleteid="6121">
              <RESULTS>
                <RESULT eventid="1108" points="221" reactiontime="+82" swimtime="00:03:01.11" resultid="6122" heatid="7280" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="256" reactiontime="+89" swimtime="00:01:10.74" resultid="6123" heatid="7355" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="262" reactiontime="+80" swimtime="00:01:26.90" resultid="6124" heatid="7420" lane="9" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="244" reactiontime="+81" swimtime="00:00:34.80" resultid="6125" heatid="7440" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="1625" points="181" reactiontime="+82" swimtime="00:01:24.99" resultid="6126" heatid="7516" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="282" reactiontime="+81" swimtime="00:00:38.47" resultid="6127" heatid="7553" lane="1" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="6247">
              <RESULTS>
                <RESULT eventid="1156" points="252" swimtime="00:11:41.62" resultid="6248" heatid="7296" lane="0" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:20.66" />
                    <SPLIT distance="150" swimtime="00:02:03.94" />
                    <SPLIT distance="200" swimtime="00:02:47.43" />
                    <SPLIT distance="250" swimtime="00:03:31.56" />
                    <SPLIT distance="300" swimtime="00:04:16.07" />
                    <SPLIT distance="350" swimtime="00:05:00.70" />
                    <SPLIT distance="400" swimtime="00:05:45.17" />
                    <SPLIT distance="450" swimtime="00:06:29.72" />
                    <SPLIT distance="500" swimtime="00:07:14.80" />
                    <SPLIT distance="550" swimtime="00:07:59.54" />
                    <SPLIT distance="600" swimtime="00:08:44.27" />
                    <SPLIT distance="650" swimtime="00:09:29.34" />
                    <SPLIT distance="700" swimtime="00:10:14.03" />
                    <SPLIT distance="750" swimtime="00:10:58.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="215" reactiontime="+87" swimtime="00:03:00.54" resultid="6249" heatid="7396" lane="5" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="150" swimtime="00:02:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="223" reactiontime="+87" swimtime="00:06:27.83" resultid="6250" heatid="8156" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="150" swimtime="00:02:23.28" />
                    <SPLIT distance="200" swimtime="00:03:16.22" />
                    <SPLIT distance="250" swimtime="00:04:11.30" />
                    <SPLIT distance="300" swimtime="00:05:04.93" />
                    <SPLIT distance="350" swimtime="00:05:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="235" reactiontime="+83" swimtime="00:00:40.88" resultid="6251" heatid="7551" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1737" points="234" reactiontime="+86" swimtime="00:05:44.23" resultid="6252" heatid="7579" lane="7" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:21.64" />
                    <SPLIT distance="150" swimtime="00:02:05.12" />
                    <SPLIT distance="200" swimtime="00:02:49.30" />
                    <SPLIT distance="250" swimtime="00:03:33.52" />
                    <SPLIT distance="300" swimtime="00:04:18.00" />
                    <SPLIT distance="350" swimtime="00:05:02.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-15" firstname="Mieszko" gender="M" lastname="Palmi-Kukiełko" nation="POL" athleteid="6171">
              <RESULTS>
                <RESULT eventid="1108" points="600" reactiontime="+78" swimtime="00:02:09.93" resultid="6172" heatid="7285" lane="4" entrytime="00:02:09.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                    <SPLIT distance="100" swimtime="00:00:59.63" />
                    <SPLIT distance="150" swimtime="00:01:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="537" reactiontime="+73" swimtime="00:17:22.89" resultid="6173" heatid="7302" lane="4" entrytime="00:17:07.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:02.56" />
                    <SPLIT distance="150" swimtime="00:01:37.03" />
                    <SPLIT distance="200" swimtime="00:02:12.33" />
                    <SPLIT distance="250" swimtime="00:02:47.82" />
                    <SPLIT distance="300" swimtime="00:03:23.41" />
                    <SPLIT distance="350" swimtime="00:03:59.03" />
                    <SPLIT distance="400" swimtime="00:04:34.95" />
                    <SPLIT distance="450" swimtime="00:05:10.50" />
                    <SPLIT distance="500" swimtime="00:05:46.18" />
                    <SPLIT distance="550" swimtime="00:06:21.84" />
                    <SPLIT distance="600" swimtime="00:06:57.73" />
                    <SPLIT distance="650" swimtime="00:07:33.02" />
                    <SPLIT distance="700" swimtime="00:08:08.15" />
                    <SPLIT distance="750" swimtime="00:08:43.51" />
                    <SPLIT distance="800" swimtime="00:09:18.61" />
                    <SPLIT distance="850" swimtime="00:09:54.07" />
                    <SPLIT distance="900" swimtime="00:10:29.62" />
                    <SPLIT distance="950" swimtime="00:11:04.89" />
                    <SPLIT distance="1000" swimtime="00:11:39.95" />
                    <SPLIT distance="1050" swimtime="00:12:14.49" />
                    <SPLIT distance="1100" swimtime="00:12:48.80" />
                    <SPLIT distance="1150" swimtime="00:13:23.06" />
                    <SPLIT distance="1200" swimtime="00:13:57.61" />
                    <SPLIT distance="1250" swimtime="00:14:32.62" />
                    <SPLIT distance="1300" swimtime="00:15:07.15" />
                    <SPLIT distance="1350" swimtime="00:15:41.65" />
                    <SPLIT distance="1400" swimtime="00:16:15.96" />
                    <SPLIT distance="1450" swimtime="00:16:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="609" reactiontime="+75" swimtime="00:00:59.29" resultid="6174" heatid="7390" lane="6" entrytime="00:00:58.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="576" reactiontime="+76" swimtime="00:02:10.08" resultid="6175" heatid="7398" lane="3" entrytime="00:02:11.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="150" swimtime="00:01:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="603" reactiontime="+73" swimtime="00:01:57.59" resultid="6176" heatid="7488" lane="2" entrytime="00:01:58.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="150" swimtime="00:01:27.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="599" reactiontime="+74" swimtime="00:04:39.29" resultid="6177" heatid="8158" lane="4" entrytime="00:04:38.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="200" swimtime="00:02:16.73" />
                    <SPLIT distance="250" swimtime="00:02:56.13" />
                    <SPLIT distance="300" swimtime="00:03:35.91" />
                    <SPLIT distance="350" swimtime="00:04:08.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="600" reactiontime="+71" swimtime="00:00:56.99" resultid="6178" heatid="7522" lane="2" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="517" reactiontime="+73" swimtime="00:02:11.56" resultid="6179" heatid="7536" lane="4" entrytime="00:02:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:03.64" />
                    <SPLIT distance="150" swimtime="00:01:37.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-03-10" firstname="Kartarzyna" gender="F" lastname="Sienkiewicz" nation="POL" athleteid="6208">
              <RESULTS>
                <RESULT eventid="1092" points="205" reactiontime="+80" swimtime="00:03:26.39" resultid="6209" heatid="7272" lane="1" entrytime="00:03:35.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:01:40.21" />
                    <SPLIT distance="150" swimtime="00:02:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="170" reactiontime="+87" swimtime="00:14:24.10" resultid="6210" heatid="7292" lane="6" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:32.61" />
                    <SPLIT distance="150" swimtime="00:02:25.69" />
                    <SPLIT distance="200" swimtime="00:03:19.98" />
                    <SPLIT distance="250" swimtime="00:04:14.85" />
                    <SPLIT distance="300" swimtime="00:05:10.18" />
                    <SPLIT distance="350" swimtime="00:06:05.85" />
                    <SPLIT distance="400" swimtime="00:07:02.12" />
                    <SPLIT distance="450" swimtime="00:07:57.96" />
                    <SPLIT distance="500" swimtime="00:08:54.02" />
                    <SPLIT distance="550" swimtime="00:09:50.29" />
                    <SPLIT distance="600" swimtime="00:10:45.19" />
                    <SPLIT distance="650" swimtime="00:11:41.46" />
                    <SPLIT distance="700" swimtime="00:12:36.85" />
                    <SPLIT distance="750" swimtime="00:13:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="214" reactiontime="+91" swimtime="00:01:23.93" resultid="6211" heatid="7343" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="216" reactiontime="+90" swimtime="00:01:34.04" resultid="6212" heatid="7371" lane="1" entrytime="00:01:35.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="223" reactiontime="+84" swimtime="00:00:40.19" resultid="6213" heatid="7428" lane="6" entrytime="00:00:41.98" />
                <RESULT eventid="1497" points="191" reactiontime="+88" swimtime="00:03:11.53" resultid="6214" heatid="7470" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:02:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="159" reactiontime="+93" swimtime="00:01:40.60" resultid="6215" heatid="7507" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="6216" heatid="7539" lane="1" entrytime="00:00:51.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="6180">
              <RESULTS>
                <RESULT eventid="1156" points="300" reactiontime="+97" swimtime="00:11:01.95" resultid="6181" heatid="7296" lane="2" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                    <SPLIT distance="200" swimtime="00:02:33.31" />
                    <SPLIT distance="250" swimtime="00:03:14.89" />
                    <SPLIT distance="300" swimtime="00:03:56.85" />
                    <SPLIT distance="350" swimtime="00:04:38.91" />
                    <SPLIT distance="400" swimtime="00:05:22.10" />
                    <SPLIT distance="450" swimtime="00:06:04.80" />
                    <SPLIT distance="500" swimtime="00:06:47.19" />
                    <SPLIT distance="550" swimtime="00:07:30.51" />
                    <SPLIT distance="600" swimtime="00:08:13.65" />
                    <SPLIT distance="650" swimtime="00:08:56.71" />
                    <SPLIT distance="700" swimtime="00:09:39.95" />
                    <SPLIT distance="750" swimtime="00:10:22.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="357" reactiontime="+84" swimtime="00:01:03.31" resultid="6182" heatid="7357" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6183" heatid="7440" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1513" points="325" reactiontime="+82" swimtime="00:02:24.42" resultid="6184" heatid="7481" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:46.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-15" firstname="Adam" gender="M" lastname="Szmit" nation="POL" athleteid="6114">
              <RESULTS>
                <RESULT eventid="1076" points="230" reactiontime="+99" swimtime="00:00:33.05" resultid="6115" heatid="7254" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1188" points="278" reactiontime="+96" swimtime="00:21:37.90" resultid="6116" heatid="7303" lane="7" entrytime="00:22:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:02:00.57" />
                    <SPLIT distance="200" swimtime="00:02:42.43" />
                    <SPLIT distance="250" swimtime="00:03:24.98" />
                    <SPLIT distance="300" swimtime="00:04:07.81" />
                    <SPLIT distance="350" swimtime="00:04:51.04" />
                    <SPLIT distance="400" swimtime="00:05:33.96" />
                    <SPLIT distance="450" swimtime="00:06:16.77" />
                    <SPLIT distance="500" swimtime="00:06:59.56" />
                    <SPLIT distance="600" swimtime="00:08:26.48" />
                    <SPLIT distance="700" swimtime="00:09:54.72" />
                    <SPLIT distance="750" swimtime="00:10:38.66" />
                    <SPLIT distance="850" swimtime="00:12:07.37" />
                    <SPLIT distance="1000" swimtime="00:12:50.99" />
                    <SPLIT distance="1050" swimtime="00:15:01.12" />
                    <SPLIT distance="1200" swimtime="00:17:13.19" />
                    <SPLIT distance="1250" swimtime="00:17:57.73" />
                    <SPLIT distance="1300" swimtime="00:18:42.29" />
                    <SPLIT distance="1350" swimtime="00:19:27.18" />
                    <SPLIT distance="1400" swimtime="00:20:11.19" />
                    <SPLIT distance="1450" swimtime="00:20:56.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="250" reactiontime="+85" swimtime="00:01:11.28" resultid="6117" heatid="7355" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="252" reactiontime="+96" swimtime="00:02:37.31" resultid="6118" heatid="7480" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="183" reactiontime="+90" swimtime="00:03:05.77" resultid="6119" heatid="7532" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="252" reactiontime="+97" swimtime="00:05:36.03" resultid="6120" heatid="7579" lane="5" entrytime="00:05:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="150" swimtime="00:02:02.12" />
                    <SPLIT distance="200" swimtime="00:02:45.13" />
                    <SPLIT distance="250" swimtime="00:03:28.33" />
                    <SPLIT distance="350" swimtime="00:04:52.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-18" firstname="Danuta" gender="F" lastname="Wegen" nation="POL" athleteid="6200">
              <RESULTS>
                <RESULT eventid="1059" points="118" reactiontime="+84" swimtime="00:00:46.70" resultid="6201" heatid="7234" lane="3" />
                <RESULT eventid="1207" points="110" reactiontime="+99" swimtime="00:00:53.51" resultid="6202" heatid="7306" lane="3" />
                <RESULT eventid="1272" points="103" reactiontime="+100" swimtime="00:01:46.87" resultid="6203" heatid="7340" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="97" reactiontime="+93" swimtime="00:01:59.76" resultid="6204" heatid="7452" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="85" swimtime="00:04:10.87" resultid="6205" heatid="7468" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                    <SPLIT distance="100" swimtime="00:01:59.78" />
                    <SPLIT distance="150" swimtime="00:03:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="88" reactiontime="+93" swimtime="00:04:27.87" resultid="6206" heatid="7523" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.23" />
                    <SPLIT distance="100" swimtime="00:02:08.69" />
                    <SPLIT distance="150" swimtime="00:03:19.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="84" swimtime="00:08:53.42" resultid="6207" heatid="7572" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.27" />
                    <SPLIT distance="100" swimtime="00:02:01.89" />
                    <SPLIT distance="150" swimtime="00:03:11.24" />
                    <SPLIT distance="200" swimtime="00:04:20.30" />
                    <SPLIT distance="250" swimtime="00:05:29.89" />
                    <SPLIT distance="300" swimtime="00:06:40.57" />
                    <SPLIT distance="350" swimtime="00:07:49.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Zaleska" nation="POL" athleteid="6153">
              <RESULTS>
                <RESULT eventid="1092" points="355" reactiontime="+86" swimtime="00:02:52.09" resultid="6154" heatid="7273" lane="7" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="150" swimtime="00:02:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="378" reactiontime="+93" swimtime="00:21:11.09" resultid="6155" heatid="7300" lane="3" entrytime="00:21:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                    <SPLIT distance="200" swimtime="00:02:38.94" />
                    <SPLIT distance="250" swimtime="00:03:19.77" />
                    <SPLIT distance="300" swimtime="00:04:00.82" />
                    <SPLIT distance="350" swimtime="00:04:42.29" />
                    <SPLIT distance="400" swimtime="00:05:24.00" />
                    <SPLIT distance="450" swimtime="00:06:06.03" />
                    <SPLIT distance="500" swimtime="00:06:47.87" />
                    <SPLIT distance="550" swimtime="00:07:29.86" />
                    <SPLIT distance="600" swimtime="00:08:12.18" />
                    <SPLIT distance="650" swimtime="00:08:54.17" />
                    <SPLIT distance="700" swimtime="00:09:36.70" />
                    <SPLIT distance="750" swimtime="00:10:20.23" />
                    <SPLIT distance="800" swimtime="00:11:02.97" />
                    <SPLIT distance="850" swimtime="00:11:45.95" />
                    <SPLIT distance="900" swimtime="00:12:29.49" />
                    <SPLIT distance="950" swimtime="00:13:13.22" />
                    <SPLIT distance="1000" swimtime="00:13:56.99" />
                    <SPLIT distance="1050" swimtime="00:14:40.28" />
                    <SPLIT distance="1100" swimtime="00:15:23.65" />
                    <SPLIT distance="1150" swimtime="00:16:07.06" />
                    <SPLIT distance="1200" swimtime="00:16:49.88" />
                    <SPLIT distance="1250" swimtime="00:17:33.52" />
                    <SPLIT distance="1300" swimtime="00:18:17.28" />
                    <SPLIT distance="1350" swimtime="00:19:00.31" />
                    <SPLIT distance="1400" swimtime="00:19:44.07" />
                    <SPLIT distance="1450" swimtime="00:20:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="355" reactiontime="+81" swimtime="00:00:36.24" resultid="6156" heatid="7312" lane="9" entrytime="00:00:37.50" />
                <RESULT eventid="1336" points="389" reactiontime="+80" swimtime="00:02:43.84" resultid="6157" heatid="7393" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:02:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="374" reactiontime="+80" swimtime="00:00:33.81" resultid="6158" heatid="7431" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="1561" points="353" reactiontime="+85" swimtime="00:06:06.09" resultid="6159" heatid="8151" lane="7" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:20.02" />
                    <SPLIT distance="150" swimtime="00:02:08.25" />
                    <SPLIT distance="200" swimtime="00:02:55.36" />
                    <SPLIT distance="250" swimtime="00:03:47.57" />
                    <SPLIT distance="300" swimtime="00:04:40.19" />
                    <SPLIT distance="350" swimtime="00:05:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="367" reactiontime="+83" swimtime="00:01:16.27" resultid="6160" heatid="7510" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="380" reactiontime="+81" swimtime="00:05:22.92" resultid="6161" heatid="7568" lane="8" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:15.92" />
                    <SPLIT distance="150" swimtime="00:01:56.78" />
                    <SPLIT distance="200" swimtime="00:02:37.78" />
                    <SPLIT distance="250" swimtime="00:03:18.34" />
                    <SPLIT distance="300" swimtime="00:03:58.81" />
                    <SPLIT distance="350" swimtime="00:04:36.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-28" firstname="Maciej" gender="M" lastname="Zembrzuski" nation="POL" athleteid="6253">
              <RESULTS>
                <RESULT eventid="1108" points="436" reactiontime="+83" swimtime="00:02:24.57" resultid="6254" heatid="7284" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                    <SPLIT distance="150" swimtime="00:01:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="365" reactiontime="+85" swimtime="00:10:20.25" resultid="6255" heatid="7295" lane="3" entrytime="00:10:34.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                    <SPLIT distance="200" swimtime="00:02:24.70" />
                    <SPLIT distance="250" swimtime="00:03:02.82" />
                    <SPLIT distance="300" swimtime="00:03:41.32" />
                    <SPLIT distance="350" swimtime="00:04:20.59" />
                    <SPLIT distance="400" swimtime="00:04:59.66" />
                    <SPLIT distance="450" swimtime="00:05:39.91" />
                    <SPLIT distance="500" swimtime="00:06:20.39" />
                    <SPLIT distance="550" swimtime="00:07:00.53" />
                    <SPLIT distance="600" swimtime="00:07:40.62" />
                    <SPLIT distance="650" swimtime="00:08:20.83" />
                    <SPLIT distance="700" swimtime="00:09:01.25" />
                    <SPLIT distance="750" swimtime="00:09:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="574" reactiontime="+81" swimtime="00:00:54.06" resultid="6256" heatid="7365" lane="1" entrytime="00:00:57.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="605" reactiontime="+78" swimtime="00:00:25.71" resultid="6257" heatid="7450" lane="6" entrytime="00:00:26.35" />
                <RESULT eventid="1513" points="527" reactiontime="+79" swimtime="00:02:03.01" resultid="6258" heatid="7487" lane="2" entrytime="00:02:04.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="150" swimtime="00:01:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="6259" heatid="7521" lane="9" entrytime="00:01:01.01" />
                <RESULT eventid="1737" points="437" reactiontime="+82" swimtime="00:04:39.52" resultid="6260" heatid="7574" lane="7" entrytime="00:04:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:42.16" />
                    <SPLIT distance="200" swimtime="00:02:18.25" />
                    <SPLIT distance="250" swimtime="00:02:53.93" />
                    <SPLIT distance="300" swimtime="00:03:29.21" />
                    <SPLIT distance="350" swimtime="00:04:05.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-18" firstname="Jacek" gender="M" lastname="Łuczak" nation="POL" athleteid="6185">
              <RESULTS>
                <RESULT eventid="1076" points="389" reactiontime="+70" swimtime="00:00:27.75" resultid="6186" heatid="7261" lane="8" entrytime="00:00:28.03" />
                <RESULT eventid="1256" points="307" reactiontime="+73" swimtime="00:02:57.99" resultid="6187" heatid="7336" lane="5" entrytime="00:03:08.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:25.38" />
                    <SPLIT distance="150" swimtime="00:02:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="331" reactiontime="+71" swimtime="00:01:04.95" resultid="6188" heatid="7360" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="356" reactiontime="+67" swimtime="00:01:18.42" resultid="6189" heatid="7422" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="396" reactiontime="+71" swimtime="00:00:34.38" resultid="6190" heatid="7558" lane="1" entrytime="00:00:34.81" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="PSTRĄGI" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="547" reactiontime="+75" swimtime="00:01:50.55" resultid="6265" heatid="7406" lane="1" entrytime="00:01:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                    <SPLIT distance="100" swimtime="00:00:59.93" />
                    <SPLIT distance="150" swimtime="00:01:24.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6171" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6089" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="6253" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="6144" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="SANDACZE" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="527" reactiontime="+75" swimtime="00:01:41.23" resultid="6269" heatid="7496" lane="7" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="100" swimtime="00:00:51.04" />
                    <SPLIT distance="150" swimtime="00:01:17.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6089" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="6253" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6144" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="6171" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WĘGORZE" number="2">
              <RESULTS>
                <RESULT eventid="1391" points="357" reactiontime="+67" swimtime="00:02:07.46" resultid="6266" heatid="7405" lane="9" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:36.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6135" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6185" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="6232" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="6121" number="4" reactiontime="-6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="ŁOSOSIE" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="381" reactiontime="+80" swimtime="00:01:52.83" resultid="6270" heatid="7495" lane="9" entrytime="00:01:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:00:56.86" />
                    <SPLIT distance="150" swimtime="00:01:23.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6180" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="6135" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="6185" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="6191" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="KARPIE" number="3">
              <RESULTS>
                <RESULT eventid="1545" points="241" reactiontime="+83" swimtime="00:02:11.42" resultid="6271" heatid="7494" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="150" swimtime="00:01:37.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6121" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="6114" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="6105" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="6097" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="SUMY" number="3">
              <RESULTS>
                <RESULT eventid="1391" points="247" reactiontime="+66" swimtime="00:02:24.13" resultid="6267" heatid="7404" lane="8" entrytime="00:02:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:52.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6191" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="6097" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="6247" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="6114" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="PŁOTKI" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="404" reactiontime="+82" swimtime="00:02:07.02" resultid="6268" heatid="7491" lane="9" entrytime="00:02:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:02.25" />
                    <SPLIT distance="150" swimtime="00:01:34.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6128" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="6223" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="6153" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="6162" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="STYNKI" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="381" reactiontime="+77" swimtime="00:02:21.19" resultid="6264" heatid="7401" lane="0" entrytime="00:02:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6162" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6153" number="2" />
                    <RELAYPOSITION athleteid="6128" number="3" />
                    <RELAYPOSITION athleteid="6223" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="CIERNICZKI" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="509" reactiontime="+81" swimtime="00:02:00.72" resultid="6272" heatid="7565" lane="2" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:36.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6153" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="6171" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="6128" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="6253" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="OKONKI" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="494" reactiontime="+81" swimtime="00:01:51.11" resultid="6261" heatid="7289" lane="5" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                    <SPLIT distance="100" swimtime="00:00:49.87" />
                    <SPLIT distance="150" swimtime="00:01:22.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6253" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="6171" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="6153" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="6128" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="KIEŁBIKI" number="2">
              <RESULTS>
                <RESULT eventid="1705" points="425" reactiontime="+77" swimtime="00:02:08.12" resultid="6273" heatid="7564" lane="5" entrytime="00:02:11.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.94" />
                    <SPLIT distance="150" swimtime="00:01:36.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6162" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6089" number="2" />
                    <RELAYPOSITION athleteid="6144" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="6223" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="SZCZUPACZKI" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="399" reactiontime="+72" swimtime="00:01:59.30" resultid="6262" heatid="7288" lane="3" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:52.42" />
                    <SPLIT distance="150" swimtime="00:01:24.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6089" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6144" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="6223" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="6238" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="LESZCZYKI" number="3">
              <RESULTS>
                <RESULT eventid="1124" points="360" reactiontime="+67" swimtime="00:02:03.54" resultid="6263" heatid="7288" lane="8" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                    <SPLIT distance="100" swimtime="00:00:53.65" />
                    <SPLIT distance="150" swimtime="00:01:26.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6135" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="6232" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="6162" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="6208" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="ZŁOTE RYBKI" number="3">
              <RESULTS>
                <RESULT eventid="1705" points="251" reactiontime="+77" swimtime="00:02:32.66" resultid="6274" heatid="7563" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:57.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6191" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6097" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="6208" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="6238" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ASGDY" nation="POL" region="10" clubid="2897" name="AquaStars Gdynia">
          <CONTACT name="MARIUSZ GOLON" />
          <ATHLETES>
            <ATHLETE birthdate="1978-10-20" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="2898">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2899" heatid="7255" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1224" points="323" reactiontime="+77" swimtime="00:00:32.37" resultid="2900" heatid="7322" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="397" reactiontime="+82" swimtime="00:01:08.37" resultid="2901" heatid="7385" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="372" reactiontime="+80" swimtime="00:01:17.31" resultid="2902" heatid="7416" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="448" reactiontime="+79" swimtime="00:00:28.42" resultid="2903" heatid="7445" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1689" points="421" reactiontime="+82" swimtime="00:00:33.68" resultid="2904" heatid="7555" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AQUNI" nation="SVK" region="ZSO" clubid="4361" name="Aquatics Nitra">
          <ATHLETES>
            <ATHLETE birthdate="1994-09-06" firstname="Martina" gender="F" lastname="Bábiková" nation="SVK" license="SVK23949" athleteid="4377">
              <RESULTS>
                <RESULT eventid="1240" points="185" reactiontime="+97" swimtime="00:03:55.78" resultid="4378" heatid="7329" lane="7" entrytime="00:03:47.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:50.08" />
                    <SPLIT distance="150" swimtime="00:02:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="191" reactiontime="+97" swimtime="00:01:48.25" resultid="4379" heatid="7409" lane="4" entrytime="00:01:51.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="138" reactiontime="+98" swimtime="00:01:49.26" resultid="4380" heatid="7370" lane="9" entrytime="00:01:50.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="202" reactiontime="+90" swimtime="00:00:48.67" resultid="4381" heatid="7539" lane="6" entrytime="00:00:50.63" entrycourse="SCM" />
                <RESULT eventid="1721" points="161" reactiontime="+98" swimtime="00:07:09.67" resultid="4382" heatid="7570" lane="1" entrytime="00:07:18.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:42.68" />
                    <SPLIT distance="150" swimtime="00:02:38.04" />
                    <SPLIT distance="200" swimtime="00:03:33.01" />
                    <SPLIT distance="250" swimtime="00:04:27.65" />
                    <SPLIT distance="300" swimtime="00:05:22.47" />
                    <SPLIT distance="350" swimtime="00:06:17.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="149" swimtime="00:00:43.21" resultid="4383" heatid="7236" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-08" firstname="Karol" gender="M" lastname="Lacko" nation="SVK" license="SVK16793" athleteid="4390">
              <RESULTS>
                <RESULT eventid="1513" points="401" reactiontime="+81" swimtime="00:02:14.73" resultid="4391" heatid="7484" lane="2" entrytime="00:02:15.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="398" reactiontime="+88" swimtime="00:04:48.32" resultid="4392" heatid="7575" lane="7" entrytime="00:04:50.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:45.33" />
                    <SPLIT distance="200" swimtime="00:02:21.73" />
                    <SPLIT distance="250" swimtime="00:02:57.84" />
                    <SPLIT distance="300" swimtime="00:03:34.66" />
                    <SPLIT distance="350" swimtime="00:04:11.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="383" swimtime="00:10:10.53" resultid="4393" heatid="7294" lane="0" entrytime="00:10:19.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:48.60" />
                    <SPLIT distance="200" swimtime="00:02:26.48" />
                    <SPLIT distance="250" swimtime="00:03:04.12" />
                    <SPLIT distance="300" swimtime="00:03:41.85" />
                    <SPLIT distance="350" swimtime="00:04:19.40" />
                    <SPLIT distance="400" swimtime="00:04:57.18" />
                    <SPLIT distance="450" swimtime="00:05:35.98" />
                    <SPLIT distance="500" swimtime="00:06:14.95" />
                    <SPLIT distance="550" swimtime="00:06:54.06" />
                    <SPLIT distance="600" swimtime="00:07:33.75" />
                    <SPLIT distance="650" swimtime="00:08:13.27" />
                    <SPLIT distance="700" swimtime="00:08:52.95" />
                    <SPLIT distance="750" swimtime="00:09:32.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-08" firstname="Miroslav" gender="M" lastname="Ábel" nation="SVK" license="SVK12721" athleteid="4362" firstname.en="Abel" lastname.en="Miroslav">
              <RESULTS>
                <RESULT eventid="1108" points="401" reactiontime="+86" swimtime="00:02:28.63" resultid="4363" heatid="7284" lane="9" entrytime="00:02:26.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="371" reactiontime="+76" swimtime="00:02:47.08" resultid="4364" heatid="7338" lane="2" entrytime="00:02:46.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:04.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="424" reactiontime="+80" swimtime="00:01:06.90" resultid="4365" heatid="7388" lane="7" entrytime="00:01:06.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="392" reactiontime="+77" swimtime="00:01:15.95" resultid="4366" heatid="7424" lane="8" entrytime="00:01:15.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="400" reactiontime="+69" swimtime="00:00:29.50" resultid="4367" heatid="7446" lane="6" entrytime="00:00:29.47" entrycourse="SCM" />
                <RESULT eventid="1577" points="349" reactiontime="+85" swimtime="00:05:34.28" resultid="4368" heatid="8158" lane="0" entrytime="00:05:29.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:54.13" />
                    <SPLIT distance="200" swimtime="00:02:35.87" />
                    <SPLIT distance="250" swimtime="00:03:23.33" />
                    <SPLIT distance="300" swimtime="00:04:11.71" />
                    <SPLIT distance="350" swimtime="00:04:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="402" reactiontime="+84" swimtime="00:01:05.11" resultid="4369" heatid="7520" lane="1" entrytime="00:01:03.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="398" reactiontime="+74" swimtime="00:00:34.31" resultid="4370" heatid="7559" lane="9" entrytime="00:00:33.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-01" firstname="Lucia" gender="F" lastname="Ábelová" nation="SVK" license="SVK19294" athleteid="4371">
              <RESULTS>
                <RESULT eventid="1059" points="145" reactiontime="+92" swimtime="00:00:43.61" resultid="4372" heatid="7237" lane="6" entrytime="00:00:41.86" entrycourse="SCM" />
                <RESULT eventid="1207" points="114" reactiontime="+84" swimtime="00:00:52.81" resultid="4373" heatid="7308" lane="4" entrytime="00:00:53.57" entrycourse="LCM" />
                <RESULT eventid="1304" points="145" swimtime="00:01:47.42" resultid="4374" heatid="7369" lane="4" entrytime="00:01:50.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="104" reactiontime="+98" swimtime="00:00:51.70" resultid="4375" heatid="7427" lane="7" entrytime="00:00:52.67" entrycourse="SCM" />
                <RESULT eventid="1673" points="219" reactiontime="+89" swimtime="00:00:47.31" resultid="4376" heatid="7539" lane="3" entrytime="00:00:50.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-02-03" firstname="Peter" gender="M" lastname="Čigáš" nation="SVK" license="SVK15844" athleteid="4384">
              <RESULTS>
                <RESULT eventid="1076" points="398" reactiontime="+88" swimtime="00:00:27.54" resultid="4385" heatid="7263" lane="5" entrytime="00:00:27.22" entrycourse="SCM" />
                <RESULT eventid="1224" points="368" reactiontime="+72" swimtime="00:00:30.99" resultid="4386" heatid="7325" lane="8" entrytime="00:00:31.07" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4387" heatid="7362" lane="1" entrytime="00:01:00.89" entrycourse="SCM" />
                <RESULT eventid="1481" points="388" reactiontime="+77" swimtime="00:01:06.96" resultid="4388" heatid="7466" lane="5" entrytime="00:01:05.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="342" reactiontime="+78" swimtime="00:02:30.96" resultid="4389" heatid="7535" lane="6" entrytime="00:02:26.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:52.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZRAC" nation="POL" region="11" clubid="2114" name="AZS PWSZ Racibórz">
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="2115">
              <RESULTS>
                <RESULT eventid="1108" points="194" reactiontime="+93" swimtime="00:03:09.10" resultid="2116" heatid="7279" lane="4" entrytime="00:03:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:24.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="185" reactiontime="+98" swimtime="00:03:30.83" resultid="2117" heatid="7335" lane="3" entrytime="00:03:23.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:41.14" />
                    <SPLIT distance="150" swimtime="00:02:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="148" swimtime="00:03:24.32" resultid="2118" heatid="7396" lane="7" entrytime="00:03:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:37.40" />
                    <SPLIT distance="150" swimtime="00:02:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="222" reactiontime="+92" swimtime="00:01:31.72" resultid="2119" heatid="7419" lane="2" entrytime="00:01:30.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="185" swimtime="00:06:52.97" resultid="2120" heatid="8156" lane="1" entrytime="00:06:45.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:40.58" />
                    <SPLIT distance="150" swimtime="00:02:34.86" />
                    <SPLIT distance="200" swimtime="00:03:26.76" />
                    <SPLIT distance="250" swimtime="00:04:23.18" />
                    <SPLIT distance="300" swimtime="00:05:18.99" />
                    <SPLIT distance="350" swimtime="00:06:06.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="150" reactiontime="+97" swimtime="00:01:30.38" resultid="2121" heatid="7515" lane="2" entrytime="00:01:30.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="239" reactiontime="+90" swimtime="00:00:40.65" resultid="2122" heatid="7552" lane="8" entrytime="00:00:40.55" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZKIE" nation="POL" region="12" clubid="2769" name="AZS UJK Kielce">
          <ATHLETES>
            <ATHLETE birthdate="1996-11-24" firstname="Paulina" gender="F" lastname="Majos" nation="POL" athleteid="2768">
              <RESULTS>
                <RESULT eventid="1059" points="405" reactiontime="+82" swimtime="00:00:30.97" resultid="2770" heatid="7242" lane="4" entrytime="00:00:31.20" />
                <RESULT eventid="1140" points="425" reactiontime="+86" swimtime="00:10:37.42" resultid="2771" heatid="7290" lane="7" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                    <SPLIT distance="200" swimtime="00:02:29.87" />
                    <SPLIT distance="250" swimtime="00:03:09.86" />
                    <SPLIT distance="300" swimtime="00:03:50.44" />
                    <SPLIT distance="350" swimtime="00:04:31.15" />
                    <SPLIT distance="400" swimtime="00:05:12.25" />
                    <SPLIT distance="450" swimtime="00:05:53.12" />
                    <SPLIT distance="500" swimtime="00:06:34.09" />
                    <SPLIT distance="550" swimtime="00:07:15.11" />
                    <SPLIT distance="600" swimtime="00:07:56.23" />
                    <SPLIT distance="650" swimtime="00:08:37.02" />
                    <SPLIT distance="700" swimtime="00:09:17.76" />
                    <SPLIT distance="750" swimtime="00:09:58.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BPMYS" nation="POL" region="11" clubid="2329" name="Baza Pływania Mysłowice">
          <CONTACT city="Mysłowice" email="kisielmonika@onet.pl" name="Kisiel" phone="511987305" street="Stawowa" zip="41-400" />
          <ATHLETES>
            <ATHLETE birthdate="1996-05-27" firstname="Monika" gender="F" lastname="Kisiel" nation="POL" athleteid="2330">
              <RESULTS>
                <RESULT eventid="1207" points="470" reactiontime="+77" swimtime="00:00:33.01" resultid="2331" heatid="7313" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1465" points="454" reactiontime="+80" swimtime="00:01:11.57" resultid="2332" heatid="7458" lane="8" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="429" reactiontime="+75" swimtime="00:02:38.07" resultid="2333" heatid="7528" lane="6" entrytime="00:02:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CMUJKR" nation="POL" region="06" clubid="6302" name="Collegium Medicum UJ Masters Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT email="mariuszbaranik@gmail.com" name="Mariusz Baranik" phone="69812822" state="MAL" street="Białopradnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="6303">
              <RESULTS>
                <RESULT eventid="1076" points="474" reactiontime="+75" swimtime="00:00:25.97" resultid="6304" heatid="7264" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1288" points="467" reactiontime="+77" swimtime="00:00:57.92" resultid="6305" heatid="7363" lane="7" entrytime="00:00:59.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="410" reactiontime="+78" swimtime="00:01:07.61" resultid="6306" heatid="7387" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="6307" heatid="7423" lane="7" entrytime="00:01:18.00" />
                <RESULT eventid="1449" points="454" reactiontime="+72" swimtime="00:00:28.29" resultid="6308" heatid="7447" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1625" points="380" reactiontime="+75" swimtime="00:01:06.36" resultid="6309" heatid="7519" lane="0" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="420" reactiontime="+69" swimtime="00:00:33.69" resultid="6310" heatid="7557" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="6492">
              <RESULTS>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="6494" heatid="7304" lane="3" entrytime="00:24:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="11" clubid="4184" name="CSiR MOS Dąbrowa Grn.">
          <CONTACT email="mariuszwaliczek@interia.pl" name="Waliczek Mariusz" />
          <ATHLETES>
            <ATHLETE birthdate="1997-10-21" firstname="Patryk" gender="M" lastname="Droś" nation="POL" athleteid="4185">
              <RESULTS>
                <RESULT eventid="1288" points="648" reactiontime="+68" swimtime="00:00:51.91" resultid="4186" heatid="7367" lane="2" entrytime="00:00:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="583" reactiontime="+71" swimtime="00:01:00.14" resultid="4187" heatid="7390" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="626" reactiontime="+69" swimtime="00:01:05.00" resultid="4188" heatid="7425" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="580" reactiontime="+71" swimtime="00:01:59.12" resultid="4189" heatid="7488" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                    <SPLIT distance="150" swimtime="00:01:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="695" reactiontime="+69" swimtime="00:00:28.50" resultid="4190" heatid="7561" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-03-23" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="4207">
              <RESULTS>
                <RESULT eventid="1224" points="348" reactiontime="+66" swimtime="00:00:31.59" resultid="4208" heatid="7326" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="4209" heatid="7394" lane="8" />
                <RESULT eventid="1481" points="350" reactiontime="+71" swimtime="00:01:09.32" resultid="4210" heatid="7465" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="4211" heatid="8153" lane="9" />
                <RESULT eventid="1657" points="253" reactiontime="+73" swimtime="00:02:46.86" resultid="4212" heatid="7534" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-01" firstname="Dawid" gender="M" lastname="Nowodworski" nation="POL" license="102711200028" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1076" points="646" reactiontime="+83" swimtime="00:00:23.43" resultid="4200" heatid="7270" lane="5" entrytime="00:00:23.00" />
                <RESULT eventid="1224" points="588" reactiontime="+78" swimtime="00:00:26.52" resultid="4201" heatid="7326" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1320" points="677" reactiontime="+77" swimtime="00:00:57.22" resultid="4202" heatid="7390" lane="5" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="683" reactiontime="+78" swimtime="00:01:03.14" resultid="4203" heatid="7425" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="695" reactiontime="+72" swimtime="00:00:24.55" resultid="4204" heatid="7451" lane="6" entrytime="00:00:24.80" />
                <RESULT eventid="1625" points="619" reactiontime="+76" swimtime="00:00:56.39" resultid="4205" heatid="7522" lane="1" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="709" reactiontime="+70" swimtime="00:00:28.31" resultid="4206" heatid="7561" lane="3" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-08-24" firstname="Wiktoria" gender="F" lastname="Szlachcic" nation="POL" athleteid="4213">
              <RESULTS>
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="4214" heatid="7313" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1240" points="333" reactiontime="+82" swimtime="00:03:14.06" resultid="4215" heatid="7327" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4216" heatid="7473" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="1561" points="301" reactiontime="+83" swimtime="00:06:26.13" resultid="4217" heatid="8149" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:15.55" />
                    <SPLIT distance="200" swimtime="00:03:05.23" />
                    <SPLIT distance="250" swimtime="00:04:00.61" />
                    <SPLIT distance="300" swimtime="00:04:55.93" />
                    <SPLIT distance="350" swimtime="00:05:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="4218" heatid="7528" lane="8" entrytime="00:02:40.00" />
                <RESULT eventid="1721" points="329" reactiontime="+92" swimtime="00:05:38.53" resultid="4219" heatid="7572" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                    <SPLIT distance="200" swimtime="00:02:43.37" />
                    <SPLIT distance="250" swimtime="00:03:26.66" />
                    <SPLIT distance="300" swimtime="00:04:10.79" />
                    <SPLIT distance="350" swimtime="00:04:55.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-22" firstname="Anna" gender="F" lastname="Teresko" nation="POL" athleteid="4191">
              <RESULTS>
                <RESULT eventid="1207" points="551" reactiontime="+76" swimtime="00:00:31.30" resultid="4192" heatid="7314" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="4193" heatid="7376" lane="2" entrytime="00:01:08.00" />
                <RESULT eventid="1336" points="532" reactiontime="+80" swimtime="00:02:27.59" resultid="4194" heatid="7393" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                    <SPLIT distance="150" swimtime="00:01:48.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="545" reactiontime="+78" swimtime="00:01:07.37" resultid="4195" heatid="7458" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="648" reactiontime="+68" swimtime="00:02:07.61" resultid="4196" heatid="7474" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="100" swimtime="00:01:02.44" />
                    <SPLIT distance="150" swimtime="00:01:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="568" reactiontime="+70" swimtime="00:01:05.92" resultid="4197" heatid="7511" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="535" reactiontime="+77" swimtime="00:02:26.87" resultid="4198" heatid="7528" lane="4" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEGLI" nation="POL" region="11" clubid="2503" name="Delfin 92 Gliwice">
          <CONTACT email="cupialsport@op.pl" name="Cupiał" phone="605065587" />
          <ATHLETES>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="2504">
              <RESULTS>
                <RESULT eventid="1076" points="35" reactiontime="+79" swimtime="00:01:01.39" resultid="2505" heatid="7247" lane="2" entrytime="00:01:06.38" />
                <RESULT eventid="1224" points="27" swimtime="00:01:13.41" resultid="2506" heatid="7316" lane="2" entrytime="00:01:16.28" />
                <RESULT eventid="1256" points="42" reactiontime="+92" swimtime="00:05:43.21" resultid="2507" heatid="7332" lane="6" entrytime="00:05:56.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.65" />
                    <SPLIT distance="100" swimtime="00:02:42.14" />
                    <SPLIT distance="150" swimtime="00:04:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="48" swimtime="00:02:32.65" resultid="2508" heatid="7415" lane="1" entrytime="00:02:33.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="22" swimtime="00:02:51.90" resultid="2509" heatid="7460" lane="9" entrytime="00:02:44.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="30" swimtime="00:05:36.26" resultid="2510" heatid="7529" lane="6" entrytime="00:05:48.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.22" />
                    <SPLIT distance="100" swimtime="00:02:43.06" />
                    <SPLIT distance="150" swimtime="00:04:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="64" reactiontime="+99" swimtime="00:01:03.04" resultid="2511" heatid="7547" lane="9" entrytime="00:01:05.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00105" nation="POL" region="05" clubid="3609" name="Delfin Masters Łódz">
          <CONTACT email="cewa@poczta.fm" name="Ewa Kadłubiec" phone="604627966" />
          <ATHLETES>
            <ATHLETE birthdate="1971-02-25" firstname="Jacek" gender="M" lastname="Kadłubiec" nation="POL" athleteid="3610">
              <RESULTS>
                <RESULT eventid="1256" points="288" reactiontime="+87" swimtime="00:03:01.88" resultid="3611" heatid="7337" lane="4" entrytime="00:02:57.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="299" reactiontime="+91" swimtime="00:01:23.10" resultid="3612" heatid="7422" lane="9" entrytime="00:01:20.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-15" firstname="Grzegorz" gender="M" lastname="Kędziora" nation="POL" athleteid="3622">
              <RESULTS>
                <RESULT eventid="1449" points="383" reactiontime="+88" swimtime="00:00:29.94" resultid="3623" heatid="7439" lane="9" entrytime="00:00:38.13" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="3624" heatid="7515" lane="6" entrytime="00:01:30.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-14" firstname="Piotr" gender="M" lastname="Lewiński" nation="POL" athleteid="3618">
              <RESULTS>
                <RESULT eventid="1156" points="172" reactiontime="+99" swimtime="00:13:16.22" resultid="3619" heatid="7298" lane="4" entrytime="00:12:30.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:26.80" />
                    <SPLIT distance="150" swimtime="00:02:14.27" />
                    <SPLIT distance="200" swimtime="00:03:03.66" />
                    <SPLIT distance="250" swimtime="00:03:54.06" />
                    <SPLIT distance="300" swimtime="00:04:43.73" />
                    <SPLIT distance="450" swimtime="00:07:16.02" />
                    <SPLIT distance="600" swimtime="00:09:51.52" />
                    <SPLIT distance="650" swimtime="00:10:42.43" />
                    <SPLIT distance="750" swimtime="00:12:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="142" reactiontime="+88" swimtime="00:00:42.54" resultid="3620" heatid="7318" lane="5" entrytime="00:00:45.13" />
                <RESULT eventid="1513" points="202" reactiontime="+93" swimtime="00:02:49.35" resultid="3621" heatid="7479" lane="1" entrytime="00:02:50.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:05.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-05-06" firstname="Krzysztof" gender="M" lastname="Połomka" nation="POL" athleteid="3613">
              <RESULTS>
                <RESULT eventid="1076" points="279" reactiontime="+84" swimtime="00:00:30.98" resultid="3614" heatid="7256" lane="3" entrytime="00:00:31.18" />
                <RESULT eventid="1224" points="202" reactiontime="+77" swimtime="00:00:37.83" resultid="3615" heatid="7320" lane="4" entrytime="00:00:38.01" />
                <RESULT eventid="1288" points="259" reactiontime="+84" swimtime="00:01:10.45" resultid="3616" heatid="7356" lane="9" entrytime="00:01:11.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="212" reactiontime="+76" swimtime="00:01:21.85" resultid="3617" heatid="7462" lane="3" entrytime="00:01:30.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Grzegorz" gender="M" lastname="Rogalski" nation="POL" athleteid="3632">
              <RESULTS>
                <RESULT eventid="1076" points="396" reactiontime="+87" swimtime="00:00:27.57" resultid="3633" heatid="7257" lane="2" entrytime="00:00:30.13" />
                <RESULT eventid="1224" points="274" reactiontime="+79" swimtime="00:00:34.17" resultid="3634" heatid="7321" lane="3" entrytime="00:00:36.13" />
                <RESULT eventid="1449" points="370" reactiontime="+73" swimtime="00:00:30.27" resultid="3635" heatid="7441" lane="3" entrytime="00:00:33.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-08" firstname="Tomasz" gender="M" lastname="Wiaderny" nation="POL" athleteid="3625">
              <RESULTS>
                <RESULT eventid="1076" points="201" reactiontime="+78" swimtime="00:00:34.54" resultid="3626" heatid="7251" lane="6" entrytime="00:00:36.93" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3627" heatid="7319" lane="4" entrytime="00:00:41.36" />
                <RESULT eventid="1288" points="166" reactiontime="+95" swimtime="00:01:21.70" resultid="3656" heatid="7350" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="349" reactiontime="+82" swimtime="00:01:56.11" resultid="3638" heatid="7492" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:00:58.29" />
                    <SPLIT distance="150" swimtime="00:01:28.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3622" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3613" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3610" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3632" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RSUSZ" nation="HUN" clubid="5911" name="Dr. Regele Szenior Úszóklub">
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Ferenc" gender="M" lastname="Bagdi" nation="HUN" athleteid="5910">
              <RESULTS>
                <RESULT eventid="1108" points="347" reactiontime="+91" swimtime="00:02:35.88" resultid="5912" heatid="7282" lane="5" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:59.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="314" reactiontime="+93" swimtime="00:10:52.21" resultid="5913" heatid="7295" lane="9" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:49.73" />
                    <SPLIT distance="200" swimtime="00:02:29.90" />
                    <SPLIT distance="250" swimtime="00:03:10.38" />
                    <SPLIT distance="300" swimtime="00:03:51.56" />
                    <SPLIT distance="350" swimtime="00:04:32.87" />
                    <SPLIT distance="400" swimtime="00:05:14.44" />
                    <SPLIT distance="450" swimtime="00:05:55.85" />
                    <SPLIT distance="500" swimtime="00:06:37.56" />
                    <SPLIT distance="550" swimtime="00:07:19.52" />
                    <SPLIT distance="600" swimtime="00:08:02.18" />
                    <SPLIT distance="650" swimtime="00:08:45.03" />
                    <SPLIT distance="700" swimtime="00:09:27.43" />
                    <SPLIT distance="750" swimtime="00:10:10.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="389" reactiontime="+78" swimtime="00:01:01.56" resultid="5914" heatid="7359" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="357" reactiontime="+81" swimtime="00:01:10.82" resultid="5915" heatid="7385" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="327" reactiontime="+81" swimtime="00:01:20.67" resultid="5916" heatid="7420" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="361" reactiontime="+84" swimtime="00:02:19.44" resultid="5917" heatid="7483" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:41.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DSPDA" nation="POL" region="11" clubid="5896" name="Dąbrowska Szkoła Pływania">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="5895">
              <RESULTS>
                <RESULT eventid="1224" points="228" reactiontime="+70" swimtime="00:00:36.37" resultid="5897" heatid="7318" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1256" points="305" reactiontime="+83" swimtime="00:02:58.33" resultid="5898" heatid="7333" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:23.87" />
                    <SPLIT distance="150" swimtime="00:02:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="361" reactiontime="+82" swimtime="00:01:18.08" resultid="5899" heatid="7416" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="252" reactiontime="+75" swimtime="00:01:17.38" resultid="5900" heatid="7461" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5901" heatid="7530" lane="3" entrytime="00:04:00.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5902" heatid="7550" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-03-24" firstname="Kinga" gender="F" lastname="Pluta" nation="POL" athleteid="5903">
              <RESULTS>
                <RESULT eventid="1207" points="307" reactiontime="+82" swimtime="00:00:38.04" resultid="5904" heatid="7309" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1240" points="370" reactiontime="+86" swimtime="00:03:07.29" resultid="5905" heatid="7329" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:16.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="414" reactiontime="+86" swimtime="00:01:23.66" resultid="5906" heatid="7409" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="414" reactiontime="+80" swimtime="00:00:32.70" resultid="5907" heatid="7428" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="5908" heatid="7525" lane="1" entrytime="00:04:00.00" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5909" heatid="7541" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EULVI" nation="UKR" clubid="4239" name="Euro Lviv">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua, riff.lviv@gmail.com" fax="+48 537 723 854" internet="www.mastersswim.com.ua" name="Ruslan Friauf" phone="+38 067 673 4796" zip="79000" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-29" firstname="Sergii" gender="M" lastname="Abdulaiev" nation="UKR" athleteid="4240">
              <RESULTS>
                <RESULT eventid="1076" points="468" swimtime="00:00:26.08" resultid="4241" heatid="7268" lane="0" entrytime="00:00:25.50" />
                <RESULT eventid="1224" points="477" reactiontime="+72" swimtime="00:00:28.43" resultid="4242" heatid="7326" lane="2" entrytime="00:00:28.90" />
                <RESULT eventid="1320" points="474" reactiontime="+84" swimtime="00:01:04.44" resultid="4243" heatid="7389" lane="7" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="460" reactiontime="+83" swimtime="00:01:03.32" resultid="4244" heatid="7467" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="407" reactiontime="+85" swimtime="00:00:34.07" resultid="4245" heatid="7560" lane="8" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="4274">
              <RESULTS>
                <RESULT eventid="1224" points="177" reactiontime="+90" swimtime="00:00:39.55" resultid="4275" heatid="7320" lane="2" entrytime="00:00:39.50" />
                <RESULT eventid="1320" points="229" reactiontime="+89" swimtime="00:01:22.04" resultid="4276" heatid="7381" lane="5" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="4277" heatid="7463" lane="9" entrytime="00:01:27.50" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="4278" heatid="7532" lane="9" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-18" firstname="Vladyslav" gender="M" lastname="Horovoy" nation="UKR" athleteid="4259">
              <RESULTS>
                <RESULT eventid="1108" points="515" reactiontime="+74" swimtime="00:02:16.70" resultid="4260" heatid="7285" lane="1" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="546" reactiontime="+76" swimtime="00:02:27.01" resultid="4261" heatid="7339" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:09.90" />
                    <SPLIT distance="150" swimtime="00:01:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="544" reactiontime="+77" swimtime="00:01:01.56" resultid="4262" heatid="7389" lane="1" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="593" reactiontime="+71" swimtime="00:01:06.19" resultid="4263" heatid="7425" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="505" reactiontime="+73" swimtime="00:02:04.76" resultid="4264" heatid="7487" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="100" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="572" reactiontime="+69" swimtime="00:00:30.41" resultid="4265" heatid="7560" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="4266" heatid="7573" lane="3" entrytime="00:04:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="4252">
              <RESULTS>
                <RESULT eventid="1076" points="485" reactiontime="+69" swimtime="00:00:25.77" resultid="4253" heatid="7266" lane="4" entrytime="00:00:26.25" />
                <RESULT eventid="1156" points="344" reactiontime="+75" swimtime="00:10:32.84" resultid="4254" heatid="7295" lane="8" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                    <SPLIT distance="200" swimtime="00:02:26.95" />
                    <SPLIT distance="250" swimtime="00:03:06.29" />
                    <SPLIT distance="300" swimtime="00:03:46.25" />
                    <SPLIT distance="350" swimtime="00:04:26.60" />
                    <SPLIT distance="400" swimtime="00:05:06.53" />
                    <SPLIT distance="450" swimtime="00:05:46.73" />
                    <SPLIT distance="500" swimtime="00:06:27.29" />
                    <SPLIT distance="550" swimtime="00:07:07.48" />
                    <SPLIT distance="600" swimtime="00:07:48.77" />
                    <SPLIT distance="650" swimtime="00:08:29.81" />
                    <SPLIT distance="700" swimtime="00:09:11.11" />
                    <SPLIT distance="750" swimtime="00:09:52.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="478" reactiontime="+74" swimtime="00:00:57.46" resultid="4255" heatid="7364" lane="0" entrytime="00:00:58.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="403" reactiontime="+70" swimtime="00:00:29.43" resultid="4256" heatid="7446" lane="9" entrytime="00:00:29.85" />
                <RESULT eventid="1689" points="453" reactiontime="+71" swimtime="00:00:32.87" resultid="4257" heatid="7559" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1737" points="368" reactiontime="+72" swimtime="00:04:55.97" resultid="4258" heatid="7577" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:10.51" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                    <SPLIT distance="200" swimtime="00:02:26.91" />
                    <SPLIT distance="250" swimtime="00:03:05.02" />
                    <SPLIT distance="300" swimtime="00:03:42.72" />
                    <SPLIT distance="350" swimtime="00:04:20.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-02-27" firstname="Olena" gender="F" lastname="Pereyaslova" nation="UKR" athleteid="4267">
              <RESULTS>
                <RESULT eventid="1059" points="304" reactiontime="+99" swimtime="00:00:34.08" resultid="4268" heatid="7240" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1272" points="286" reactiontime="+88" swimtime="00:01:16.19" resultid="4269" heatid="7344" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="196" reactiontime="+93" swimtime="00:01:47.30" resultid="4270" heatid="7410" lane="5" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="252" reactiontime="+92" swimtime="00:02:54.63" resultid="4271" heatid="7471" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="204" reactiontime="+79" swimtime="00:00:48.51" resultid="4272" heatid="7540" lane="0" entrytime="00:00:48.00" />
                <RESULT eventid="1721" points="243" reactiontime="+90" swimtime="00:06:14.62" resultid="4273" heatid="7569" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:15.52" />
                    <SPLIT distance="200" swimtime="00:03:04.14" />
                    <SPLIT distance="250" swimtime="00:03:52.59" />
                    <SPLIT distance="300" swimtime="00:04:41.42" />
                    <SPLIT distance="350" swimtime="00:05:29.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="4246">
              <RESULTS>
                <RESULT eventid="1076" points="471" reactiontime="+88" swimtime="00:00:26.03" resultid="4247" heatid="7267" lane="5" entrytime="00:00:25.73" />
                <RESULT eventid="1288" points="467" reactiontime="+83" swimtime="00:00:57.92" resultid="4248" heatid="7364" lane="2" entrytime="00:00:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="413" reactiontime="+80" swimtime="00:02:25.32" resultid="4249" heatid="7398" lane="7" entrytime="00:02:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="504" reactiontime="+77" swimtime="00:00:27.32" resultid="4250" heatid="7449" lane="3" entrytime="00:00:27.34" />
                <RESULT eventid="1625" points="439" reactiontime="+89" swimtime="00:01:03.25" resultid="4251" heatid="7520" lane="0" entrytime="00:01:03.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="527" reactiontime="+84" swimtime="00:01:51.91" resultid="4279" heatid="7406" lane="2" entrytime="00:01:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                    <SPLIT distance="150" swimtime="00:01:26.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4240" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4259" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4246" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4252" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="496" reactiontime="+75" swimtime="00:01:43.29" resultid="4280" heatid="7496" lane="2" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.59" />
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="150" swimtime="00:01:17.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4259" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4252" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="4240" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4246" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11314" nation="POL" region="14" clubid="2773" name="Fundacja Hasten Warszawa " shortname="Hasten Warszawa ">
          <CONTACT email="hasten@hasten.pl" name="Bochyńska-Knapik Sonia" phone="507929874" />
          <ATHLETES>
            <ATHLETE birthdate="1993-01-10" firstname="Magdalena" gender="F" lastname="Baranowska" nation="POL" athleteid="2776">
              <RESULTS>
                <RESULT eventid="1059" points="530" reactiontime="+88" swimtime="00:00:28.32" resultid="2777" heatid="7245" lane="2" entrytime="00:00:27.49" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2778" heatid="7348" lane="6" entrytime="00:00:59.99" />
                <RESULT eventid="1433" points="511" reactiontime="+79" swimtime="00:00:30.49" resultid="2779" heatid="7434" lane="2" entrytime="00:00:29.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-10" firstname="Sonia" gender="F" lastname="Bochyńska-Knapik" nation="POL" athleteid="2780">
              <RESULTS>
                <RESULT eventid="1207" points="536" reactiontime="+70" swimtime="00:00:31.60" resultid="2781" heatid="7314" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1433" points="518" reactiontime="+71" swimtime="00:00:30.34" resultid="2782" heatid="7434" lane="9" entrytime="00:00:30.50" />
                <RESULT eventid="1465" points="461" reactiontime="+67" swimtime="00:01:11.23" resultid="2783" heatid="7458" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-20" firstname="Mirela" gender="F" lastname="Olczak" nation="POL" athleteid="2784">
              <RESULTS>
                <RESULT eventid="1304" points="522" reactiontime="+72" swimtime="00:01:10.16" resultid="2785" heatid="7376" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="543" reactiontime="+72" swimtime="00:00:29.87" resultid="2786" heatid="7434" lane="3" entrytime="00:00:29.49" />
                <RESULT eventid="1608" points="492" reactiontime="+71" swimtime="00:01:09.17" resultid="2787" heatid="7511" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-04" firstname="Natalia" gender="F" lastname="Pawlaczek" nation="POL" athleteid="2774">
              <RESULTS>
                <RESULT eventid="1272" points="648" reactiontime="+74" swimtime="00:00:58.05" resultid="2775" heatid="7348" lane="4" entrytime="00:00:58.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="TEAM HASTEN &apos;90" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="590" reactiontime="+77" swimtime="00:01:51.96" resultid="2788" heatid="7491" lane="4" entrytime="00:01:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:00:57.38" />
                    <SPLIT distance="150" swimtime="00:01:25.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2776" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2784" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2780" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2774" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="542" reactiontime="+64" swimtime="00:02:05.56" resultid="2789" heatid="7401" lane="4" entrytime="00:02:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:39.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2780" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2776" number="2" />
                    <RELAYPOSITION athleteid="2784" number="3" />
                    <RELAYPOSITION athleteid="2774" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAGDY" nation="POL" region="10" clubid="4055" name="Gdynia Masters">
          <CONTACT name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Jan" gender="M" lastname="Boboli" nation="POL" athleteid="4064">
              <RESULTS>
                <RESULT eventid="1076" points="154" reactiontime="+86" swimtime="00:00:37.73" resultid="4065" heatid="7250" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1224" points="39" reactiontime="+87" swimtime="00:01:05.22" resultid="4066" heatid="7317" lane="0" entrytime="00:01:00.00" />
                <RESULT eventid="1689" points="46" reactiontime="+90" swimtime="00:01:10.41" resultid="4067" heatid="7547" lane="7" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="4129">
              <RESULTS>
                <RESULT eventid="1059" points="84" swimtime="00:00:52.33" resultid="4130" heatid="7235" lane="7" entrytime="00:00:57.00" />
                <RESULT eventid="1207" points="80" reactiontime="+72" swimtime="00:00:59.41" resultid="4131" heatid="7307" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="1465" points="70" reactiontime="+82" swimtime="00:02:12.97" resultid="4132" heatid="7453" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="68" reactiontime="+73" swimtime="00:04:50.89" resultid="4133" heatid="7524" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.94" />
                    <SPLIT distance="100" swimtime="00:02:23.68" />
                    <SPLIT distance="150" swimtime="00:03:38.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Ewa" gender="F" lastname="Gawlik" nation="POL" athleteid="4120">
              <RESULTS>
                <RESULT eventid="1059" points="154" swimtime="00:00:42.75" resultid="4121" heatid="7236" lane="4" entrytime="00:00:43.20" />
                <RESULT comment="Rekord Polski Masters kategoria J" eventid="1140" points="145" reactiontime="+86" swimtime="00:15:11.93" resultid="4122" heatid="7292" lane="1" entrytime="00:15:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.06" />
                    <SPLIT distance="100" swimtime="00:01:45.61" />
                    <SPLIT distance="150" swimtime="00:02:43.13" />
                    <SPLIT distance="200" swimtime="00:03:40.97" />
                    <SPLIT distance="250" swimtime="00:04:38.05" />
                    <SPLIT distance="300" swimtime="00:05:35.91" />
                    <SPLIT distance="350" swimtime="00:06:33.59" />
                    <SPLIT distance="400" swimtime="00:07:31.05" />
                    <SPLIT distance="450" swimtime="00:08:28.37" />
                    <SPLIT distance="500" swimtime="00:09:25.78" />
                    <SPLIT distance="550" swimtime="00:10:23.66" />
                    <SPLIT distance="600" swimtime="00:11:21.24" />
                    <SPLIT distance="650" swimtime="00:12:19.67" />
                    <SPLIT distance="700" swimtime="00:13:18.04" />
                    <SPLIT distance="750" swimtime="00:14:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="139" reactiontime="+96" swimtime="00:01:36.93" resultid="4123" heatid="7342" lane="8" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="121" reactiontime="+95" swimtime="00:01:54.12" resultid="4124" heatid="7369" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="113" reactiontime="+82" swimtime="00:00:50.40" resultid="4125" heatid="7427" lane="3" entrytime="00:00:50.50" />
                <RESULT eventid="1497" points="132" reactiontime="+89" swimtime="00:03:36.59" resultid="4126" heatid="7469" lane="1" entrytime="00:03:34.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:43.34" />
                    <SPLIT distance="150" swimtime="00:02:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="99" reactiontime="+93" swimtime="00:01:57.77" resultid="4127" heatid="7508" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="147" reactiontime="+93" swimtime="00:07:22.28" resultid="4128" heatid="7570" lane="9" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                    <SPLIT distance="150" swimtime="00:02:38.66" />
                    <SPLIT distance="200" swimtime="00:03:34.53" />
                    <SPLIT distance="250" swimtime="00:04:31.23" />
                    <SPLIT distance="300" swimtime="00:05:28.19" />
                    <SPLIT distance="350" swimtime="00:06:25.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="4088">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="4089" heatid="7237" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="4090" heatid="7308" lane="1" entrytime="00:00:57.00" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="4091" heatid="7369" lane="8" entrytime="00:02:08.00" />
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="4092" heatid="7408" lane="5" entrytime="00:02:09.00" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4093" heatid="7453" lane="3" entrytime="00:02:04.00" />
                <RESULT eventid="1673" points="130" reactiontime="+95" swimtime="00:00:56.33" resultid="4094" heatid="7538" lane="7" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="4068">
              <RESULTS>
                <RESULT eventid="1256" points="202" reactiontime="+90" swimtime="00:03:24.46" resultid="4069" heatid="7335" lane="1" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="240" reactiontime="+86" swimtime="00:01:29.48" resultid="4070" heatid="7419" lane="8" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="240" reactiontime="+92" swimtime="00:00:40.60" resultid="4071" heatid="7551" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="4081">
              <RESULTS>
                <RESULT eventid="1092" points="134" swimtime="00:03:58.02" resultid="4082" heatid="7272" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                    <SPLIT distance="100" swimtime="00:01:56.74" />
                    <SPLIT distance="150" swimtime="00:03:03.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="142" swimtime="00:04:17.35" resultid="4083" heatid="7328" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.86" />
                    <SPLIT distance="100" swimtime="00:02:02.63" />
                    <SPLIT distance="150" swimtime="00:03:10.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="136" swimtime="00:01:49.62" resultid="4084" heatid="7370" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="141" reactiontime="+93" swimtime="00:01:59.68" resultid="4085" heatid="7409" lane="6" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="99" swimtime="00:00:52.66" resultid="4086" heatid="7427" lane="6" entrytime="00:00:51.01" />
                <RESULT eventid="1608" points="95" reactiontime="+93" swimtime="00:01:59.53" resultid="4087" heatid="7508" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="Mazurek" nation="POL" athleteid="4113">
              <RESULTS>
                <RESULT eventid="1059" points="167" swimtime="00:00:41.56" resultid="4114" heatid="7238" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1304" points="154" reactiontime="+98" swimtime="00:01:45.31" resultid="4115" heatid="7371" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="175" swimtime="00:01:51.47" resultid="4116" heatid="7411" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="131" reactiontime="+95" swimtime="00:00:47.89" resultid="4117" heatid="7428" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1608" points="118" reactiontime="+94" swimtime="00:01:51.07" resultid="4118" heatid="7508" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="197" reactiontime="+98" swimtime="00:00:49.05" resultid="4119" heatid="7542" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="4107">
              <RESULTS>
                <RESULT eventid="1188" points="97" swimtime="00:30:41.46" resultid="4108" heatid="7304" lane="0" entrytime="00:29:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:51.87" />
                    <SPLIT distance="150" swimtime="00:02:53.73" />
                    <SPLIT distance="200" swimtime="00:03:57.07" />
                    <SPLIT distance="250" swimtime="00:05:00.70" />
                    <SPLIT distance="300" swimtime="00:06:03.77" />
                    <SPLIT distance="350" swimtime="00:07:07.45" />
                    <SPLIT distance="400" swimtime="00:08:11.58" />
                    <SPLIT distance="450" swimtime="00:09:14.65" />
                    <SPLIT distance="500" swimtime="00:10:17.15" />
                    <SPLIT distance="550" swimtime="00:11:20.09" />
                    <SPLIT distance="600" swimtime="00:12:22.27" />
                    <SPLIT distance="650" swimtime="00:13:25.01" />
                    <SPLIT distance="700" swimtime="00:14:27.71" />
                    <SPLIT distance="750" swimtime="00:15:29.97" />
                    <SPLIT distance="800" swimtime="00:16:31.83" />
                    <SPLIT distance="850" swimtime="00:17:32.87" />
                    <SPLIT distance="900" swimtime="00:18:34.07" />
                    <SPLIT distance="950" swimtime="00:19:35.35" />
                    <SPLIT distance="1000" swimtime="00:20:36.76" />
                    <SPLIT distance="1050" swimtime="00:21:38.51" />
                    <SPLIT distance="1100" swimtime="00:22:39.19" />
                    <SPLIT distance="1150" swimtime="00:23:39.64" />
                    <SPLIT distance="1200" swimtime="00:24:40.86" />
                    <SPLIT distance="1250" swimtime="00:25:42.02" />
                    <SPLIT distance="1300" swimtime="00:26:42.47" />
                    <SPLIT distance="1350" swimtime="00:27:44.26" />
                    <SPLIT distance="1400" swimtime="00:28:45.10" />
                    <SPLIT distance="1450" swimtime="00:29:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="35" swimtime="00:05:30.51" resultid="4109" heatid="7395" lane="7" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.01" />
                    <SPLIT distance="100" swimtime="00:02:29.86" />
                    <SPLIT distance="150" swimtime="00:04:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="4110" heatid="8154" lane="3" entrytime="00:08:40.00" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="4111" heatid="7513" lane="6" entrytime="00:02:15.00" />
                <RESULT eventid="1689" points="147" swimtime="00:00:47.83" resultid="4112" heatid="7549" lane="3" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="4056">
              <RESULTS>
                <RESULT eventid="1059" points="211" swimtime="00:00:38.50" resultid="4057" heatid="7237" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1207" points="161" reactiontime="+85" swimtime="00:00:47.11" resultid="4058" heatid="7309" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1272" points="186" reactiontime="+97" swimtime="00:01:27.89" resultid="4059" heatid="7342" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="132" reactiontime="+82" swimtime="00:01:47.93" resultid="4060" heatid="7454" lane="8" entrytime="00:01:44.00" />
                <RESULT eventid="1497" points="147" swimtime="00:03:29.16" resultid="4061" heatid="7469" lane="5" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:38.78" />
                    <SPLIT distance="150" swimtime="00:02:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="132" reactiontime="+90" swimtime="00:03:54.01" resultid="4062" heatid="7525" lane="6" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.16" />
                    <SPLIT distance="100" swimtime="00:01:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="4063" heatid="7570" lane="2" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="Radkowiak" nation="POL" athleteid="4072">
              <RESULTS>
                <RESULT eventid="1059" points="194" swimtime="00:00:39.60" resultid="4073" heatid="7237" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1092" points="120" swimtime="00:04:06.66" resultid="4074" heatid="7272" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                    <SPLIT distance="100" swimtime="00:02:02.27" />
                    <SPLIT distance="150" swimtime="00:03:09.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="95" reactiontime="+96" swimtime="00:00:56.19" resultid="4075" heatid="7308" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="4076" heatid="7328" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1400" points="159" reactiontime="+96" swimtime="00:01:54.87" resultid="4077" heatid="7409" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="112" reactiontime="+98" swimtime="00:08:56.79" resultid="4078" heatid="8149" lane="6" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.50" />
                    <SPLIT distance="100" swimtime="00:02:02.16" />
                    <SPLIT distance="150" swimtime="00:03:18.34" />
                    <SPLIT distance="200" swimtime="00:04:31.04" />
                    <SPLIT distance="250" swimtime="00:05:43.18" />
                    <SPLIT distance="300" swimtime="00:06:56.07" />
                    <SPLIT distance="350" swimtime="00:07:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="4079" heatid="7508" lane="8" entrytime="00:02:00.00" />
                <RESULT eventid="1673" points="175" reactiontime="+93" swimtime="00:00:50.99" resultid="4080" heatid="7538" lane="4" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="4098">
              <RESULTS>
                <RESULT eventid="1076" points="72" swimtime="00:00:48.60" resultid="4099" heatid="7249" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1108" points="61" reactiontime="+80" swimtime="00:04:38.01" resultid="4100" heatid="7277" lane="4" entrytime="00:04:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.34" />
                    <SPLIT distance="100" swimtime="00:02:23.51" />
                    <SPLIT distance="150" swimtime="00:03:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="85" swimtime="00:04:32.73" resultid="4101" heatid="7333" lane="7" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.46" />
                    <SPLIT distance="100" swimtime="00:02:12.18" />
                    <SPLIT distance="150" swimtime="00:03:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="63" swimtime="00:02:06.07" resultid="4102" heatid="7378" lane="7" entrytime="00:01:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="95" reactiontime="+96" swimtime="00:02:01.66" resultid="4103" heatid="7416" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="39" reactiontime="+89" swimtime="00:02:23.65" resultid="4104" heatid="7460" lane="4" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="39" reactiontime="+91" swimtime="00:05:09.89" resultid="4105" heatid="7530" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:30.71" />
                    <SPLIT distance="150" swimtime="00:03:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="127" reactiontime="+98" swimtime="00:00:50.12" resultid="4106" heatid="7548" lane="1" entrytime="00:00:51.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Anna" gender="F" lastname="Walczak" nation="POL" athleteid="4095">
              <RESULTS>
                <RESULT eventid="1059" points="88" swimtime="00:00:51.54" resultid="4096" heatid="7235" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1207" points="105" reactiontime="+53" swimtime="00:00:54.31" resultid="4097" heatid="7308" lane="0" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="110" swimtime="00:02:50.28" resultid="4135" heatid="7493" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                    <SPLIT distance="100" swimtime="00:01:26.78" />
                    <SPLIT distance="150" swimtime="00:02:15.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4107" number="1" />
                    <RELAYPOSITION athleteid="4064" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4098" number="3" reactiontime="+96" />
                    <RELAYPOSITION athleteid="4068" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S1 - Pływak utraciły kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 13:47)" eventid="1391" reactiontime="+94" status="DSQ" swimtime="00:03:18.16" resultid="4136" heatid="7403" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="100" swimtime="00:01:37.55" />
                    <SPLIT distance="150" swimtime="00:02:40.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4098" number="1" reactiontime="+94" status="DSQ" />
                    <RELAYPOSITION athleteid="4068" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="4107" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="4064" number="4" reactiontime="-13" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="175" swimtime="00:02:47.76" resultid="4140" heatid="7490" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:26.39" />
                    <SPLIT distance="150" swimtime="00:02:06.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4081" number="1" />
                    <RELAYPOSITION athleteid="4113" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4072" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="4056" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="155" reactiontime="+88" swimtime="00:03:10.55" resultid="4141" heatid="7400" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.29" />
                    <SPLIT distance="150" swimtime="00:02:27.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4056" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="4072" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4113" number="3" />
                    <RELAYPOSITION athleteid="4081" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" status="WDR" swimtime="00:00:00.00" resultid="4142" heatid="7399" lane="5" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4095" number="1" />
                    <RELAYPOSITION athleteid="4120" number="2" />
                    <RELAYPOSITION athleteid="4129" number="3" />
                    <RELAYPOSITION athleteid="4088" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="4143" heatid="7490" lane="9" entrytime="00:03:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4095" number="1" />
                    <RELAYPOSITION athleteid="4120" number="2" />
                    <RELAYPOSITION athleteid="4129" number="3" />
                    <RELAYPOSITION athleteid="4088" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="125" reactiontime="+74" swimtime="00:03:12.41" resultid="4134" heatid="7563" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                    <SPLIT distance="150" swimtime="00:02:23.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4095" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4068" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4113" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4098" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1124" points="140" swimtime="00:02:48.94" resultid="4137" heatid="7287" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:29.41" />
                    <SPLIT distance="150" swimtime="00:02:14.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4081" number="1" />
                    <RELAYPOSITION athleteid="4098" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4120" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4068" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="142" reactiontime="+86" swimtime="00:03:04.57" resultid="4138" heatid="7562" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                    <SPLIT distance="100" swimtime="00:01:35.84" />
                    <SPLIT distance="150" swimtime="00:02:26.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4056" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="4107" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4072" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4064" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="148" reactiontime="+97" swimtime="00:02:46.01" resultid="4139" heatid="7287" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:08.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4072" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="4107" number="2" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4113" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4064" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="GWWRO" nation="POL" region="01" clubid="6415" name="Grupa Wodna Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1980-09-05" firstname="Tomasz" gender="M" lastname="Spychalski " nation="POL" athleteid="6414">
              <RESULTS>
                <RESULT eventid="1188" points="303" swimtime="00:21:01.66" resultid="6416" heatid="7302" lane="0" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                    <SPLIT distance="200" swimtime="00:02:27.42" />
                    <SPLIT distance="250" swimtime="00:03:08.15" />
                    <SPLIT distance="300" swimtime="00:03:49.80" />
                    <SPLIT distance="350" swimtime="00:04:31.97" />
                    <SPLIT distance="400" swimtime="00:05:14.33" />
                    <SPLIT distance="450" swimtime="00:05:56.57" />
                    <SPLIT distance="500" swimtime="00:06:39.39" />
                    <SPLIT distance="550" swimtime="00:07:22.35" />
                    <SPLIT distance="600" swimtime="00:08:05.86" />
                    <SPLIT distance="650" swimtime="00:08:49.53" />
                    <SPLIT distance="700" swimtime="00:09:33.24" />
                    <SPLIT distance="750" swimtime="00:10:17.26" />
                    <SPLIT distance="800" swimtime="00:11:01.12" />
                    <SPLIT distance="850" swimtime="00:11:45.04" />
                    <SPLIT distance="900" swimtime="00:12:28.65" />
                    <SPLIT distance="950" swimtime="00:13:11.93" />
                    <SPLIT distance="1000" swimtime="00:13:54.94" />
                    <SPLIT distance="1050" swimtime="00:14:38.67" />
                    <SPLIT distance="1100" swimtime="00:15:21.65" />
                    <SPLIT distance="1150" swimtime="00:16:05.33" />
                    <SPLIT distance="1200" swimtime="00:16:48.24" />
                    <SPLIT distance="1250" swimtime="00:17:32.00" />
                    <SPLIT distance="1300" swimtime="00:18:14.92" />
                    <SPLIT distance="1350" swimtime="00:18:57.31" />
                    <SPLIT distance="1400" swimtime="00:19:40.28" />
                    <SPLIT distance="1450" swimtime="00:20:22.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="IKKON" nation="POL" region="14" clubid="5187" name="IKS Konstancin">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1999-09-11" firstname="Maciej" gender="M" lastname="Pecyna" nation="POL" athleteid="5188">
              <RESULTS>
                <RESULT eventid="1288" points="625" reactiontime="+77" swimtime="00:00:52.55" resultid="5189" heatid="7366" lane="8" entrytime="00:00:56.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="574" reactiontime="+75" swimtime="00:00:26.17" resultid="5190" heatid="7450" lane="3" entrytime="00:00:26.10" />
                <RESULT eventid="1513" points="588" reactiontime="+77" swimtime="00:01:58.59" resultid="5191" heatid="7488" lane="8" entrytime="00:02:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:58.99" />
                    <SPLIT distance="150" swimtime="00:01:29.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ILKAI" nation="LTU" clubid="5752" name="Ilgaplaukiai Kaisiadorys">
          <ATHLETES>
            <ATHLETE birthdate="1966-11-04" firstname="Vaidotas" gender="M" lastname="Gumbis" nation="LTU" athleteid="5751">
              <RESULTS>
                <RESULT eventid="1076" points="405" reactiontime="+94" swimtime="00:00:27.38" resultid="5753" heatid="7264" lane="9" entrytime="00:00:27.13" />
                <RESULT eventid="1288" points="423" reactiontime="+73" swimtime="00:00:59.85" resultid="5754" heatid="7362" lane="2" entrytime="00:01:00.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="400" reactiontime="+67" swimtime="00:02:14.76" resultid="5755" heatid="7483" lane="5" entrytime="00:02:18.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:04.66" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="5756" heatid="7584" lane="3" entrytime="00:04:53.03" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ISBIA" nation="POL" region="09" clubid="6339" name="Iswim Białystok">
          <CONTACT email="biuro@isiwm.bialystok.pl" internet="www.iswim.bialystok.pl" name="SEBSTAIN HUMBLA" phone="782997050" street="WIERZBOWA 3" street2="Białystok" />
          <ATHLETES>
            <ATHLETE birthdate="1979-11-12" firstname="Piotr" gender="M" lastname="Buczko" nation="POL" athleteid="6340">
              <RESULTS>
                <RESULT eventid="1076" points="449" reactiontime="+78" swimtime="00:00:26.45" resultid="6341" heatid="7263" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6342" heatid="7445" lane="4" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-12" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="6343">
              <RESULTS>
                <RESULT eventid="1076" points="423" reactiontime="+76" swimtime="00:00:26.97" resultid="6344" heatid="7261" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1224" points="340" reactiontime="+72" swimtime="00:00:31.83" resultid="6345" heatid="7324" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1320" points="305" reactiontime="+72" swimtime="00:01:14.59" resultid="6346" heatid="7385" lane="1" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="431" reactiontime="+70" swimtime="00:00:28.78" resultid="6347" heatid="7446" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1689" points="451" reactiontime="+70" swimtime="00:00:32.92" resultid="6348" heatid="7559" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-01" firstname="Justyna" gender="F" lastname="Hermanowicz" nation="POL" athleteid="6389">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="6390" heatid="7241" lane="7" entrytime="00:00:32.90" />
                <RESULT eventid="1272" points="317" reactiontime="+97" swimtime="00:01:13.67" resultid="6391" heatid="7346" lane="3" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="290" reactiontime="+96" swimtime="00:02:46.71" resultid="6392" heatid="7474" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:02:00.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="6393" heatid="7567" lane="5" entrytime="00:05:19.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-24" firstname="Sebastian" gender="M" lastname="Humbla" nation="POL" athleteid="6370">
              <RESULTS>
                <RESULT eventid="1076" points="506" reactiontime="+76" swimtime="00:00:25.42" resultid="6371" heatid="7266" lane="9" entrytime="00:00:26.60" />
                <RESULT eventid="1224" points="379" reactiontime="+70" swimtime="00:00:30.70" resultid="6372" heatid="7324" lane="4" entrytime="00:00:31.38" />
                <RESULT eventid="1320" points="474" reactiontime="+71" swimtime="00:01:04.44" resultid="6373" heatid="7388" lane="8" entrytime="00:01:06.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="477" reactiontime="+74" swimtime="00:00:27.82" resultid="6374" heatid="7448" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1689" points="478" reactiontime="+70" swimtime="00:00:32.28" resultid="6375" heatid="7559" lane="5" entrytime="00:00:33.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-17" firstname="Magdalena" gender="F" lastname="Iwaniuk Mróz" nation="POL" athleteid="6400">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="6410" heatid="7242" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="6411" heatid="7347" lane="7" entrytime="00:01:06.00" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="6412" heatid="7373" lane="2" entrytime="00:01:22.90" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="6413" heatid="7430" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-12" firstname="Piotr" gender="M" lastname="Iłendo" nation="POL" athleteid="6349">
              <RESULTS>
                <RESULT eventid="1076" points="527" reactiontime="+68" swimtime="00:00:25.08" resultid="6350" heatid="7268" lane="4" entrytime="00:00:25.20" />
                <RESULT eventid="1288" points="552" reactiontime="+71" swimtime="00:00:54.77" resultid="6351" heatid="7366" lane="1" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="540" reactiontime="+64" swimtime="00:02:01.97" resultid="6352" heatid="7487" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                    <SPLIT distance="100" swimtime="00:00:58.53" />
                    <SPLIT distance="150" swimtime="00:01:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="436" reactiontime="+71" swimtime="00:02:19.27" resultid="6353" heatid="7536" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="150" swimtime="00:01:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-21" firstname="Ewa" gender="F" lastname="Markowska" nation="POL" athleteid="6354">
              <RESULTS>
                <RESULT eventid="1140" points="152" reactiontime="+95" swimtime="00:14:57.92" resultid="6355" heatid="7292" lane="2" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                    <SPLIT distance="100" swimtime="00:01:35.68" />
                    <SPLIT distance="150" swimtime="00:02:31.28" />
                    <SPLIT distance="200" swimtime="00:03:28.25" />
                    <SPLIT distance="250" swimtime="00:04:23.94" />
                    <SPLIT distance="300" swimtime="00:05:21.62" />
                    <SPLIT distance="350" swimtime="00:06:19.63" />
                    <SPLIT distance="400" swimtime="00:07:18.54" />
                    <SPLIT distance="450" swimtime="00:08:16.96" />
                    <SPLIT distance="500" swimtime="00:09:14.25" />
                    <SPLIT distance="550" swimtime="00:10:12.76" />
                    <SPLIT distance="600" swimtime="00:11:12.33" />
                    <SPLIT distance="650" swimtime="00:12:10.43" />
                    <SPLIT distance="700" swimtime="00:13:08.87" />
                    <SPLIT distance="750" swimtime="00:14:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="6356" heatid="7392" lane="2" entrytime="00:03:40.00" />
                <RESULT eventid="1561" points="153" swimtime="00:08:04.06" resultid="6357" heatid="8150" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.80" />
                    <SPLIT distance="100" swimtime="00:02:06.25" />
                    <SPLIT distance="150" swimtime="00:03:12.38" />
                    <SPLIT distance="200" swimtime="00:04:16.01" />
                    <SPLIT distance="250" swimtime="00:05:11.38" />
                    <SPLIT distance="300" swimtime="00:06:10.38" />
                    <SPLIT distance="350" swimtime="00:07:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="6358" heatid="7570" lane="5" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-10" firstname="Dawid" gender="M" lastname="Perkowski" nation="POL" athleteid="6359">
              <RESULTS>
                <RESULT eventid="1076" points="536" reactiontime="+65" swimtime="00:00:24.93" resultid="6360" heatid="7268" lane="5" entrytime="00:00:25.30" />
                <RESULT eventid="1352" points="475" reactiontime="+62" swimtime="00:02:18.70" resultid="6361" heatid="7398" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:03.72" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="557" reactiontime="+65" swimtime="00:00:26.43" resultid="6362" heatid="7451" lane="0" entrytime="00:00:25.90" />
                <RESULT eventid="1625" points="548" reactiontime="+66" swimtime="00:00:58.74" resultid="6363" heatid="7521" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-09-27" firstname="Józef" gender="M" lastname="Sawicki" nation="POL" athleteid="6364">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="6365" heatid="7265" lane="5" entrytime="00:00:26.99" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="6366" heatid="7297" lane="0" entrytime="00:12:30.00" />
                <RESULT eventid="1288" points="443" reactiontime="+67" swimtime="00:00:58.95" resultid="6367" heatid="7363" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu. (Time: 19:26)" eventid="1513" reactiontime="+52" status="DSQ" swimtime="00:02:13.97" resultid="6368" heatid="7485" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:05.29" />
                    <SPLIT distance="150" swimtime="00:01:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="370" reactiontime="+77" swimtime="00:04:55.61" resultid="6369" heatid="7576" lane="3" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:46.66" />
                    <SPLIT distance="250" swimtime="00:03:03.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Agnieszka" gender="F" lastname="Stefanowska" nation="POL" athleteid="6394">
              <RESULTS>
                <RESULT eventid="1172" points="212" swimtime="00:25:41.67" resultid="6395" heatid="7300" lane="0" entrytime="00:26:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="150" swimtime="00:02:23.34" />
                    <SPLIT distance="200" swimtime="00:03:14.51" />
                    <SPLIT distance="250" swimtime="00:04:05.93" />
                    <SPLIT distance="300" swimtime="00:04:57.48" />
                    <SPLIT distance="350" swimtime="00:05:49.62" />
                    <SPLIT distance="400" swimtime="00:06:41.23" />
                    <SPLIT distance="450" swimtime="00:07:32.87" />
                    <SPLIT distance="500" swimtime="00:08:24.20" />
                    <SPLIT distance="550" swimtime="00:09:16.71" />
                    <SPLIT distance="600" swimtime="00:10:09.04" />
                    <SPLIT distance="650" swimtime="00:11:00.42" />
                    <SPLIT distance="700" swimtime="00:11:52.97" />
                    <SPLIT distance="750" swimtime="00:12:45.88" />
                    <SPLIT distance="800" swimtime="00:13:37.11" />
                    <SPLIT distance="850" swimtime="00:14:28.91" />
                    <SPLIT distance="900" swimtime="00:15:21.00" />
                    <SPLIT distance="950" swimtime="00:16:12.95" />
                    <SPLIT distance="1000" swimtime="00:17:04.89" />
                    <SPLIT distance="1050" swimtime="00:17:57.46" />
                    <SPLIT distance="1100" swimtime="00:18:50.54" />
                    <SPLIT distance="1150" swimtime="00:19:42.33" />
                    <SPLIT distance="1200" swimtime="00:20:34.06" />
                    <SPLIT distance="1250" swimtime="00:21:26.13" />
                    <SPLIT distance="1300" swimtime="00:22:17.59" />
                    <SPLIT distance="1350" swimtime="00:23:09.61" />
                    <SPLIT distance="1400" swimtime="00:24:00.96" />
                    <SPLIT distance="1450" swimtime="00:24:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="126" reactiontime="+93" swimtime="00:03:58.02" resultid="6396" heatid="7392" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                    <SPLIT distance="100" swimtime="00:01:46.89" />
                    <SPLIT distance="150" swimtime="00:02:51.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="169" swimtime="00:00:44.07" resultid="6397" heatid="7429" lane="0" entrytime="00:00:39.90" />
                <RESULT eventid="1608" points="159" reactiontime="+99" swimtime="00:01:40.79" resultid="6398" heatid="7509" lane="9" entrytime="00:01:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="6399" heatid="7570" lane="4" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-16" firstname="Karol" gender="M" lastname="Traciecki" nation="POL" athleteid="6385">
              <RESULTS>
                <RESULT eventid="1320" points="297" reactiontime="+74" swimtime="00:01:15.32" resultid="6386" heatid="7383" lane="4" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="308" reactiontime="+66" swimtime="00:01:22.29" resultid="6387" heatid="7422" lane="5" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="309" reactiontime="+72" swimtime="00:00:37.31" resultid="6388" heatid="7556" lane="2" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-17" firstname="Filip" gender="M" lastname="Walczuk" nation="POL" athleteid="6376">
              <RESULTS>
                <RESULT eventid="1076" points="427" reactiontime="+93" swimtime="00:00:26.89" resultid="6377" heatid="7264" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="6378" heatid="7359" lane="9" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-13" firstname="Dawid" gender="M" lastname="Świderski" nation="POL" athleteid="6379">
              <RESULTS>
                <RESULT eventid="1076" points="477" reactiontime="+73" swimtime="00:00:25.92" resultid="6380" heatid="7267" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="6381" heatid="7388" lane="0" entrytime="00:01:07.00" />
                <RESULT eventid="1352" points="410" reactiontime="+81" swimtime="00:02:25.65" resultid="6382" heatid="7395" lane="4" entrytime="00:03:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:47.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="483" reactiontime="+74" swimtime="00:00:27.72" resultid="6383" heatid="7448" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1625" points="478" reactiontime="+76" swimtime="00:01:01.49" resultid="6384" heatid="7520" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kategoria C" eventid="1545" points="500" reactiontime="+78" swimtime="00:01:43.00" resultid="6408" heatid="7496" lane="8" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.83" />
                    <SPLIT distance="100" swimtime="00:00:52.40" />
                    <SPLIT distance="150" swimtime="00:01:17.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6379" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="6376" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6370" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="6340" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="420" reactiontime="+85" swimtime="00:02:00.72" resultid="6875" heatid="7406" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:03.82" />
                    <SPLIT distance="150" swimtime="00:01:33.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6340" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="6370" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="6379" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="6376" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utraciły kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 20:10)" eventid="1545" reactiontime="+75" status="DSQ" swimtime="00:01:47.83" resultid="6405" heatid="7495" lane="4" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="100" swimtime="00:00:53.95" />
                    <SPLIT distance="150" swimtime="00:01:23.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6343" number="1" reactiontime="+75" status="DSQ" />
                    <RELAYPOSITION athleteid="6364" number="2" reactiontime="-19" status="DSQ" />
                    <RELAYPOSITION athleteid="6385" number="3" reactiontime="+46" status="DSQ" />
                    <RELAYPOSITION athleteid="6349" number="4" reactiontime="-3" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" status="DNS" swimtime="00:00:00.00" resultid="6876" heatid="7405" lane="4" entrytime="00:01:57.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6349" number="1" />
                    <RELAYPOSITION athleteid="6385" number="2" />
                    <RELAYPOSITION athleteid="6343" number="3" />
                    <RELAYPOSITION athleteid="6364" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="240" reactiontime="+86" swimtime="00:02:44.72" resultid="6406" heatid="7401" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6400" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="6354" number="2" />
                    <RELAYPOSITION athleteid="6394" number="3" />
                    <RELAYPOSITION athleteid="6389" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S1 - Pływak utraciły kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 20:09)" eventid="1529" reactiontime="+85" status="DSQ" swimtime="00:02:15.22" resultid="6407" heatid="7491" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:43.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6400" number="1" reactiontime="+85" status="DSQ" />
                    <RELAYPOSITION athleteid="6394" number="2" reactiontime="+53" status="DSQ" />
                    <RELAYPOSITION athleteid="6354" number="3" reactiontime="+58" status="DSQ" />
                    <RELAYPOSITION athleteid="6389" number="4" reactiontime="-87" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="6877" heatid="7289" lane="8" entrytime="00:01:58.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6340" number="1" />
                    <RELAYPOSITION athleteid="6400" number="2" />
                    <RELAYPOSITION athleteid="6389" number="3" />
                    <RELAYPOSITION athleteid="6376" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="329" reactiontime="+70" swimtime="00:02:19.64" resultid="6878" heatid="7565" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6349" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="6354" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="6364" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="6389" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="315" reactiontime="+72" swimtime="00:02:09.12" resultid="6409" heatid="7288" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="100" swimtime="00:01:03.64" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6343" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="6354" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="6394" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="6385" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="325" reactiontime="+77" swimtime="00:02:20.09" resultid="6879" heatid="7565" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6376" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="6343" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="6400" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="6394" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="JKKRA" nation="POL" region="06" clubid="2654" name="JK Team Kraków">
          <CONTACT name="Joanna Kwatera" phone="790611187" />
          <ATHLETES>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="2655">
              <RESULTS>
                <RESULT eventid="1240" points="291" reactiontime="+74" swimtime="00:03:22.93" resultid="2656" heatid="7330" lane="5" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:02:28.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="K3LVI" nation="UKR" clubid="4035" name="K3 Swim Lviv">
          <CONTACT city="Lviv" email="valentunakvita28@gmail.com" name="Kvita Valentyna" phone="+38 093 679 8731" />
          <ATHLETES>
            <ATHLETE birthdate="1988-06-28" firstname="Valentyna" gender="F" lastname="Kvita" nation="UKR" athleteid="4036">
              <RESULTS>
                <RESULT eventid="1059" points="552" reactiontime="+78" swimtime="00:00:27.94" resultid="4037" heatid="7244" lane="3" entrytime="00:00:28.80" />
                <RESULT eventid="1092" points="500" reactiontime="+84" swimtime="00:02:33.49" resultid="4038" heatid="7275" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:57.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="593" reactiontime="+77" swimtime="00:00:59.81" resultid="4039" heatid="7348" lane="9" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="523" reactiontime="+79" swimtime="00:01:10.10" resultid="4040" heatid="7375" lane="4" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="458" reactiontime="+81" swimtime="00:01:20.85" resultid="4041" heatid="7413" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="542" reactiontime="+83" swimtime="00:02:15.44" resultid="4042" heatid="7474" lane="9" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="150" swimtime="00:01:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="499" reactiontime="+70" swimtime="00:00:36.00" resultid="4043" heatid="7544" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1721" points="467" reactiontime="+79" swimtime="00:05:01.35" resultid="4044" heatid="7566" lane="8" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:46.66" />
                    <SPLIT distance="200" swimtime="00:02:25.03" />
                    <SPLIT distance="250" swimtime="00:03:04.18" />
                    <SPLIT distance="300" swimtime="00:03:43.42" />
                    <SPLIT distance="350" swimtime="00:04:22.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KATAK" nation="LTU" clubid="4220" name="Kauno Takas">
          <CONTACT city="Kaunas" internet="klubastakas.lt" name="Ramune Ivanauskaite" />
          <ATHLETES>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="Ivanauskaite" nation="LTU" athleteid="4221">
              <RESULTS>
                <RESULT eventid="1092" points="257" reactiontime="+94" swimtime="00:03:11.43" resultid="4222" heatid="7273" lane="1" entrytime="00:03:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:33.72" />
                    <SPLIT distance="150" swimtime="00:02:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="234" reactiontime="+100" swimtime="00:00:41.65" resultid="4223" heatid="7310" lane="7" entrytime="00:00:42.70" />
                <RESULT eventid="1240" points="295" swimtime="00:03:22.15" resultid="4224" heatid="7330" lane="0" entrytime="00:03:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="100" swimtime="00:01:38.07" />
                    <SPLIT distance="150" swimtime="00:02:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="270" reactiontime="+82" swimtime="00:01:36.38" resultid="4225" heatid="7410" lane="6" entrytime="00:01:43.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="242" reactiontime="+98" swimtime="00:01:28.19" resultid="4226" heatid="7455" lane="1" entrytime="00:01:33.20" />
                <RESULT eventid="1641" points="271" swimtime="00:03:04.16" resultid="4227" heatid="7526" lane="1" entrytime="00:03:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="150" swimtime="00:02:17.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-05-07" firstname="Jolanta" gender="F" lastname="Kozak" nation="LTU" athleteid="4228">
              <RESULTS>
                <RESULT eventid="1140" points="83" swimtime="00:18:15.23" resultid="4229" heatid="7292" lane="9" entrytime="00:17:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.56" />
                    <SPLIT distance="100" swimtime="00:02:14.23" />
                    <SPLIT distance="150" swimtime="00:03:28.73" />
                    <SPLIT distance="200" swimtime="00:04:42.71" />
                    <SPLIT distance="250" swimtime="00:05:56.97" />
                    <SPLIT distance="300" swimtime="00:07:11.63" />
                    <SPLIT distance="350" swimtime="00:08:27.15" />
                    <SPLIT distance="400" swimtime="00:09:42.12" />
                    <SPLIT distance="450" swimtime="00:10:56.24" />
                    <SPLIT distance="500" swimtime="00:12:09.59" />
                    <SPLIT distance="550" swimtime="00:13:24.94" />
                    <SPLIT distance="600" swimtime="00:14:38.67" />
                    <SPLIT distance="650" swimtime="00:15:53.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="67" reactiontime="+81" swimtime="00:01:03.01" resultid="4230" heatid="7308" lane="9" entrytime="00:00:59.50" />
                <RESULT eventid="1272" points="67" swimtime="00:02:03.17" resultid="4231" heatid="7341" lane="2" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="63" swimtime="00:04:37.48" resultid="4232" heatid="7468" lane="6" entrytime="00:04:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.07" />
                    <SPLIT distance="100" swimtime="00:02:14.12" />
                    <SPLIT distance="150" swimtime="00:03:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="4233" heatid="7571" lane="3" entrytime="00:08:21.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="Yliene" nation="LTU" athleteid="4234">
              <RESULTS>
                <RESULT eventid="1059" points="105" swimtime="00:00:48.49" resultid="4235" heatid="7236" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1207" points="104" reactiontime="+86" swimtime="00:00:54.44" resultid="4236" heatid="7309" lane="9" entrytime="00:00:53.00" />
                <RESULT eventid="1465" points="81" reactiontime="+93" swimtime="00:02:07.05" resultid="4237" heatid="7453" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="81" reactiontime="+91" swimtime="00:04:34.75" resultid="4238" heatid="7524" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.74" />
                    <SPLIT distance="100" swimtime="00:02:14.37" />
                    <SPLIT distance="150" swimtime="00:03:27.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00306" nation="POL" region="06" clubid="4764" name="Korona Masters  Kraków ">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="4765">
              <RESULTS>
                <RESULT eventid="1433" points="272" reactiontime="+98" swimtime="00:00:37.59" resultid="4766" heatid="7430" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1561" points="222" swimtime="00:07:07.33" resultid="4767" heatid="8150" lane="8" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                    <SPLIT distance="100" swimtime="00:01:40.66" />
                    <SPLIT distance="150" swimtime="00:02:36.98" />
                    <SPLIT distance="200" swimtime="00:03:33.69" />
                    <SPLIT distance="250" swimtime="00:04:32.77" />
                    <SPLIT distance="300" swimtime="00:05:32.26" />
                    <SPLIT distance="350" swimtime="00:06:21.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="198" reactiontime="+97" swimtime="00:01:33.55" resultid="4768" heatid="7509" lane="7" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="4842">
              <RESULTS>
                <RESULT eventid="1076" points="77" swimtime="00:00:47.47" resultid="4843" heatid="7248" lane="2" entrytime="00:00:47.00" />
                <RESULT eventid="1224" points="45" reactiontime="+76" swimtime="00:01:02.17" resultid="4844" heatid="7317" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1288" points="70" swimtime="00:01:48.63" resultid="4845" heatid="7350" lane="3" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="57" reactiontime="+99" swimtime="00:02:23.72" resultid="4846" heatid="7415" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="56" swimtime="00:04:19.44" resultid="4847" heatid="7475" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.34" />
                    <SPLIT distance="100" swimtime="00:01:55.59" />
                    <SPLIT distance="150" swimtime="00:03:09.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="51" reactiontime="+75" swimtime="00:04:43.35" resultid="4848" heatid="7530" lane="9" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.41" />
                    <SPLIT distance="100" swimtime="00:02:14.68" />
                    <SPLIT distance="150" swimtime="00:03:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="68" reactiontime="+97" swimtime="00:01:01.82" resultid="4849" heatid="7547" lane="6" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="4820">
              <RESULTS>
                <RESULT eventid="1059" points="266" swimtime="00:00:35.61" resultid="4821" heatid="7239" lane="8" entrytime="00:00:35.71" />
                <RESULT eventid="1092" points="190" swimtime="00:03:31.96" resultid="4822" heatid="7272" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:40.18" />
                    <SPLIT distance="150" swimtime="00:02:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="188" reactiontime="+91" swimtime="00:00:44.78" resultid="4823" heatid="7310" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1336" points="137" swimtime="00:03:51.58" resultid="4824" heatid="7392" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                    <SPLIT distance="100" swimtime="00:01:46.43" />
                    <SPLIT distance="150" swimtime="00:02:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="164" swimtime="00:00:44.47" resultid="4825" heatid="7428" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1561" points="163" swimtime="00:07:53.18" resultid="4826" heatid="8149" lane="4" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.35" />
                    <SPLIT distance="100" swimtime="00:01:53.48" />
                    <SPLIT distance="150" swimtime="00:02:55.84" />
                    <SPLIT distance="200" swimtime="00:03:57.99" />
                    <SPLIT distance="250" swimtime="00:04:21.98" />
                    <SPLIT distance="300" swimtime="00:05:02.18" />
                    <SPLIT distance="350" swimtime="00:06:04.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="137" swimtime="00:01:45.75" resultid="4827" heatid="7507" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="203" reactiontime="+96" swimtime="00:00:48.52" resultid="4828" heatid="7539" lane="8" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="4769">
              <RESULTS>
                <RESULT eventid="1059" points="305" swimtime="00:00:34.03" resultid="4770" heatid="7240" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1140" points="279" reactiontime="+94" swimtime="00:12:12.90" resultid="4771" heatid="7291" lane="7" entrytime="00:12:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:09.74" />
                    <SPLIT distance="200" swimtime="00:02:56.16" />
                    <SPLIT distance="250" swimtime="00:03:42.96" />
                    <SPLIT distance="300" swimtime="00:04:29.46" />
                    <SPLIT distance="350" swimtime="00:05:16.85" />
                    <SPLIT distance="400" swimtime="00:06:03.40" />
                    <SPLIT distance="450" swimtime="00:06:50.19" />
                    <SPLIT distance="500" swimtime="00:07:37.13" />
                    <SPLIT distance="550" swimtime="00:08:23.78" />
                    <SPLIT distance="600" swimtime="00:09:10.76" />
                    <SPLIT distance="650" swimtime="00:09:57.92" />
                    <SPLIT distance="700" swimtime="00:10:44.21" />
                    <SPLIT distance="750" swimtime="00:11:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="304" reactiontime="+91" swimtime="00:01:14.67" resultid="4772" heatid="7344" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="211" reactiontime="+93" swimtime="00:03:20.74" resultid="4773" heatid="7393" lane="9" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:33.20" />
                    <SPLIT distance="150" swimtime="00:02:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="301" reactiontime="+85" swimtime="00:02:44.71" resultid="4774" heatid="7471" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:03.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="250" swimtime="00:06:50.67" resultid="4775" heatid="8150" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:01:35.80" />
                    <SPLIT distance="150" swimtime="00:02:29.91" />
                    <SPLIT distance="200" swimtime="00:03:22.15" />
                    <SPLIT distance="250" swimtime="00:04:20.23" />
                    <SPLIT distance="300" swimtime="00:05:20.75" />
                    <SPLIT distance="350" swimtime="00:06:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="235" swimtime="00:01:28.43" resultid="4776" heatid="7509" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="286" reactiontime="+91" swimtime="00:05:54.87" resultid="4777" heatid="7568" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="150" swimtime="00:02:07.04" />
                    <SPLIT distance="200" swimtime="00:02:52.82" />
                    <SPLIT distance="250" swimtime="00:03:38.91" />
                    <SPLIT distance="300" swimtime="00:04:25.52" />
                    <SPLIT distance="350" swimtime="00:05:11.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="4778">
              <RESULTS>
                <RESULT eventid="1076" points="195" swimtime="00:00:34.93" resultid="4779" heatid="7253" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1156" points="113" swimtime="00:15:15.62" resultid="4780" heatid="7299" lane="3" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                    <SPLIT distance="100" swimtime="00:01:42.95" />
                    <SPLIT distance="150" swimtime="00:02:38.92" />
                    <SPLIT distance="200" swimtime="00:03:34.87" />
                    <SPLIT distance="250" swimtime="00:04:30.94" />
                    <SPLIT distance="300" swimtime="00:05:26.30" />
                    <SPLIT distance="350" swimtime="00:06:22.97" />
                    <SPLIT distance="400" swimtime="00:07:19.26" />
                    <SPLIT distance="450" swimtime="00:08:15.65" />
                    <SPLIT distance="500" swimtime="00:09:12.21" />
                    <SPLIT distance="550" swimtime="00:10:11.31" />
                    <SPLIT distance="600" swimtime="00:11:11.20" />
                    <SPLIT distance="650" swimtime="00:12:12.32" />
                    <SPLIT distance="700" swimtime="00:13:13.90" />
                    <SPLIT distance="750" swimtime="00:14:15.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="197" swimtime="00:01:17.21" resultid="4781" heatid="7354" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="49" swimtime="00:04:55.48" resultid="4782" heatid="7395" lane="8" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.51" />
                    <SPLIT distance="100" swimtime="00:02:22.29" />
                    <SPLIT distance="150" swimtime="00:03:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="128" swimtime="00:03:16.77" resultid="4783" heatid="7478" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:24.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNF" swimtime="00:00:00.00" resultid="4784" heatid="8154" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.92" />
                    <SPLIT distance="100" swimtime="00:02:19.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="73" swimtime="00:01:54.79" resultid="4785" heatid="7514" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="117" swimtime="00:07:13.85" resultid="4786" heatid="7582" lane="6" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                    <SPLIT distance="100" swimtime="00:01:41.10" />
                    <SPLIT distance="150" swimtime="00:02:35.58" />
                    <SPLIT distance="200" swimtime="00:03:30.64" />
                    <SPLIT distance="250" swimtime="00:04:26.85" />
                    <SPLIT distance="300" swimtime="00:05:23.27" />
                    <SPLIT distance="350" swimtime="00:06:18.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz-Musiał" nation="POL" athleteid="4787">
              <RESULTS>
                <RESULT eventid="1092" points="77" reactiontime="+99" swimtime="00:04:45.90" resultid="4788" heatid="7271" lane="1" entrytime="00:04:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.32" />
                    <SPLIT distance="100" swimtime="00:02:19.09" />
                    <SPLIT distance="150" swimtime="00:03:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="103" reactiontime="+96" swimtime="00:32:36.56" resultid="4789" heatid="7301" lane="2" entrytime="00:31:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                    <SPLIT distance="100" swimtime="00:01:51.00" />
                    <SPLIT distance="150" swimtime="00:02:54.69" />
                    <SPLIT distance="200" swimtime="00:03:59.96" />
                    <SPLIT distance="250" swimtime="00:05:06.53" />
                    <SPLIT distance="300" swimtime="00:06:11.66" />
                    <SPLIT distance="350" swimtime="00:07:18.16" />
                    <SPLIT distance="400" swimtime="00:08:21.94" />
                    <SPLIT distance="450" swimtime="00:09:26.12" />
                    <SPLIT distance="500" swimtime="00:10:32.79" />
                    <SPLIT distance="550" swimtime="00:11:37.93" />
                    <SPLIT distance="600" swimtime="00:12:43.36" />
                    <SPLIT distance="650" swimtime="00:13:48.21" />
                    <SPLIT distance="700" swimtime="00:14:52.88" />
                    <SPLIT distance="750" swimtime="00:15:59.40" />
                    <SPLIT distance="800" swimtime="00:17:03.73" />
                    <SPLIT distance="850" swimtime="00:18:08.10" />
                    <SPLIT distance="900" swimtime="00:19:13.33" />
                    <SPLIT distance="950" swimtime="00:20:18.83" />
                    <SPLIT distance="1000" swimtime="00:21:25.32" />
                    <SPLIT distance="1050" swimtime="00:22:32.58" />
                    <SPLIT distance="1100" swimtime="00:23:38.37" />
                    <SPLIT distance="1150" swimtime="00:24:43.70" />
                    <SPLIT distance="1200" swimtime="00:25:52.42" />
                    <SPLIT distance="1250" swimtime="00:27:00.83" />
                    <SPLIT distance="1300" swimtime="00:28:08.34" />
                    <SPLIT distance="1350" swimtime="00:29:14.76" />
                    <SPLIT distance="1400" swimtime="00:30:22.48" />
                    <SPLIT distance="1450" swimtime="00:31:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="81" reactiontime="+74" swimtime="00:00:59.21" resultid="4790" heatid="7307" lane="4" entrytime="00:01:01.00" />
                <RESULT eventid="1304" points="81" swimtime="00:02:10.50" resultid="4791" heatid="7369" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="82" reactiontime="+93" swimtime="00:02:23.49" resultid="4792" heatid="7408" lane="0" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="67" swimtime="00:01:00.01" resultid="4793" heatid="7426" lane="3" />
                <RESULT eventid="1608" points="59" reactiontime="+90" swimtime="00:02:20.13" resultid="4794" heatid="7507" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="99" reactiontime="+99" swimtime="00:08:24.85" resultid="4795" heatid="7571" lane="6" entrytime="00:08:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.81" />
                    <SPLIT distance="100" swimtime="00:01:54.64" />
                    <SPLIT distance="150" swimtime="00:02:59.47" />
                    <SPLIT distance="200" swimtime="00:04:04.70" />
                    <SPLIT distance="250" swimtime="00:05:09.58" />
                    <SPLIT distance="300" swimtime="00:06:15.60" />
                    <SPLIT distance="350" swimtime="00:07:21.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="4796">
              <RESULTS>
                <RESULT eventid="1076" points="324" reactiontime="+93" swimtime="00:00:29.48" resultid="4797" heatid="7257" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1224" points="267" reactiontime="+85" swimtime="00:00:34.49" resultid="4798" heatid="7322" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="326" reactiontime="+93" swimtime="00:01:13.01" resultid="4799" heatid="7383" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="351" reactiontime="+89" swimtime="00:00:30.83" resultid="4800" heatid="7443" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1481" points="282" reactiontime="+83" swimtime="00:01:14.50" resultid="4801" heatid="7464" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="313" reactiontime="+93" swimtime="00:01:10.79" resultid="4802" heatid="7519" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="343" reactiontime="+93" swimtime="00:00:36.07" resultid="4803" heatid="7555" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="4829">
              <RESULTS>
                <RESULT eventid="1076" points="185" reactiontime="+87" swimtime="00:00:35.52" resultid="4830" heatid="7249" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1224" points="84" reactiontime="+78" swimtime="00:00:50.56" resultid="4831" heatid="7318" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1320" points="98" reactiontime="+84" swimtime="00:01:48.81" resultid="4832" heatid="7378" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="78" reactiontime="+90" swimtime="00:01:54.07" resultid="4833" heatid="7461" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="104" reactiontime="+86" swimtime="00:00:53.60" resultid="4834" heatid="7546" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="4804">
              <RESULTS>
                <RESULT eventid="1076" points="260" reactiontime="+86" swimtime="00:00:31.74" resultid="4805" heatid="7256" lane="6" entrytime="00:00:31.19" />
                <RESULT eventid="1156" points="240" reactiontime="+72" swimtime="00:11:53.22" resultid="4806" heatid="7297" lane="8" entrytime="00:12:28.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:18.16" />
                    <SPLIT distance="150" swimtime="00:02:03.08" />
                    <SPLIT distance="200" swimtime="00:02:49.15" />
                    <SPLIT distance="250" swimtime="00:03:34.54" />
                    <SPLIT distance="300" swimtime="00:04:19.86" />
                    <SPLIT distance="350" swimtime="00:05:05.33" />
                    <SPLIT distance="400" swimtime="00:05:51.54" />
                    <SPLIT distance="450" swimtime="00:06:37.67" />
                    <SPLIT distance="500" swimtime="00:07:23.80" />
                    <SPLIT distance="550" swimtime="00:08:09.63" />
                    <SPLIT distance="600" swimtime="00:08:55.02" />
                    <SPLIT distance="650" swimtime="00:09:40.62" />
                    <SPLIT distance="700" swimtime="00:10:26.21" />
                    <SPLIT distance="750" swimtime="00:11:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="246" reactiontime="+97" swimtime="00:03:11.62" resultid="4807" heatid="7336" lane="7" entrytime="00:03:18.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:31.75" />
                    <SPLIT distance="150" swimtime="00:02:21.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="213" reactiontime="+83" swimtime="00:01:24.07" resultid="4808" heatid="7381" lane="7" entrytime="00:01:24.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="235" reactiontime="+87" swimtime="00:01:30.04" resultid="4809" heatid="7420" lane="8" entrytime="00:01:28.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="195" reactiontime="+71" swimtime="00:00:37.47" resultid="4810" heatid="7439" lane="0" entrytime="00:00:38.11" />
                <RESULT eventid="1689" points="295" reactiontime="+89" swimtime="00:00:37.92" resultid="4811" heatid="7554" lane="9" entrytime="00:00:38.88" />
                <RESULT eventid="1737" points="246" reactiontime="+97" swimtime="00:05:38.62" resultid="4812" heatid="7580" lane="5" entrytime="00:05:57.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:01:58.86" />
                    <SPLIT distance="200" swimtime="00:02:42.75" />
                    <SPLIT distance="250" swimtime="00:03:26.80" />
                    <SPLIT distance="300" swimtime="00:04:11.06" />
                    <SPLIT distance="350" swimtime="00:04:55.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-10-20" firstname="Janusz" gender="M" lastname="Toporski" nation="POL" athleteid="4835">
              <RESULTS>
                <RESULT eventid="1256" points="218" reactiontime="+84" swimtime="00:03:19.57" resultid="4836" heatid="7334" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                    <SPLIT distance="100" swimtime="00:01:37.54" />
                    <SPLIT distance="150" swimtime="00:02:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="121" reactiontime="+81" swimtime="00:03:38.40" resultid="4837" heatid="7395" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                    <SPLIT distance="100" swimtime="00:01:44.11" />
                    <SPLIT distance="150" swimtime="00:02:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="193" reactiontime="+89" swimtime="00:01:36.07" resultid="4838" heatid="7416" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="132" reactiontime="+88" swimtime="00:00:42.68" resultid="4839" heatid="7436" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1625" points="126" reactiontime="+80" swimtime="00:01:35.84" resultid="4840" heatid="7513" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="177" reactiontime="+74" swimtime="00:00:44.97" resultid="4841" heatid="7547" lane="2" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="4813">
              <RESULTS>
                <RESULT eventid="1076" points="73" swimtime="00:00:48.41" resultid="4814" heatid="7248" lane="7" entrytime="00:00:47.00" />
                <RESULT eventid="1188" points="69" swimtime="00:34:24.01" resultid="4815" heatid="7305" lane="5" entrytime="00:36:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.02" />
                    <SPLIT distance="100" swimtime="00:02:07.76" />
                    <SPLIT distance="150" swimtime="00:03:15.79" />
                    <SPLIT distance="200" swimtime="00:04:24.91" />
                    <SPLIT distance="250" swimtime="00:05:34.24" />
                    <SPLIT distance="300" swimtime="00:06:44.99" />
                    <SPLIT distance="350" swimtime="00:07:52.77" />
                    <SPLIT distance="400" swimtime="00:09:02.63" />
                    <SPLIT distance="450" swimtime="00:10:11.63" />
                    <SPLIT distance="500" swimtime="00:11:21.45" />
                    <SPLIT distance="550" swimtime="00:12:30.79" />
                    <SPLIT distance="600" swimtime="00:13:39.05" />
                    <SPLIT distance="650" swimtime="00:14:48.29" />
                    <SPLIT distance="700" swimtime="00:15:57.50" />
                    <SPLIT distance="750" swimtime="00:17:06.62" />
                    <SPLIT distance="800" swimtime="00:18:15.47" />
                    <SPLIT distance="850" swimtime="00:19:24.20" />
                    <SPLIT distance="900" swimtime="00:20:32.54" />
                    <SPLIT distance="950" swimtime="00:21:40.95" />
                    <SPLIT distance="1000" swimtime="00:22:50.74" />
                    <SPLIT distance="1050" swimtime="00:24:00.87" />
                    <SPLIT distance="1100" swimtime="00:25:10.20" />
                    <SPLIT distance="1150" swimtime="00:26:20.81" />
                    <SPLIT distance="1200" swimtime="00:27:31.32" />
                    <SPLIT distance="1250" swimtime="00:28:41.94" />
                    <SPLIT distance="1300" swimtime="00:29:52.41" />
                    <SPLIT distance="1350" swimtime="00:31:02.18" />
                    <SPLIT distance="1400" swimtime="00:32:11.77" />
                    <SPLIT distance="1450" swimtime="00:33:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="61" reactiontime="+96" swimtime="00:01:53.64" resultid="4816" heatid="7350" lane="4" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="60" swimtime="00:04:13.52" resultid="4817" heatid="7476" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="100" swimtime="00:02:02.00" />
                    <SPLIT distance="150" swimtime="00:03:09.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="51" swimtime="00:01:07.67" resultid="4818" heatid="7546" lane="4" entrytime="00:01:07.00" />
                <RESULT eventid="1737" points="58" swimtime="00:09:08.01" resultid="4819" heatid="7583" lane="0" entrytime="00:08:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.11" />
                    <SPLIT distance="100" swimtime="00:02:09.36" />
                    <SPLIT distance="150" swimtime="00:03:20.43" />
                    <SPLIT distance="200" swimtime="00:04:30.73" />
                    <SPLIT distance="250" swimtime="00:05:41.98" />
                    <SPLIT distance="300" swimtime="00:06:53.13" />
                    <SPLIT distance="350" swimtime="00:08:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="246" reactiontime="+91" swimtime="00:02:10.41" resultid="4852" heatid="7494" lane="9" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:41.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4804" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="4835" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4778" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4796" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="210" reactiontime="+75" swimtime="00:02:32.10" resultid="4853" heatid="7403" lane="4" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:01:57.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4796" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4835" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4804" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="4778" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="309" reactiontime="+87" swimtime="00:02:09.97" resultid="4850" heatid="7287" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4804" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="4769" number="2" />
                    <RELAYPOSITION athleteid="4820" number="3" reactiontime="-6" />
                    <RELAYPOSITION athleteid="4796" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="281" reactiontime="+76" swimtime="00:02:27.16" resultid="4851" heatid="7564" lane="9" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:01:50.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4769" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4804" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4796" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4820" number="4" reactiontime="+81" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="15" clubid="2094" name="KS Extreme Team Oborniki" shortname="Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANWOL@POCZTA.ONET.PL" name="WOLNIEWICZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="2095">
              <RESULTS>
                <RESULT eventid="1076" points="160" swimtime="00:00:37.28" resultid="2096" heatid="7252" lane="9" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1188" points="103" reactiontime="+99" swimtime="00:30:05.68" resultid="2097" heatid="7304" lane="9" entrytime="00:30:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                    <SPLIT distance="100" swimtime="00:01:45.95" />
                    <SPLIT distance="150" swimtime="00:02:44.18" />
                    <SPLIT distance="200" swimtime="00:03:44.07" />
                    <SPLIT distance="250" swimtime="00:04:43.34" />
                    <SPLIT distance="300" swimtime="00:05:42.93" />
                    <SPLIT distance="350" swimtime="00:06:41.78" />
                    <SPLIT distance="400" swimtime="00:07:41.63" />
                    <SPLIT distance="450" swimtime="00:08:41.13" />
                    <SPLIT distance="500" swimtime="00:09:41.22" />
                    <SPLIT distance="550" swimtime="00:10:41.54" />
                    <SPLIT distance="600" swimtime="00:11:41.44" />
                    <SPLIT distance="650" swimtime="00:12:41.47" />
                    <SPLIT distance="700" swimtime="00:13:41.76" />
                    <SPLIT distance="750" swimtime="00:14:43.27" />
                    <SPLIT distance="800" swimtime="00:15:44.05" />
                    <SPLIT distance="850" swimtime="00:16:44.91" />
                    <SPLIT distance="900" swimtime="00:17:46.55" />
                    <SPLIT distance="950" swimtime="00:18:48.01" />
                    <SPLIT distance="1000" swimtime="00:19:49.31" />
                    <SPLIT distance="1050" swimtime="00:20:51.64" />
                    <SPLIT distance="1100" swimtime="00:21:53.43" />
                    <SPLIT distance="1150" swimtime="00:22:55.09" />
                    <SPLIT distance="1200" swimtime="00:23:57.39" />
                    <SPLIT distance="1250" swimtime="00:24:58.63" />
                    <SPLIT distance="1300" swimtime="00:25:59.36" />
                    <SPLIT distance="1350" swimtime="00:27:01.66" />
                    <SPLIT distance="1400" swimtime="00:28:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="138" reactiontime="+98" swimtime="00:01:26.81" resultid="2098" heatid="7352" lane="6" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="102" reactiontime="+96" swimtime="00:03:32.44" resultid="2099" heatid="7477" lane="2" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:37.96" />
                    <SPLIT distance="150" swimtime="00:02:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="97" swimtime="00:07:41.14" resultid="2100" heatid="7582" lane="1" entrytime="00:07:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:41.68" />
                    <SPLIT distance="150" swimtime="00:02:41.18" />
                    <SPLIT distance="200" swimtime="00:03:41.03" />
                    <SPLIT distance="250" swimtime="00:04:41.60" />
                    <SPLIT distance="300" swimtime="00:05:42.12" />
                    <SPLIT distance="350" swimtime="00:06:44.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="3747" name="KS Górnik Radlin" shortname="Górnik Radlin">
          <ATHLETES>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="3748">
              <RESULTS>
                <RESULT eventid="1272" points="461" reactiontime="+86" swimtime="00:01:05.02" resultid="3749" heatid="7347" lane="0" entrytime="00:01:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="400" reactiontime="+92" swimtime="00:00:33.07" resultid="3750" heatid="7433" lane="0" entrytime="00:00:32.74" />
                <RESULT eventid="1608" points="357" reactiontime="+84" swimtime="00:01:16.92" resultid="3751" heatid="7510" lane="6" entrytime="00:01:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="390" reactiontime="+85" swimtime="00:00:39.08" resultid="3752" heatid="7544" lane="9" entrytime="00:00:38.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-22" firstname="Ryszard" gender="M" lastname="Kubica" nation="POL" license="100211700343" athleteid="3753">
              <RESULTS>
                <RESULT eventid="1076" points="359" reactiontime="+81" swimtime="00:00:28.48" resultid="3754" heatid="7259" lane="8" entrytime="00:00:29.43" />
                <RESULT eventid="1188" points="284" reactiontime="+97" swimtime="00:21:29.97" resultid="3755" heatid="7302" lane="1" entrytime="00:19:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                    <SPLIT distance="200" swimtime="00:02:34.65" />
                    <SPLIT distance="250" swimtime="00:03:16.47" />
                    <SPLIT distance="300" swimtime="00:03:58.18" />
                    <SPLIT distance="350" swimtime="00:04:40.27" />
                    <SPLIT distance="400" swimtime="00:05:23.21" />
                    <SPLIT distance="450" swimtime="00:06:06.46" />
                    <SPLIT distance="500" swimtime="00:06:49.87" />
                    <SPLIT distance="550" swimtime="00:07:33.55" />
                    <SPLIT distance="600" swimtime="00:08:17.30" />
                    <SPLIT distance="650" swimtime="00:09:01.07" />
                    <SPLIT distance="700" swimtime="00:09:45.06" />
                    <SPLIT distance="750" swimtime="00:10:29.21" />
                    <SPLIT distance="800" swimtime="00:11:12.94" />
                    <SPLIT distance="850" swimtime="00:11:56.50" />
                    <SPLIT distance="900" swimtime="00:12:40.71" />
                    <SPLIT distance="950" swimtime="00:13:24.77" />
                    <SPLIT distance="1000" swimtime="00:14:08.94" />
                    <SPLIT distance="1050" swimtime="00:14:53.03" />
                    <SPLIT distance="1100" swimtime="00:15:37.24" />
                    <SPLIT distance="1150" swimtime="00:16:21.51" />
                    <SPLIT distance="1200" swimtime="00:17:05.82" />
                    <SPLIT distance="1250" swimtime="00:17:49.93" />
                    <SPLIT distance="1300" swimtime="00:18:34.14" />
                    <SPLIT distance="1350" swimtime="00:19:18.76" />
                    <SPLIT distance="1400" swimtime="00:20:02.94" />
                    <SPLIT distance="1450" swimtime="00:20:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="239" reactiontime="+69" swimtime="00:00:35.79" resultid="3756" heatid="7321" lane="2" entrytime="00:00:36.88" />
                <RESULT eventid="1288" points="355" reactiontime="+81" swimtime="00:01:03.41" resultid="3757" heatid="7359" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="333" reactiontime="+81" swimtime="00:00:31.36" resultid="3758" heatid="7441" lane="4" entrytime="00:00:33.08" />
                <RESULT eventid="1513" points="303" reactiontime="+91" swimtime="00:02:27.86" resultid="3759" heatid="7482" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.58" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="271" reactiontime="+92" swimtime="00:01:14.27" resultid="3760" heatid="7517" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="284" reactiontime="+92" swimtime="00:05:22.55" resultid="3761" heatid="7578" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                    <SPLIT distance="200" swimtime="00:02:37.70" />
                    <SPLIT distance="250" swimtime="00:03:19.69" />
                    <SPLIT distance="300" swimtime="00:04:01.66" />
                    <SPLIT distance="350" swimtime="00:04:43.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKOWA" nation="POL" region="14" clubid="4281" name="KS Mako Warszawa" shortname="Mako Warszawa">
          <CONTACT city="Warszawa" email="ania.plywanie@gmail.com" name="Anna Dabrowska" phone="601480280" />
          <ATHLETES>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="4288">
              <RESULTS>
                <RESULT eventid="1076" points="154" reactiontime="+76" swimtime="00:00:37.74" resultid="4289" heatid="7250" lane="4" entrytime="00:00:38.02" />
                <RESULT eventid="1320" points="109" reactiontime="+72" swimtime="00:01:44.90" resultid="4290" heatid="7379" lane="9" entrytime="00:01:43.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="185" reactiontime="+75" swimtime="00:01:37.56" resultid="4291" heatid="7418" lane="0" entrytime="00:01:39.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="98" reactiontime="+74" swimtime="00:03:35.19" resultid="4292" heatid="7477" lane="9" entrytime="00:03:28.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="150" swimtime="00:02:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="212" reactiontime="+70" swimtime="00:00:42.33" resultid="4293" heatid="7551" lane="0" entrytime="00:00:42.02" />
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="4294" heatid="7584" lane="5" entrytime="00:07:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-12-14" firstname="Ada" gender="F" lastname="Andruszkiewicz" nation="POL" athleteid="4300">
              <RESULTS>
                <RESULT eventid="1272" points="254" reactiontime="+79" swimtime="00:01:19.30" resultid="4301" heatid="7343" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="214" reactiontime="+93" swimtime="00:01:34.37" resultid="4302" heatid="7368" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="220" reactiontime="+78" swimtime="00:01:31.13" resultid="4303" heatid="7454" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="217" reactiontime="+81" swimtime="00:03:18.20" resultid="4304" heatid="7523" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:38.29" />
                    <SPLIT distance="150" swimtime="00:02:29.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="4319">
              <RESULTS>
                <RESULT eventid="1092" points="298" reactiontime="+78" swimtime="00:03:02.42" resultid="4320" heatid="7272" lane="3" entrytime="00:03:20.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:02:19.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="298" reactiontime="+85" swimtime="00:11:57.00" resultid="4321" heatid="7291" lane="9" entrytime="00:13:07.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:08.24" />
                    <SPLIT distance="200" swimtime="00:02:53.26" />
                    <SPLIT distance="250" swimtime="00:03:37.24" />
                    <SPLIT distance="300" swimtime="00:04:22.18" />
                    <SPLIT distance="350" swimtime="00:05:07.33" />
                    <SPLIT distance="400" swimtime="00:05:52.33" />
                    <SPLIT distance="450" swimtime="00:06:37.32" />
                    <SPLIT distance="500" swimtime="00:07:23.19" />
                    <SPLIT distance="550" swimtime="00:08:09.01" />
                    <SPLIT distance="600" swimtime="00:08:54.84" />
                    <SPLIT distance="650" swimtime="00:09:41.21" />
                    <SPLIT distance="700" swimtime="00:10:27.41" />
                    <SPLIT distance="750" swimtime="00:11:12.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="343" reactiontime="+79" swimtime="00:03:12.21" resultid="4322" heatid="7330" lane="3" entrytime="00:03:24.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:32.89" />
                    <SPLIT distance="150" swimtime="00:02:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="302" reactiontime="+80" swimtime="00:01:24.21" resultid="4323" heatid="7371" lane="4" entrytime="00:01:32.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="375" reactiontime="+77" swimtime="00:01:26.41" resultid="4324" heatid="7411" lane="6" entrytime="00:01:36.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="266" reactiontime="+90" swimtime="00:06:42.14" resultid="4325" heatid="8150" lane="0" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:37.06" />
                    <SPLIT distance="150" swimtime="00:02:33.43" />
                    <SPLIT distance="200" swimtime="00:03:26.27" />
                    <SPLIT distance="250" swimtime="00:04:18.36" />
                    <SPLIT distance="300" swimtime="00:05:11.18" />
                    <SPLIT distance="350" swimtime="00:05:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="398" reactiontime="+72" swimtime="00:00:38.80" resultid="4326" heatid="7542" lane="5" entrytime="00:00:41.95" />
                <RESULT eventid="1721" points="299" reactiontime="+81" swimtime="00:05:49.60" resultid="4327" heatid="7569" lane="0" entrytime="00:06:22.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="150" swimtime="00:02:08.14" />
                    <SPLIT distance="200" swimtime="00:02:52.41" />
                    <SPLIT distance="250" swimtime="00:03:36.47" />
                    <SPLIT distance="300" swimtime="00:04:20.98" />
                    <SPLIT distance="350" swimtime="00:05:05.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarosław" gender="M" lastname="Bystry" nation="POL" athleteid="4313">
              <RESULTS>
                <RESULT eventid="1076" points="382" reactiontime="+74" swimtime="00:00:27.92" resultid="4314" heatid="7263" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1288" points="388" reactiontime="+67" swimtime="00:01:01.59" resultid="4315" heatid="7362" lane="9" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="302" reactiontime="+65" swimtime="00:01:14.87" resultid="4316" heatid="7384" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="310" reactiontime="+68" swimtime="00:00:32.11" resultid="4317" heatid="7445" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1689" points="333" reactiontime="+69" swimtime="00:00:36.41" resultid="4318" heatid="7556" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-27" firstname="Rafał" gender="M" lastname="Domeracki" nation="POL" athleteid="4328">
              <RESULTS>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="4329" heatid="7303" lane="4" entrytime="00:21:12.30" />
                <RESULT eventid="1288" status="WDR" swimtime="00:00:00.00" resultid="4330" heatid="7352" lane="5" entrytime="00:01:11.60" />
                <RESULT eventid="1513" status="WDR" swimtime="00:00:00.00" resultid="4331" heatid="7481" lane="2" entrytime="00:02:32.50" />
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="4332" heatid="7578" lane="5" entrytime="00:05:21.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-10" firstname="Karolina" gender="F" lastname="Drach" nation="POL" athleteid="4333">
              <RESULTS>
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="4334" heatid="7309" lane="2" entrytime="00:00:45.53" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4335" heatid="7342" lane="4" entrytime="00:01:25.60" />
                <RESULT eventid="1465" points="126" reactiontime="+87" swimtime="00:01:49.51" resultid="4336" heatid="7454" lane="9" entrytime="00:01:45.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-08" firstname="Siergiej" gender="M" lastname="Kulinicz" nation="POL" athleteid="4309">
              <RESULTS>
                <RESULT eventid="1076" points="356" reactiontime="+88" swimtime="00:00:28.56" resultid="4310" heatid="7258" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4311" heatid="7355" lane="7" entrytime="00:01:12.99" />
                <RESULT eventid="1449" points="242" reactiontime="+84" swimtime="00:00:34.89" resultid="4312" heatid="7439" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-20" firstname="Tomasz" gender="M" lastname="Matras" nation="POL" athleteid="4344">
              <RESULTS>
                <RESULT eventid="1076" points="359" reactiontime="+99" swimtime="00:00:28.48" resultid="4345" heatid="7262" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4346" heatid="7360" lane="9" entrytime="00:01:04.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="4305">
              <RESULTS>
                <RESULT eventid="1288" points="181" swimtime="00:01:19.41" resultid="4306" heatid="7352" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach. (Time: 12:23)" eventid="1320" status="DSQ" swimtime="00:01:33.40" resultid="4307" heatid="7379" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="185" reactiontime="+60" swimtime="00:01:37.57" resultid="4308" heatid="7418" lane="7" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-07-28" firstname="Marek" gender="M" lastname="Piórkowski" nation="POL" athleteid="4295">
              <RESULTS>
                <RESULT eventid="1076" points="135" swimtime="00:00:39.47" resultid="4296" heatid="7249" lane="6" entrytime="00:00:40.22" />
                <RESULT eventid="1224" points="103" reactiontime="+82" swimtime="00:00:47.35" resultid="4297" heatid="7318" lane="9" entrytime="00:00:52.00" />
                <RESULT eventid="1288" points="99" swimtime="00:01:36.94" resultid="4298" heatid="7350" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="87" reactiontime="+95" swimtime="00:01:50.29" resultid="4299" heatid="7459" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="4282">
              <RESULTS>
                <RESULT eventid="1076" points="661" reactiontime="+63" swimtime="00:00:23.25" resultid="4283" heatid="7270" lane="3" entrytime="00:00:23.00" />
                <RESULT eventid="1256" points="656" reactiontime="+64" swimtime="00:02:18.23" resultid="4284" heatid="7339" lane="4" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:06.15" />
                    <SPLIT distance="150" swimtime="00:01:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="689" reactiontime="+65" swimtime="00:00:56.90" resultid="4285" heatid="7390" lane="3" entrytime="00:00:57.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="746" reactiontime="+63" swimtime="00:01:01.31" resultid="4286" heatid="7425" lane="4" entrytime="00:01:01.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="736" reactiontime="+64" swimtime="00:00:27.96" resultid="4287" heatid="7561" lane="4" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-05-06" firstname="Monika" gender="F" lastname="Winnicka" nation="POL" athleteid="4337">
              <RESULTS>
                <RESULT eventid="1059" points="291" reactiontime="+83" swimtime="00:00:34.60" resultid="4338" heatid="7241" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="4339" heatid="7311" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4340" heatid="7346" lane="1" entrytime="00:01:09.69" />
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="4341" heatid="7455" lane="2" entrytime="00:01:30.64" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4342" heatid="7472" lane="6" entrytime="00:02:36.40" />
                <RESULT eventid="1721" status="WDR" swimtime="00:00:00.00" resultid="4343" heatid="7567" lane="2" entrytime="00:05:30.55" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1391" points="201" reactiontime="+98" swimtime="00:02:34.25" resultid="4351" heatid="7404" lane="9" entrytime="00:02:32.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4295" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="4288" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4313" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4305" number="4" reactiontime="+92" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1391" status="WDR" swimtime="00:00:00.00" resultid="4352" heatid="7403" lane="7" entrytime="00:02:06.54">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4282" number="1" />
                    <RELAYPOSITION athleteid="4305" number="2" />
                    <RELAYPOSITION athleteid="4313" number="3" />
                    <RELAYPOSITION athleteid="4344" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1545" points="385" reactiontime="+60" swimtime="00:01:52.36" resultid="4353" heatid="7495" lane="6" entrytime="00:01:48.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.30" />
                    <SPLIT distance="100" swimtime="00:00:51.18" />
                    <SPLIT distance="150" swimtime="00:01:25.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4282" number="1" reactiontime="+60" status="DSQ" />
                    <RELAYPOSITION athleteid="4309" number="2" reactiontime="+38" status="DSQ" />
                    <RELAYPOSITION athleteid="4344" number="3" reactiontime="+91" status="DSQ" />
                    <RELAYPOSITION athleteid="4313" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1545" status="WDR" swimtime="00:00:00.00" resultid="4354" heatid="7493" lane="5" entrytime="00:02:24.20">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4328" number="1" />
                    <RELAYPOSITION athleteid="4305" number="2" />
                    <RELAYPOSITION athleteid="4288" number="3" />
                    <RELAYPOSITION athleteid="4295" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utraciły kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 13:31)" eventid="1368" reactiontime="+79" status="DSQ" swimtime="00:02:39.72" resultid="4348" heatid="7400" lane="2" entrytime="00:02:39.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:17.86" />
                    <SPLIT distance="150" swimtime="00:01:59.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4337" number="1" reactiontime="+79" status="DSQ" />
                    <RELAYPOSITION athleteid="4319" number="2" reactiontime="-6" status="DSQ" />
                    <RELAYPOSITION athleteid="4300" number="3" reactiontime="+65" status="DSQ" />
                    <RELAYPOSITION athleteid="4333" number="4" reactiontime="+64" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1529" points="288" reactiontime="+78" swimtime="00:02:22.17" resultid="4349" heatid="7490" lane="5" entrytime="00:02:16.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:48.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4337" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4319" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="4333" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="4300" number="4" reactiontime="+3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="349" reactiontime="+69" swimtime="00:02:04.76" resultid="4347" heatid="7288" lane="6" entrytime="00:02:03.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:35.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4313" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4337" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4319" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="4309" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1705" points="378" reactiontime="+80" status="EXH" swimtime="00:02:13.22" resultid="4350" heatid="7564" lane="7" entrytime="00:02:12.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4300" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4282" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="4313" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4319" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="14" clubid="2834" name="KS Niezrzeszeni.pl" shortname="Niezrzeszeni.pl">
          <CONTACT name="KS_Niezrzeszeni_pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="2835">
              <RESULTS>
                <RESULT eventid="1108" points="159" reactiontime="+88" swimtime="00:03:22.20" resultid="2836" heatid="7279" lane="2" entrytime="00:03:28.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="194" reactiontime="+97" swimtime="00:12:45.44" resultid="2837" heatid="7298" lane="3" entrytime="00:12:37.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="150" swimtime="00:02:18.19" />
                    <SPLIT distance="200" swimtime="00:03:06.91" />
                    <SPLIT distance="250" swimtime="00:03:56.47" />
                    <SPLIT distance="300" swimtime="00:04:45.13" />
                    <SPLIT distance="350" swimtime="00:05:34.26" />
                    <SPLIT distance="400" swimtime="00:06:23.60" />
                    <SPLIT distance="450" swimtime="00:07:13.13" />
                    <SPLIT distance="500" swimtime="00:08:02.12" />
                    <SPLIT distance="550" swimtime="00:08:50.98" />
                    <SPLIT distance="600" swimtime="00:09:39.74" />
                    <SPLIT distance="650" swimtime="00:10:28.47" />
                    <SPLIT distance="700" swimtime="00:11:16.46" />
                    <SPLIT distance="750" swimtime="00:12:02.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="153" reactiontime="+71" swimtime="00:00:41.53" resultid="2838" heatid="7316" lane="0" />
                <RESULT eventid="1256" points="135" reactiontime="+89" swimtime="00:03:54.04" resultid="2839" heatid="7334" lane="1" entrytime="00:03:51.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                    <SPLIT distance="100" swimtime="00:01:51.31" />
                    <SPLIT distance="150" swimtime="00:02:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="200" reactiontime="+75" swimtime="00:02:49.66" resultid="2840" heatid="7478" lane="6" entrytime="00:02:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                    <SPLIT distance="150" swimtime="00:02:05.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="168" reactiontime="+66" swimtime="00:03:11.10" resultid="2841" heatid="7532" lane="2" entrytime="00:03:09.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:33.69" />
                    <SPLIT distance="150" swimtime="00:02:23.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="188" swimtime="00:06:10.11" resultid="2842" heatid="7581" lane="5" entrytime="00:06:15.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:28.78" />
                    <SPLIT distance="150" swimtime="00:02:17.00" />
                    <SPLIT distance="200" swimtime="00:03:05.42" />
                    <SPLIT distance="250" swimtime="00:03:53.32" />
                    <SPLIT distance="300" swimtime="00:04:41.73" />
                    <SPLIT distance="350" swimtime="00:05:28.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00914" nation="POL" region="14" clubid="2889" name="KS Polonia Warszawa" shortname="Polonia Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Lucjan" gender="M" lastname="Prządło" nation="POL" athleteid="2888">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2890" heatid="7248" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1224" status="WDR" swimtime="00:00:00.00" resultid="2891" heatid="7316" lane="4" entrytime="00:01:05.00" />
                <RESULT eventid="1256" status="WDR" swimtime="00:00:00.00" resultid="2892" entrytime="00:05:15.00" />
                <RESULT eventid="1417" status="WDR" swimtime="00:00:00.00" resultid="2893" heatid="7414" lane="5" entrytime="00:02:05.00" />
                <RESULT eventid="1481" status="WDR" swimtime="00:00:00.00" resultid="2894" heatid="7460" lane="1" entrytime="00:02:15.00" />
                <RESULT eventid="1657" status="WDR" swimtime="00:00:00.00" resultid="2895" heatid="7529" lane="5" entrytime="00:05:15.00" />
                <RESULT eventid="1689" status="WDR" swimtime="00:00:00.00" resultid="2896" heatid="7547" lane="1" entrytime="00:01:00.01" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PRRZE" nation="POL" region="08" clubid="3640" name="KS Prestige Rzeszów" shortname="Prestige Rzeszów">
          <ATHLETES>
            <ATHLETE birthdate="1995-12-15" firstname="Justyna" gender="F" lastname="Gałuszka" nation="POL" athleteid="3639">
              <RESULTS>
                <RESULT eventid="1240" points="328" reactiontime="+86" swimtime="00:03:15.09" resultid="5298" heatid="7327" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:35.49" />
                    <SPLIT distance="150" swimtime="00:02:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="358" reactiontime="+84" swimtime="00:01:19.58" resultid="5299" heatid="7368" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="349" reactiontime="+83" swimtime="00:01:28.51" resultid="5300" heatid="7407" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="5301" heatid="7430" lane="4" entrytime="00:00:36.80" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5302" heatid="7537" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="01" clubid="3699" name="KS Rekin Świebodzice" shortname="Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="3700">
              <RESULTS>
                <RESULT eventid="1059" points="535" reactiontime="+78" swimtime="00:00:28.24" resultid="3701" heatid="7244" lane="2" entrytime="00:00:29.50" entrycourse="SCM" />
                <RESULT eventid="1240" points="428" reactiontime="+75" swimtime="00:02:58.50" resultid="3702" heatid="7327" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:10.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="500" reactiontime="+75" swimtime="00:01:03.29" resultid="3703" heatid="7347" lane="2" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="490" reactiontime="+75" swimtime="00:01:19.06" resultid="3704" heatid="7413" lane="0" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="438" reactiontime="+75" swimtime="00:02:25.33" resultid="3705" heatid="7473" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                    <SPLIT distance="150" swimtime="00:01:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="503" reactiontime="+72" swimtime="00:00:35.89" resultid="3706" heatid="7544" lane="3" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="3707">
              <RESULTS>
                <RESULT eventid="1092" points="360" reactiontime="+73" swimtime="00:02:51.23" resultid="3708" heatid="7274" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="373" reactiontime="+76" swimtime="00:21:17.15" resultid="3709" heatid="7300" lane="2" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                    <SPLIT distance="200" swimtime="00:02:45.41" />
                    <SPLIT distance="250" swimtime="00:03:28.28" />
                    <SPLIT distance="300" swimtime="00:04:11.40" />
                    <SPLIT distance="350" swimtime="00:04:54.90" />
                    <SPLIT distance="400" swimtime="00:05:38.14" />
                    <SPLIT distance="450" swimtime="00:06:21.41" />
                    <SPLIT distance="500" swimtime="00:07:04.85" />
                    <SPLIT distance="550" swimtime="00:07:48.47" />
                    <SPLIT distance="600" swimtime="00:08:32.12" />
                    <SPLIT distance="650" swimtime="00:09:15.51" />
                    <SPLIT distance="700" swimtime="00:09:58.93" />
                    <SPLIT distance="750" swimtime="00:10:41.74" />
                    <SPLIT distance="800" swimtime="00:11:24.69" />
                    <SPLIT distance="850" swimtime="00:12:07.69" />
                    <SPLIT distance="900" swimtime="00:12:50.53" />
                    <SPLIT distance="950" swimtime="00:13:33.21" />
                    <SPLIT distance="1000" swimtime="00:14:15.84" />
                    <SPLIT distance="1050" swimtime="00:14:58.53" />
                    <SPLIT distance="1100" swimtime="00:15:41.04" />
                    <SPLIT distance="1150" swimtime="00:16:24.33" />
                    <SPLIT distance="1200" swimtime="00:17:06.98" />
                    <SPLIT distance="1250" swimtime="00:17:49.27" />
                    <SPLIT distance="1300" swimtime="00:18:31.85" />
                    <SPLIT distance="1350" swimtime="00:19:13.54" />
                    <SPLIT distance="1400" swimtime="00:19:55.45" />
                    <SPLIT distance="1450" swimtime="00:20:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="350" reactiontime="+71" swimtime="00:03:10.79" resultid="3710" heatid="7331" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="150" swimtime="00:02:20.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="271" reactiontime="+75" swimtime="00:03:04.71" resultid="3711" heatid="7393" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="150" swimtime="00:02:15.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="385" reactiontime="+70" swimtime="00:02:31.77" resultid="3712" heatid="7470" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="355" reactiontime="+76" swimtime="00:06:05.36" resultid="3713" heatid="8151" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:02:14.25" />
                    <SPLIT distance="200" swimtime="00:03:00.27" />
                    <SPLIT distance="250" swimtime="00:03:50.19" />
                    <SPLIT distance="300" swimtime="00:04:41.30" />
                    <SPLIT distance="350" swimtime="00:05:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="364" reactiontime="+70" swimtime="00:00:39.99" resultid="3714" heatid="7543" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1721" points="385" reactiontime="+70" swimtime="00:05:21.29" resultid="3715" heatid="7567" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                    <SPLIT distance="200" swimtime="00:02:39.34" />
                    <SPLIT distance="250" swimtime="00:03:20.40" />
                    <SPLIT distance="300" swimtime="00:04:02.13" />
                    <SPLIT distance="350" swimtime="00:04:42.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="3716">
              <RESULTS>
                <RESULT eventid="1076" points="519" reactiontime="+85" swimtime="00:00:25.20" resultid="3717" heatid="7268" lane="7" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1108" points="520" reactiontime="+81" swimtime="00:02:16.33" resultid="3718" heatid="7285" lane="3" entrytime="00:02:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:01:02.93" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="498" reactiontime="+64" swimtime="00:00:28.03" resultid="3719" heatid="7316" lane="8" />
                <RESULT eventid="1320" points="514" reactiontime="+79" swimtime="00:01:02.71" resultid="3720" heatid="7389" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="512" reactiontime="+77" swimtime="00:00:27.17" resultid="3721" heatid="7447" lane="4" entrytime="00:00:28.90" />
                <RESULT eventid="1481" points="508" reactiontime="+63" swimtime="00:01:01.22" resultid="3722" heatid="7467" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="514" reactiontime="+81" swimtime="00:01:00.01" resultid="3723" heatid="7520" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="501" reactiontime="+63" swimtime="00:02:12.94" resultid="3724" heatid="7536" lane="5" entrytime="00:02:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:38.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="5193" name="KU AZS UAM Poznań" shortname="AZS UAM Poznań">
          <CONTACT email="swimteamuam@gmail.com" name="Sterczyński" phone="693840114" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-13" firstname="Kamil" gender="M" lastname="Bernaś" nation="POL" athleteid="5203">
              <RESULTS>
                <RESULT eventid="1076" points="398" reactiontime="+72" swimtime="00:00:27.54" resultid="5204" heatid="7264" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1288" points="368" reactiontime="+71" swimtime="00:01:02.71" resultid="5205" heatid="7361" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="328" reactiontime="+73" swimtime="00:01:12.83" resultid="5206" heatid="7384" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="348" reactiontime="+68" swimtime="00:00:30.91" resultid="5207" heatid="7447" lane="0" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-12" firstname="Joanna" gender="F" lastname="Chomicz" nation="POL" athleteid="5208">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="5209" heatid="7242" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="5210" heatid="7313" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="5211" heatid="7432" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5212" heatid="7545" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="5213">
              <RESULTS>
                <RESULT eventid="1076" points="345" reactiontime="+79" swimtime="00:00:28.87" resultid="5214" heatid="7259" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1288" points="306" reactiontime="+73" swimtime="00:01:06.64" resultid="5215" heatid="7359" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="266" reactiontime="+77" swimtime="00:01:18.10" resultid="5216" heatid="7384" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="282" reactiontime="+81" swimtime="00:00:33.13" resultid="5217" heatid="7441" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-05-10" firstname="Tomasz" gender="M" lastname="Juszkiewicz" nation="POL" athleteid="5194">
              <RESULTS>
                <RESULT eventid="1224" points="111" reactiontime="+69" swimtime="00:00:46.13" resultid="5195" heatid="7319" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1288" points="190" reactiontime="+92" swimtime="00:01:18.04" resultid="5196" heatid="7354" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="155" reactiontime="+96" swimtime="00:00:40.44" resultid="5197" heatid="7438" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="5198" heatid="7462" lane="8" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-27" firstname="Bartosz" gender="M" lastname="Kaczmarek" nation="POL" athleteid="5218">
              <RESULTS>
                <RESULT eventid="1076" points="354" swimtime="00:00:28.62" resultid="5219" heatid="7262" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1224" points="263" reactiontime="+78" swimtime="00:00:34.66" resultid="5220" heatid="7320" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1288" points="302" reactiontime="+75" swimtime="00:01:06.97" resultid="5221" heatid="7360" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="236" reactiontime="+92" swimtime="00:01:19.02" resultid="5222" heatid="7463" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="288" reactiontime="+73" swimtime="00:02:30.34" resultid="5223" heatid="7481" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-19" firstname="Damian" gender="M" lastname="Kowalik" nation="POL" athleteid="5224">
              <RESULTS>
                <RESULT eventid="1076" points="493" reactiontime="+67" swimtime="00:00:25.63" resultid="5225" heatid="7269" lane="1" entrytime="00:00:25.00" />
                <RESULT eventid="1320" points="505" reactiontime="+58" swimtime="00:01:03.08" resultid="5226" heatid="7390" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="549" reactiontime="+56" swimtime="00:00:26.56" resultid="5227" heatid="7450" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1625" points="478" reactiontime="+57" swimtime="00:01:01.49" resultid="5228" heatid="7521" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" athleteid="5229">
              <RESULTS>
                <RESULT eventid="1076" points="566" reactiontime="+65" swimtime="00:00:24.49" resultid="5230" heatid="7269" lane="8" entrytime="00:00:25.00" />
                <RESULT eventid="1224" points="557" reactiontime="+66" swimtime="00:00:26.99" resultid="5231" heatid="7326" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1449" points="621" reactiontime="+62" swimtime="00:00:25.49" resultid="5232" heatid="7451" lane="2" entrytime="00:00:25.00" />
                <RESULT eventid="1481" points="553" reactiontime="+65" swimtime="00:00:59.54" resultid="5233" heatid="7467" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="576" reactiontime="+62" swimtime="00:00:57.76" resultid="5234" heatid="7522" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-01" firstname="Dariusz" gender="M" lastname="Perkowski" nation="POL" athleteid="5199">
              <RESULTS>
                <RESULT eventid="1076" points="254" swimtime="00:00:31.96" resultid="5200" heatid="7258" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1288" points="175" reactiontime="+75" swimtime="00:01:20.25" resultid="5201" heatid="7355" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="183" reactiontime="+73" swimtime="00:00:38.29" resultid="5202" heatid="7441" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-05" firstname="Marek" gender="M" lastname="Serafin" nation="POL" athleteid="5235">
              <RESULTS>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="5236" heatid="7321" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1288" points="250" reactiontime="+82" swimtime="00:01:11.26" resultid="5237" heatid="7356" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="166" swimtime="00:00:39.50" resultid="5238" heatid="7439" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1513" points="208" reactiontime="+76" swimtime="00:02:47.67" resultid="5239" heatid="7480" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:22.06" />
                    <SPLIT distance="150" swimtime="00:02:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5240" heatid="7533" lane="8" entrytime="00:03:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Sterczyńska" nation="POL" athleteid="5241">
              <RESULTS>
                <RESULT eventid="1059" points="600" reactiontime="+82" swimtime="00:00:27.18" resultid="5242" heatid="7245" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1272" points="619" reactiontime="+78" swimtime="00:00:58.96" resultid="5243" heatid="7348" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="567" reactiontime="+77" swimtime="00:01:08.24" resultid="5244" heatid="7376" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="498" reactiontime="+76" swimtime="00:00:30.75" resultid="5245" heatid="7434" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1673" points="495" reactiontime="+78" swimtime="00:00:36.08" resultid="5246" heatid="7545" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" athleteid="5247">
              <RESULTS>
                <RESULT eventid="1076" points="438" reactiontime="+76" swimtime="00:00:26.67" resultid="5248" heatid="7267" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5249" heatid="7284" lane="5" entrytime="00:02:25.00" />
                <RESULT eventid="1320" points="465" reactiontime="+67" swimtime="00:01:04.84" resultid="5250" heatid="7389" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="461" reactiontime="+66" swimtime="00:00:28.14" resultid="5251" heatid="7446" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1657" points="379" reactiontime="+66" swimtime="00:02:25.88" resultid="5252" heatid="7536" lane="7" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:45.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-20" firstname="Krzysztof" gender="M" lastname="Strzelczyk" nation="POL" athleteid="5253">
              <RESULTS>
                <RESULT eventid="1076" points="177" reactiontime="+96" swimtime="00:00:36.06" resultid="5254" heatid="7253" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1288" points="153" reactiontime="+90" swimtime="00:01:23.95" resultid="5255" heatid="7352" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="133" reactiontime="+88" swimtime="00:01:38.31" resultid="5256" heatid="7379" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="151" reactiontime="+81" swimtime="00:00:40.83" resultid="5257" heatid="7438" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1513" points="158" reactiontime="+87" swimtime="00:03:03.57" resultid="5258" heatid="7478" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:02:16.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="185" reactiontime="+84" swimtime="00:00:44.29" resultid="5259" heatid="7550" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-10-02" firstname="Anna" gender="F" lastname="Szczucińska" nation="POL" athleteid="5260">
              <RESULTS>
                <RESULT eventid="1059" points="233" swimtime="00:00:37.25" resultid="5261" heatid="7241" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1207" points="140" reactiontime="+83" swimtime="00:00:49.33" resultid="5262" heatid="7310" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1304" points="152" reactiontime="+79" swimtime="00:01:45.71" resultid="5263" heatid="7372" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="123" reactiontime="+47" swimtime="00:00:48.98" resultid="5264" heatid="7428" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1673" points="172" reactiontime="+92" swimtime="00:00:51.35" resultid="5265" heatid="7541" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-23" firstname="Joanna" gender="F" lastname="Szymanowska" nation="POL" athleteid="5266">
              <RESULTS>
                <RESULT eventid="1272" points="312" reactiontime="+93" swimtime="00:01:14.02" resultid="5267" heatid="7346" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="292" reactiontime="+82" swimtime="00:01:33.89" resultid="5268" heatid="7411" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5269" heatid="7543" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="481" reactiontime="+61" swimtime="00:01:44.37" resultid="5270" heatid="7496" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.44" />
                    <SPLIT distance="100" swimtime="00:00:49.67" />
                    <SPLIT distance="150" swimtime="00:01:15.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5229" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5224" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="5247" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="5218" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="513" reactiontime="+67" swimtime="00:01:52.94" resultid="5272" heatid="7406" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                    <SPLIT distance="100" swimtime="00:00:59.78" />
                    <SPLIT distance="150" swimtime="00:01:25.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5229" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5247" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="5224" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="5203" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="226" reactiontime="+98" swimtime="00:02:14.18" resultid="5271" heatid="7494" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:42.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5194" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="5253" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="5199" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="5235" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1391" points="238" reactiontime="+79" swimtime="00:02:25.82" resultid="5273" heatid="7404" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5218" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="5253" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5213" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5235" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" status="WDR" swimtime="00:00:00.00" resultid="5274" heatid="7491" lane="7" entrytime="00:02:07.00" />
                <RESULT eventid="1368" status="WDR" swimtime="00:00:00.00" resultid="5275" heatid="7399" lane="3" entrytime="00:02:20.00" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="464" swimtime="00:01:53.50" resultid="5276" heatid="7289" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:29.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5260" number="1" />
                    <RELAYPOSITION athleteid="5241" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="5224" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5229" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" status="WDR" swimtime="00:00:00.00" resultid="5277" heatid="7562" lane="2" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1705" points="389" reactiontime="+64" swimtime="00:02:12.04" resultid="5278" heatid="7562" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:01:45.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5229" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5260" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5224" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="5241" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZWAR" nation="POL" region="14" clubid="2129" name="KU AZS UW Warszawa" shortname="AZS UW Warszawa">
          <CONTACT city="Warszawa" email="azsuwswimming@gmail.com" name="Eugeniusz Puzan" phone="574-504-127" state="MAZ" street="Krakowskie Przedmieњcie 24" zip="00-325" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" athleteid="2174">
              <RESULTS>
                <RESULT eventid="1076" points="514" reactiontime="+76" swimtime="00:00:25.28" resultid="2175" heatid="7268" lane="1" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1288" points="544" reactiontime="+71" swimtime="00:00:55.04" resultid="2176" heatid="7367" lane="9" entrytime="00:00:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="504" reactiontime="+76" swimtime="00:02:04.85" resultid="2177" heatid="7487" lane="0" entrytime="00:02:05.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                    <SPLIT distance="100" swimtime="00:00:59.46" />
                    <SPLIT distance="150" swimtime="00:01:31.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="2165">
              <RESULTS>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2166" heatid="7358" lane="8" entrytime="00:01:06.90" entrycourse="SCM" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="2167" heatid="7420" lane="2" entrytime="00:01:26.00" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2168" heatid="7552" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-20" firstname="Marika" gender="F" lastname="Florczak" nation="POL" athleteid="2141">
              <RESULTS>
                <RESULT eventid="1272" points="480" reactiontime="+78" swimtime="00:01:04.17" resultid="2142" heatid="7347" lane="5" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="507" reactiontime="+81" swimtime="00:02:18.47" resultid="2143" heatid="7474" lane="6" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="484" reactiontime="+77" swimtime="00:04:57.79" resultid="2144" heatid="7566" lane="7" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:48.28" />
                    <SPLIT distance="200" swimtime="00:02:26.51" />
                    <SPLIT distance="250" swimtime="00:03:04.23" />
                    <SPLIT distance="300" swimtime="00:03:42.96" />
                    <SPLIT distance="350" swimtime="00:04:21.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-05-26" firstname="Rafal" gender="M" lastname="Godlewski" nation="POL" athleteid="2153">
              <RESULTS>
                <RESULT eventid="1076" points="241" swimtime="00:00:32.53" resultid="2154" heatid="7247" lane="0" />
                <RESULT eventid="1256" points="352" reactiontime="+76" swimtime="00:02:50.12" resultid="2155" heatid="7338" lane="0" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="481" reactiontime="+72" swimtime="00:01:10.94" resultid="2156" heatid="7424" lane="0" entrytime="00:01:16.00" entrycourse="SCY">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="514" reactiontime="+74" swimtime="00:00:31.51" resultid="2157" heatid="7559" lane="3" entrytime="00:00:33.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-08-27" firstname="Edyta" gender="F" lastname="Ilcewicz" nation="POL" athleteid="2178">
              <RESULTS>
                <RESULT eventid="1272" points="520" reactiontime="+74" swimtime="00:01:02.48" resultid="2179" heatid="7348" lane="1" entrytime="00:01:00.00" entrycourse="SCY">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="488" reactiontime="+72" swimtime="00:00:30.95" resultid="2180" heatid="7434" lane="1" entrytime="00:00:30.00" entrycourse="SCY" />
                <RESULT eventid="1673" points="483" reactiontime="+75" swimtime="00:00:36.38" resultid="2181" heatid="7545" lane="1" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-17" firstname="Piotr" gender="M" lastname="Kister" nation="POL" athleteid="2158">
              <RESULTS>
                <RESULT eventid="1256" points="287" reactiontime="+77" swimtime="00:03:02.07" resultid="2159" heatid="7337" lane="7" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:02:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="307" reactiontime="+80" swimtime="00:02:40.31" resultid="2160" heatid="7397" lane="6" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="340" reactiontime="+83" swimtime="00:01:19.60" resultid="2161" heatid="7422" lane="4" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="378" reactiontime="+81" swimtime="00:00:30.06" resultid="2162" heatid="7444" lane="0" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1625" points="343" reactiontime="+82" swimtime="00:01:08.66" resultid="2163" heatid="7518" lane="7" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="358" reactiontime="+79" swimtime="00:00:35.54" resultid="2164" heatid="7556" lane="7" entrytime="00:00:36.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-08-25" firstname="Krzysztof" gender="M" lastname="Micorek" nation="POL" athleteid="2187">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2188" heatid="7269" lane="0" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2189" heatid="7390" lane="1" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2190" heatid="7450" lane="9" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2191" heatid="7560" lane="5" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="8161" heatid="7315" lane="6" late="yes" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="8162" heatid="7512" lane="9" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-08-11" firstname="Artur" gender="M" lastname="Milczarek" nation="POL" athleteid="2182">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2183" heatid="7265" lane="1" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2184" heatid="7364" lane="3" entrytime="00:00:58.00" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2185" heatid="7487" lane="1" entrytime="00:02:05.00" entrycourse="SCM" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="2186" heatid="7521" lane="2" entrytime="00:01:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-05" firstname="Yauheni" gender="M" lastname="Puzan" nation="POL" athleteid="2134">
              <RESULTS>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2135" heatid="7315" lane="5" />
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="2136" heatid="7398" lane="5" entrytime="00:02:10.00" entrycourse="SCM" />
                <RESULT eventid="1449" points="515" reactiontime="+70" swimtime="00:00:27.13" resultid="2137" heatid="7451" lane="7" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1513" points="442" reactiontime="+71" swimtime="00:02:10.45" resultid="2138" heatid="7475" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:01.42" />
                    <SPLIT distance="150" swimtime="00:01:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="534" reactiontime="+70" swimtime="00:00:59.25" resultid="2139" heatid="7522" lane="6" entrytime="00:00:56.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="385" reactiontime="+71" swimtime="00:00:34.69" resultid="2140" heatid="7546" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rebas" nation="POL" athleteid="2130">
              <RESULTS>
                <RESULT eventid="1288" points="616" reactiontime="+78" swimtime="00:00:52.80" resultid="2131" heatid="7363" lane="3" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="595" reactiontime="+76" swimtime="00:01:58.12" resultid="2132" heatid="7486" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="100" swimtime="00:00:55.69" />
                    <SPLIT distance="150" swimtime="00:01:26.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="540" reactiontime="+77" swimtime="00:00:59.01" resultid="2133" heatid="7521" lane="7" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-10" firstname="Daniel" gender="M" lastname="Rzadkowski" nation="POL" athleteid="2145">
              <RESULTS>
                <RESULT eventid="1076" points="706" reactiontime="+77" swimtime="00:00:22.75" resultid="2146" heatid="7270" lane="4" entrytime="00:00:22.50" entrycourse="SCM" />
                <RESULT eventid="1288" points="718" reactiontime="+70" swimtime="00:00:50.17" resultid="2147" heatid="7367" lane="3" entrytime="00:00:49.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-25" firstname="Michal" gender="M" lastname="Uziak" nation="POL" athleteid="2149">
              <RESULTS>
                <RESULT eventid="1076" points="391" reactiontime="+80" swimtime="00:00:27.69" resultid="2150" heatid="7263" lane="2" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1288" points="411" reactiontime="+75" swimtime="00:01:00.43" resultid="2151" heatid="7361" lane="1" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="402" reactiontime="+84" swimtime="00:02:14.60" resultid="2152" heatid="7484" lane="5" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="150" swimtime="00:01:38.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M">
              <RESULTS>
                <RESULT eventid="1545" points="596" reactiontime="+73" status="EXH" swimtime="00:01:37.16" resultid="8230" heatid="7492" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.66" />
                    <SPLIT distance="100" swimtime="00:00:48.03" />
                    <SPLIT distance="150" swimtime="00:01:12.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2145" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2130" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="2174" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="2134" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LALUB" nation="POL" region="03" clubid="2109" name="Labosport Lublin">
          <ATHLETES>
            <ATHLETE birthdate="1978-04-24" firstname="Tomasz" gender="M" lastname="Pomierny " nation="POL" athleteid="2108">
              <RESULTS>
                <RESULT eventid="1156" points="311" swimtime="00:10:54.40" resultid="2110" heatid="7296" lane="8" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:01:57.44" />
                    <SPLIT distance="200" swimtime="00:02:37.95" />
                    <SPLIT distance="250" swimtime="00:03:19.13" />
                    <SPLIT distance="300" swimtime="00:04:00.29" />
                    <SPLIT distance="350" swimtime="00:04:41.41" />
                    <SPLIT distance="400" swimtime="00:05:23.28" />
                    <SPLIT distance="450" swimtime="00:06:05.02" />
                    <SPLIT distance="500" swimtime="00:06:46.69" />
                    <SPLIT distance="550" swimtime="00:07:28.62" />
                    <SPLIT distance="600" swimtime="00:08:10.26" />
                    <SPLIT distance="650" swimtime="00:08:51.98" />
                    <SPLIT distance="700" swimtime="00:09:33.77" />
                    <SPLIT distance="750" swimtime="00:10:15.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2111" heatid="7358" lane="9" entrytime="00:01:07.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="2112" heatid="8156" lane="5" entrytime="00:06:25.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2113" heatid="7578" lane="7" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" region="04" clubid="2032" name="LC Gorzów Wlkp.">
          <CONTACT city="Os. Poznańskie" email="stan_ley@poczta.fm" name="Kaczmarek" phone="600277732" state="LUBUS" street="Liliowa 9" zip="66-446" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Kaczmarek" nation="POL" athleteid="2033">
              <RESULTS>
                <RESULT eventid="1059" points="535" reactiontime="+75" swimtime="00:00:28.23" resultid="2034" heatid="7244" lane="4" entrytime="00:00:28.12" />
                <RESULT eventid="1092" points="567" reactiontime="+79" swimtime="00:02:27.22" resultid="2035" heatid="7275" lane="4" entrytime="00:02:27.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="561" reactiontime="+77" swimtime="00:01:00.91" resultid="2036" heatid="7348" lane="8" entrytime="00:01:00.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="572" reactiontime="+76" swimtime="00:01:08.07" resultid="2037" heatid="7376" lane="3" entrytime="00:01:07.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="570" reactiontime="+81" swimtime="00:02:13.14" resultid="2038" heatid="7474" lane="3" entrytime="00:02:11.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="547" reactiontime="+79" swimtime="00:05:16.46" resultid="2039" heatid="8151" lane="4" entrytime="00:05:16.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                    <SPLIT distance="200" swimtime="00:02:34.90" />
                    <SPLIT distance="250" swimtime="00:03:18.92" />
                    <SPLIT distance="300" swimtime="00:04:03.87" />
                    <SPLIT distance="350" swimtime="00:04:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="535" reactiontime="+76" swimtime="00:00:35.16" resultid="2040" heatid="7545" lane="2" entrytime="00:00:35.94" />
                <RESULT eventid="1721" points="529" reactiontime="+79" swimtime="00:04:49.11" resultid="2041" heatid="7566" lane="5" entrytime="00:04:45.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:45.31" />
                    <SPLIT distance="200" swimtime="00:02:22.69" />
                    <SPLIT distance="250" swimtime="00:03:00.18" />
                    <SPLIT distance="300" swimtime="00:03:37.17" />
                    <SPLIT distance="350" swimtime="00:04:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" athleteid="2042">
              <RESULTS>
                <RESULT eventid="1108" points="457" reactiontime="+78" swimtime="00:02:22.23" resultid="2043" heatid="7284" lane="4" entrytime="00:02:24.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="467" reactiontime="+80" swimtime="00:09:31.36" resultid="2044" heatid="7294" lane="5" entrytime="00:09:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:02:20.45" />
                    <SPLIT distance="250" swimtime="00:02:57.29" />
                    <SPLIT distance="300" swimtime="00:03:33.51" />
                    <SPLIT distance="350" swimtime="00:04:09.80" />
                    <SPLIT distance="400" swimtime="00:04:46.03" />
                    <SPLIT distance="450" swimtime="00:05:22.20" />
                    <SPLIT distance="500" swimtime="00:05:58.56" />
                    <SPLIT distance="550" swimtime="00:06:35.24" />
                    <SPLIT distance="600" swimtime="00:07:11.59" />
                    <SPLIT distance="650" swimtime="00:07:48.16" />
                    <SPLIT distance="700" swimtime="00:08:24.51" />
                    <SPLIT distance="750" swimtime="00:09:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="419" reactiontime="+77" swimtime="00:02:40.53" resultid="2045" heatid="7339" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:01:59.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="426" reactiontime="+76" swimtime="00:02:23.79" resultid="2046" heatid="7398" lane="2" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="469" reactiontime="+75" swimtime="00:02:07.88" resultid="2047" heatid="7485" lane="3" entrytime="00:02:11.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="430" reactiontime="+79" swimtime="00:05:11.89" resultid="2048" heatid="8158" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:50.77" />
                    <SPLIT distance="200" swimtime="00:02:31.77" />
                    <SPLIT distance="250" swimtime="00:03:16.43" />
                    <SPLIT distance="300" swimtime="00:04:01.23" />
                    <SPLIT distance="350" swimtime="00:04:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="421" reactiontime="+75" swimtime="00:01:04.11" resultid="2049" heatid="7520" lane="8" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="467" reactiontime="+76" swimtime="00:04:33.57" resultid="2050" heatid="7573" lane="6" entrytime="00:04:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.56" />
                    <SPLIT distance="150" swimtime="00:01:41.85" />
                    <SPLIT distance="200" swimtime="00:02:16.92" />
                    <SPLIT distance="250" swimtime="00:02:51.91" />
                    <SPLIT distance="300" swimtime="00:03:26.85" />
                    <SPLIT distance="350" swimtime="00:04:00.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LTTWR" nation="POL" region="01" clubid="5835" name="Litwin Triathlon Team Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1994-02-04" firstname="Paulina" gender="F" lastname="Krajcarska" nation="POL" athleteid="5841">
              <RESULTS>
                <RESULT eventid="1059" points="318" reactiontime="+86" swimtime="00:00:33.57" resultid="5842" heatid="7239" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1272" points="295" reactiontime="+87" swimtime="00:01:15.47" resultid="5843" heatid="7343" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="302" reactiontime="+78" swimtime="00:00:36.30" resultid="5844" heatid="7429" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1497" points="286" reactiontime="+78" swimtime="00:02:47.56" resultid="5845" heatid="7472" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-07-13" firstname="Agata" gender="F" lastname="Litwin-Żurad" nation="POL" athleteid="5834">
              <RESULTS>
                <RESULT eventid="1059" points="498" reactiontime="+92" swimtime="00:00:28.92" resultid="5836" heatid="7243" lane="6" entrytime="00:00:30.99" />
                <RESULT eventid="1140" points="514" reactiontime="+95" swimtime="00:09:58.11" resultid="5837" heatid="7290" lane="6" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                    <SPLIT distance="200" swimtime="00:02:26.11" />
                    <SPLIT distance="250" swimtime="00:03:03.94" />
                    <SPLIT distance="300" swimtime="00:03:41.26" />
                    <SPLIT distance="350" swimtime="00:04:18.54" />
                    <SPLIT distance="400" swimtime="00:04:56.14" />
                    <SPLIT distance="450" swimtime="00:05:33.65" />
                    <SPLIT distance="500" swimtime="00:06:11.95" />
                    <SPLIT distance="550" swimtime="00:06:49.90" />
                    <SPLIT distance="600" swimtime="00:07:28.04" />
                    <SPLIT distance="650" swimtime="00:08:06.07" />
                    <SPLIT distance="700" swimtime="00:08:44.34" />
                    <SPLIT distance="750" swimtime="00:09:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="523" reactiontime="+93" swimtime="00:01:02.33" resultid="5838" heatid="7347" lane="3" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="469" reactiontime="+86" swimtime="00:01:10.82" resultid="5839" heatid="7458" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="500" reactiontime="+87" swimtime="00:04:54.68" resultid="5840" heatid="7566" lane="9" entrytime="00:05:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:45.16" />
                    <SPLIT distance="200" swimtime="00:02:22.94" />
                    <SPLIT distance="250" swimtime="00:03:01.08" />
                    <SPLIT distance="300" swimtime="00:03:39.11" />
                    <SPLIT distance="350" swimtime="00:04:17.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LOWAR" nation="POL" region="14" clubid="2211" name="Lochte Swimming Academy Warszawa" shortname="Lochte Swimming Academy W-wa">
          <ATHLETES>
            <ATHLETE birthdate="1993-12-12" firstname="Adam" gender="M" lastname="Dubiel" nation="POL" athleteid="3334">
              <RESULTS>
                <RESULT eventid="1288" points="682" reactiontime="+70" swimtime="00:00:51.05" resultid="6872" heatid="7349" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski masters kategoria A" eventid="1513" points="720" reactiontime="+68" swimtime="00:01:50.83" resultid="8231" heatid="7488" lane="6" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                    <SPLIT distance="100" swimtime="00:00:54.90" />
                    <SPLIT distance="150" swimtime="00:01:23.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-25" firstname="Patryk" gender="M" lastname="Gąsior" nation="POL" athleteid="5791">
              <RESULTS>
                <RESULT eventid="1352" points="634" reactiontime="+78" swimtime="00:02:05.97" resultid="5792" heatid="7398" lane="4" entrytime="00:02:05.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="100" swimtime="00:01:00.47" />
                    <SPLIT distance="150" swimtime="00:01:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="658" reactiontime="+77" swimtime="00:01:54.22" resultid="5793" heatid="7488" lane="5" entrytime="00:01:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="100" swimtime="00:00:55.98" />
                    <SPLIT distance="150" swimtime="00:01:24.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="615" reactiontime="+82" swimtime="00:04:36.83" resultid="5794" heatid="8158" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:39.39" />
                    <SPLIT distance="200" swimtime="00:02:15.35" />
                    <SPLIT distance="250" swimtime="00:02:54.40" />
                    <SPLIT distance="300" swimtime="00:03:33.14" />
                    <SPLIT distance="350" swimtime="00:04:06.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-09-20" firstname="Mateusz" gender="M" lastname="Kraśniewski" nation="POL" athleteid="2207">
              <RESULTS>
                <RESULT eventid="1076" points="319" swimtime="00:00:29.63" resultid="2208" heatid="7258" lane="2" entrytime="00:00:29.94" />
                <RESULT eventid="1449" points="271" reactiontime="+92" swimtime="00:00:33.58" resultid="2209" heatid="7443" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-09" firstname="Adam" gender="M" lastname="Markowski" nation="POL" athleteid="2512">
              <RESULTS>
                <RESULT eventid="1076" points="361" reactiontime="+92" swimtime="00:00:28.44" resultid="2513" heatid="7260" lane="8" entrytime="00:00:28.60" />
                <RESULT eventid="1288" points="335" reactiontime="+87" swimtime="00:01:04.65" resultid="2514" heatid="7354" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-20" firstname="Daria" gender="F" lastname="Sieradzka" nation="POL" athleteid="2227">
              <RESULTS>
                <RESULT eventid="1059" points="163" reactiontime="+78" swimtime="00:00:41.93" resultid="2228" heatid="7236" lane="2" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-07" firstname="Michał" gender="M" lastname="Sieńko" nation="POL" athleteid="2210">
              <RESULTS>
                <RESULT eventid="1076" points="479" reactiontime="+66" swimtime="00:00:25.88" resultid="2212" heatid="7267" lane="4" entrytime="00:00:25.73" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2213" heatid="7387" lane="4" entrytime="00:01:07.50" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2214" heatid="7559" lane="8" entrytime="00:00:33.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-11" firstname="Marta" gender="F" lastname="Smycz" nation="POL" athleteid="2743">
              <RESULTS>
                <RESULT eventid="1059" points="254" reactiontime="+92" swimtime="00:00:36.18" resultid="2744" heatid="7238" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1207" points="167" reactiontime="+47" swimtime="00:00:46.58" resultid="2745" heatid="7309" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1465" points="162" swimtime="00:01:40.90" resultid="2746" heatid="7454" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-09" firstname="Konrad" gender="M" lastname="Szymański" nation="POL" athleteid="3335" />
            <ATHLETE birthdate="1981-09-28" firstname="Łukasz" gender="M" lastname="Zandberg " nation="POL" athleteid="2238">
              <RESULTS>
                <RESULT eventid="1076" points="259" swimtime="00:00:31.76" resultid="2239" heatid="7254" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-16" firstname="Karol" gender="M" lastname="Zientarski" nation="POL" athleteid="2458">
              <RESULTS>
                <RESULT eventid="1076" points="93" reactiontime="+87" swimtime="00:00:44.67" resultid="2459" heatid="7248" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="606" reactiontime="+79" swimtime="00:01:36.66" resultid="2215" heatid="7496" lane="4" entrytime="00:01:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="100" swimtime="00:00:47.40" />
                    <SPLIT distance="150" swimtime="00:01:11.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5791" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2210" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="3334" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="3335" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="230" reactiontime="+83" swimtime="00:02:13.43" resultid="2874" heatid="7492" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="100" swimtime="00:00:56.83" />
                    <SPLIT distance="150" swimtime="00:01:26.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2512" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2207" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2238" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2458" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X">
              <RESULTS>
                <RESULT eventid="1124" points="274" reactiontime="+97" swimtime="00:02:15.31" resultid="2875" heatid="7286" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="100" swimtime="00:00:57.43" />
                    <SPLIT distance="150" swimtime="00:01:33.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2512" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="2207" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="2743" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2227" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAHAI" nation="ISR" clubid="2124" name="Maccabi Haifa Israel Club" shortname="Maccabi Haifa">
          <ATHLETES>
            <ATHLETE birthdate="1950-11-08" firstname="Ailon" gender="M" lastname="Tobis" nation="POL" athleteid="2123">
              <RESULTS>
                <RESULT eventid="1076" points="270" reactiontime="+93" swimtime="00:00:31.31" resultid="2125" heatid="7256" lane="8" entrytime="00:00:31.50" />
                <RESULT eventid="1224" points="190" reactiontime="+53" swimtime="00:00:38.65" resultid="2126" heatid="7320" lane="6" entrytime="00:00:39.20" />
                <RESULT eventid="1481" points="168" reactiontime="+89" swimtime="00:01:28.43" resultid="2127" heatid="7463" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="247" reactiontime="+89" swimtime="00:01:11.61" resultid="2128" heatid="7357" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MABIA" nation="POL" region="09" clubid="2428" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="MB" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="2473">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2474" heatid="7254" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1320" points="203" reactiontime="+98" swimtime="00:01:25.50" resultid="2475" heatid="7380" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="238" reactiontime="+87" swimtime="00:01:29.71" resultid="2476" heatid="7419" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="189" reactiontime="+96" swimtime="00:00:37.88" resultid="2477" heatid="7440" lane="9" entrytime="00:00:36.50" />
                <RESULT eventid="1689" points="281" reactiontime="+98" swimtime="00:00:38.54" resultid="2478" heatid="7553" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2479" heatid="7580" lane="7" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="2480">
              <RESULTS>
                <RESULT eventid="1092" points="425" reactiontime="+79" swimtime="00:02:42.04" resultid="2481" heatid="7274" lane="3" entrytime="00:02:45.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:15.86" />
                    <SPLIT distance="150" swimtime="00:02:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="412" reactiontime="+81" swimtime="00:20:35.40" resultid="2482" heatid="7300" lane="4" entrytime="00:19:46.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                    <SPLIT distance="200" swimtime="00:02:34.77" />
                    <SPLIT distance="250" swimtime="00:03:15.38" />
                    <SPLIT distance="300" swimtime="00:03:55.98" />
                    <SPLIT distance="350" swimtime="00:04:36.79" />
                    <SPLIT distance="400" swimtime="00:05:17.90" />
                    <SPLIT distance="450" swimtime="00:05:59.55" />
                    <SPLIT distance="500" swimtime="00:06:41.13" />
                    <SPLIT distance="550" swimtime="00:07:22.24" />
                    <SPLIT distance="600" swimtime="00:08:03.95" />
                    <SPLIT distance="650" swimtime="00:08:45.79" />
                    <SPLIT distance="700" swimtime="00:09:27.30" />
                    <SPLIT distance="750" swimtime="00:10:08.97" />
                    <SPLIT distance="800" swimtime="00:10:50.65" />
                    <SPLIT distance="850" swimtime="00:11:32.25" />
                    <SPLIT distance="900" swimtime="00:12:14.28" />
                    <SPLIT distance="950" swimtime="00:12:56.40" />
                    <SPLIT distance="1000" swimtime="00:13:38.52" />
                    <SPLIT distance="1050" swimtime="00:14:20.94" />
                    <SPLIT distance="1100" swimtime="00:15:02.97" />
                    <SPLIT distance="1150" swimtime="00:15:44.24" />
                    <SPLIT distance="1200" swimtime="00:16:26.12" />
                    <SPLIT distance="1250" swimtime="00:17:08.64" />
                    <SPLIT distance="1300" swimtime="00:17:51.03" />
                    <SPLIT distance="1350" swimtime="00:18:33.66" />
                    <SPLIT distance="1400" swimtime="00:19:15.91" />
                    <SPLIT distance="1450" swimtime="00:19:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="486" reactiontime="+83" swimtime="00:02:20.39" resultid="2483" heatid="7474" lane="7" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="480" reactiontime="+79" swimtime="00:04:58.56" resultid="2484" heatid="7566" lane="2" entrytime="00:04:56.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                    <SPLIT distance="200" swimtime="00:02:27.30" />
                    <SPLIT distance="250" swimtime="00:03:05.77" />
                    <SPLIT distance="300" swimtime="00:03:44.32" />
                    <SPLIT distance="350" swimtime="00:04:22.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="2461">
              <RESULTS>
                <RESULT eventid="1076" points="236" reactiontime="+91" swimtime="00:00:32.77" resultid="2462" heatid="7255" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="1224" points="213" reactiontime="+72" swimtime="00:00:37.18" resultid="2463" heatid="7321" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1256" points="199" reactiontime="+96" swimtime="00:03:25.77" resultid="2464" heatid="7335" lane="5" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:36.91" />
                    <SPLIT distance="150" swimtime="00:02:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="209" reactiontime="+79" swimtime="00:01:22.24" resultid="2465" heatid="7463" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="151" reactiontime="+97" swimtime="00:07:21.45" resultid="2466" heatid="8156" lane="0" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:44.76" />
                    <SPLIT distance="150" swimtime="00:02:37.73" />
                    <SPLIT distance="200" swimtime="00:03:30.53" />
                    <SPLIT distance="250" swimtime="00:04:34.36" />
                    <SPLIT distance="300" swimtime="00:05:39.58" />
                    <SPLIT distance="350" swimtime="00:06:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="185" reactiontime="+79" swimtime="00:03:05.13" resultid="2467" heatid="7532" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:30.51" />
                    <SPLIT distance="150" swimtime="00:02:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2468" heatid="7581" lane="2" entrytime="00:06:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="2469">
              <RESULTS>
                <RESULT eventid="1059" points="239" reactiontime="+85" swimtime="00:00:36.90" resultid="2470" heatid="7238" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1272" points="216" reactiontime="+90" swimtime="00:01:23.65" resultid="2471" heatid="7342" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="159" swimtime="00:03:23.71" resultid="2472" heatid="7469" lane="3" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:35.59" />
                    <SPLIT distance="150" swimtime="00:02:29.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MACZE" nation="POL" region="11" clubid="2000" name="Masters Częstochowa">
          <ATHLETES>
            <ATHLETE birthdate="1951-06-06" firstname="Jolanta" gender="F" lastname="Lipińska" nation="POL" athleteid="2071">
              <RESULTS>
                <RESULT eventid="1240" points="30" swimtime="00:07:11.59" resultid="2072" heatid="7327" lane="2" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.27" />
                    <SPLIT distance="100" swimtime="00:03:34.59" />
                    <SPLIT distance="150" swimtime="00:05:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="21" swimtime="00:03:24.67" resultid="2073" heatid="7368" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="29" swimtime="00:03:21.35" resultid="2074" heatid="7407" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="25" reactiontime="+94" swimtime="00:03:07.54" resultid="2075" heatid="7452" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="29" reactiontime="+78" swimtime="00:06:24.90" resultid="2076" heatid="7524" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.55" />
                    <SPLIT distance="100" swimtime="00:03:09.20" />
                    <SPLIT distance="150" swimtime="00:04:49.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="40" swimtime="00:01:22.88" resultid="2077" heatid="7537" lane="6" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="1999">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2001" heatid="7252" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="2002" heatid="7298" lane="9" entrytime="00:13:43.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2003" heatid="7479" lane="9" entrytime="00:02:54.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="2004" heatid="8153" lane="1" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="2005" heatid="7514" lane="4" entrytime="00:01:41.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2006" heatid="7582" lane="4" entrytime="00:06:35.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" nation="POL" region="03" clubid="2747" name="Masters Kraśnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" internet="www.masterskrasnik.cba.pl" name="MIchalczyk" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-204" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="2755">
              <RESULTS>
                <RESULT eventid="1076" points="93" reactiontime="+91" swimtime="00:00:44.67" resultid="2756" heatid="7250" lane="9" entrytime="00:00:49.10" />
                <RESULT eventid="1108" points="79" reactiontime="+92" swimtime="00:04:15.06" resultid="2757" heatid="7277" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.27" />
                    <SPLIT distance="100" swimtime="00:02:02.55" />
                    <SPLIT distance="150" swimtime="00:03:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="79" reactiontime="+94" swimtime="00:00:51.66" resultid="2758" heatid="7317" lane="6" entrytime="00:00:55.45" />
                <RESULT eventid="1320" points="84" reactiontime="+95" swimtime="00:01:54.59" resultid="2759" heatid="7378" lane="9" entrytime="00:01:58.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="59" reactiontime="+85" swimtime="00:00:55.83" resultid="2760" heatid="7436" lane="3" entrytime="00:00:59.10" />
                <RESULT eventid="1625" points="41" swimtime="00:02:18.44" resultid="2761" heatid="7513" lane="8" entrytime="00:02:15.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="2748">
              <RESULTS>
                <RESULT eventid="1108" points="92" swimtime="00:04:02.23" resultid="2749" heatid="7278" lane="9" entrytime="00:04:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                    <SPLIT distance="100" swimtime="00:01:57.66" />
                    <SPLIT distance="150" swimtime="00:03:09.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="107" reactiontime="+90" swimtime="00:00:46.70" resultid="2750" heatid="7317" lane="3" entrytime="00:00:53.20" />
                <RESULT eventid="1320" points="104" reactiontime="+98" swimtime="00:01:46.75" resultid="2751" heatid="7377" lane="4" entrytime="00:01:59.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="84" reactiontime="+92" swimtime="00:01:51.39" resultid="2752" heatid="7461" lane="8" entrytime="00:01:58.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="2753" heatid="8154" lane="1" entrytime="00:08:50.40" />
                <RESULT eventid="1657" points="92" reactiontime="+90" swimtime="00:03:53.15" resultid="2754" heatid="7530" lane="2" entrytime="00:04:14.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                    <SPLIT distance="100" swimtime="00:01:51.84" />
                    <SPLIT distance="150" swimtime="00:02:55.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="2762">
              <RESULTS>
                <RESULT eventid="1156" points="76" swimtime="00:17:24.70" resultid="2763" heatid="7299" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.80" />
                    <SPLIT distance="100" swimtime="00:02:07.55" />
                    <SPLIT distance="150" swimtime="00:03:12.82" />
                    <SPLIT distance="200" swimtime="00:04:18.53" />
                    <SPLIT distance="250" swimtime="00:05:25.59" />
                    <SPLIT distance="300" swimtime="00:06:32.94" />
                    <SPLIT distance="350" swimtime="00:07:40.30" />
                    <SPLIT distance="400" swimtime="00:08:46.53" />
                    <SPLIT distance="450" swimtime="00:09:53.77" />
                    <SPLIT distance="500" swimtime="00:11:00.39" />
                    <SPLIT distance="550" swimtime="00:12:07.12" />
                    <SPLIT distance="600" swimtime="00:13:12.83" />
                    <SPLIT distance="650" swimtime="00:14:18.49" />
                    <SPLIT distance="700" swimtime="00:15:22.27" />
                    <SPLIT distance="750" swimtime="00:16:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="44" swimtime="00:05:06.01" resultid="2764" heatid="7395" lane="0" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.61" />
                    <SPLIT distance="100" swimtime="00:02:19.07" />
                    <SPLIT distance="150" swimtime="00:03:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="2765" heatid="8154" lane="2" entrytime="00:08:45.00" />
                <RESULT eventid="1625" points="55" swimtime="00:02:06.30" resultid="2766" heatid="7513" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="151" swimtime="00:00:47.36" resultid="2767" heatid="7549" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKK" nation="POL" region="07" clubid="2454" name="Masters Kędzierzyn-Koźle">
          <ATHLETES>
            <ATHLETE birthdate="1948-11-01" firstname="Stanisław" gender="M" lastname="Zajfert" nation="POL" athleteid="2453">
              <RESULTS>
                <RESULT eventid="1224" points="113" reactiontime="+90" swimtime="00:00:45.91" resultid="2455" heatid="7318" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1481" points="110" reactiontime="+90" swimtime="00:01:41.96" resultid="2456" heatid="7462" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="113" reactiontime="+95" swimtime="00:03:37.97" resultid="2457" heatid="7531" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.17" />
                    <SPLIT distance="100" swimtime="00:01:50.44" />
                    <SPLIT distance="150" swimtime="00:02:47.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOST" nation="POL" region="14" clubid="2516" name="Masters Ostrołęka">
          <ATHLETES>
            <ATHLETE birthdate="1990-12-06" firstname="Adam" gender="M" lastname="Janczewski" nation="POL" athleteid="2515">
              <RESULTS>
                <RESULT eventid="1108" points="466" swimtime="00:02:21.31" resultid="2517" heatid="7285" lane="0" entrytime="00:02:23.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="387" reactiontime="+90" swimtime="00:10:08.01" resultid="2518" heatid="7295" lane="2" entrytime="00:10:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                    <SPLIT distance="200" swimtime="00:02:25.74" />
                    <SPLIT distance="250" swimtime="00:03:03.73" />
                    <SPLIT distance="300" swimtime="00:03:41.72" />
                    <SPLIT distance="350" swimtime="00:04:20.73" />
                    <SPLIT distance="400" swimtime="00:04:59.93" />
                    <SPLIT distance="450" swimtime="00:05:39.17" />
                    <SPLIT distance="500" swimtime="00:06:19.11" />
                    <SPLIT distance="550" swimtime="00:06:58.07" />
                    <SPLIT distance="600" swimtime="00:07:37.38" />
                    <SPLIT distance="650" swimtime="00:08:16.00" />
                    <SPLIT distance="700" swimtime="00:08:54.81" />
                    <SPLIT distance="750" swimtime="00:09:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2519" heatid="7389" lane="8" entrytime="00:01:03.50" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2520" heatid="7487" lane="9" entrytime="00:02:05.76" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2521" heatid="7574" lane="1" entrytime="00:04:44.85" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOZ" nation="POL" region="15" clubid="2217" name="Masters Poznań">
          <ATHLETES>
            <ATHLETE birthdate="1962-03-22" firstname="Piotr" gender="M" lastname="Burzyński" nation="POL" athleteid="2216">
              <RESULTS>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="2218" heatid="7298" lane="7" entrytime="00:13:15.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="2219" heatid="7334" lane="2" entrytime="00:03:42.00" />
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="2220" heatid="7396" lane="0" entrytime="00:03:45.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="2221" heatid="8155" lane="8" entrytime="00:07:48.00" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="2222" heatid="7514" lane="6" entrytime="00:01:45.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2223" heatid="7580" lane="9" entrytime="00:06:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-25" firstname="Joanna" gender="F" lastname="Grzeszczuk " nation="POL" athleteid="2548">
              <RESULTS>
                <RESULT eventid="1400" points="533" reactiontime="+68" swimtime="00:01:16.91" resultid="2549" heatid="7413" lane="5" entrytime="00:01:16.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="460" reactiontime="+69" swimtime="00:00:31.58" resultid="2550" heatid="7433" lane="3" entrytime="00:00:30.98" />
                <RESULT eventid="1673" points="559" reactiontime="+69" swimtime="00:00:34.65" resultid="2551" heatid="7545" lane="5" entrytime="00:00:34.08" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAWAR" nation="POL" region="14" clubid="2065" name="Masters Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1955-04-09" firstname="Anna" gender="F" lastname="Błazucka" nation="POL" athleteid="2588">
              <RESULTS>
                <RESULT eventid="1059" points="74" reactiontime="+82" swimtime="00:00:54.40" resultid="2589" heatid="7235" lane="6" entrytime="00:00:54.86" />
                <RESULT eventid="1207" points="46" reactiontime="+81" swimtime="00:01:11.39" resultid="2590" heatid="7307" lane="8" entrytime="00:01:18.78" />
                <RESULT eventid="1304" points="51" reactiontime="+96" swimtime="00:02:32.06" resultid="2591" heatid="7368" lane="4" entrytime="00:02:41.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="61" swimtime="00:02:38.38" resultid="2592" heatid="7407" lane="5" entrytime="00:02:49.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="40" reactiontime="+73" swimtime="00:02:40.27" resultid="2593" heatid="7452" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="67" reactiontime="+87" swimtime="00:01:10.31" resultid="2594" heatid="7537" lane="3" entrytime="00:01:13.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-08" firstname="Anna" gender="F" lastname="Gonet" nation="POL" athleteid="2485">
              <RESULTS>
                <RESULT eventid="1207" points="284" reactiontime="+69" swimtime="00:00:39.04" resultid="2486" heatid="7307" lane="9" />
                <RESULT eventid="1304" points="269" swimtime="00:01:27.45" resultid="2487" heatid="7368" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="2488" heatid="7452" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-11-14" firstname="Konrad" gender="M" lastname="Jajecznik" nation="POL" athleteid="2064">
              <RESULTS>
                <RESULT eventid="1076" points="190" reactiontime="+99" swimtime="00:00:35.20" resultid="2066" heatid="7252" lane="1" entrytime="00:00:35.55" />
                <RESULT eventid="1288" points="171" reactiontime="+84" swimtime="00:01:20.86" resultid="2067" heatid="7353" lane="9" entrytime="00:01:22.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="178" reactiontime="+85" swimtime="00:00:38.60" resultid="2069" heatid="7438" lane="4" entrytime="00:00:38.27" />
                <RESULT eventid="1513" points="168" reactiontime="+82" swimtime="00:02:59.93" resultid="2070" heatid="7477" lane="7" entrytime="00:03:17.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                    <SPLIT distance="150" swimtime="00:02:13.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-13" firstname="Paweł" gender="M" lastname="Kapusta" nation="POL" athleteid="6489">
              <RESULTS>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6490" heatid="7443" lane="8" entrytime="00:00:31.65" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="6491" heatid="7579" lane="6" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="2772">
              <RESULTS>
                <RESULT eventid="1256" points="201" reactiontime="+43" swimtime="00:03:24.87" resultid="2869" heatid="7332" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="100" swimtime="00:01:34.58" />
                    <SPLIT distance="150" swimtime="00:02:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="127" reactiontime="+73" swimtime="00:03:34.83" resultid="2870" heatid="7396" lane="8" entrytime="00:03:33.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:37.74" />
                    <SPLIT distance="150" swimtime="00:02:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2871" heatid="7438" lane="5" entrytime="00:00:38.60" />
                <RESULT eventid="1625" points="158" reactiontime="+60" swimtime="00:01:28.83" resultid="2872" heatid="7515" lane="7" entrytime="00:01:31.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="215" swimtime="00:00:42.14" resultid="2873" heatid="7551" lane="3" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01806" nation="POL" region="06" clubid="2240" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" license="501806600060" athleteid="2261">
              <RESULTS>
                <RESULT eventid="1092" points="82" swimtime="00:04:40.23" resultid="2262" heatid="7271" lane="7" entrytime="00:04:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.37" />
                    <SPLIT distance="100" swimtime="00:02:20.21" />
                    <SPLIT distance="150" swimtime="00:03:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="69" swimtime="00:37:13.86" resultid="2263" heatid="7301" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.69" />
                    <SPLIT distance="100" swimtime="00:02:09.16" />
                    <SPLIT distance="150" swimtime="00:03:21.03" />
                    <SPLIT distance="200" swimtime="00:04:32.93" />
                    <SPLIT distance="250" swimtime="00:05:46.75" />
                    <SPLIT distance="300" swimtime="00:07:00.63" />
                    <SPLIT distance="350" swimtime="00:08:11.23" />
                    <SPLIT distance="400" swimtime="00:09:24.78" />
                    <SPLIT distance="450" swimtime="00:10:36.52" />
                    <SPLIT distance="500" swimtime="00:11:52.84" />
                    <SPLIT distance="550" swimtime="00:13:05.91" />
                    <SPLIT distance="600" swimtime="00:14:19.77" />
                    <SPLIT distance="650" swimtime="00:15:33.08" />
                    <SPLIT distance="700" swimtime="00:16:48.55" />
                    <SPLIT distance="750" swimtime="00:18:03.79" />
                    <SPLIT distance="800" swimtime="00:19:18.42" />
                    <SPLIT distance="850" swimtime="00:20:34.54" />
                    <SPLIT distance="900" swimtime="00:21:48.56" />
                    <SPLIT distance="950" swimtime="00:23:03.94" />
                    <SPLIT distance="1000" swimtime="00:24:19.17" />
                    <SPLIT distance="1050" swimtime="00:25:35.56" />
                    <SPLIT distance="1100" swimtime="00:26:53.75" />
                    <SPLIT distance="1150" swimtime="00:28:09.88" />
                    <SPLIT distance="1200" swimtime="00:29:28.01" />
                    <SPLIT distance="1250" swimtime="00:30:45.75" />
                    <SPLIT distance="1300" swimtime="00:32:04.48" />
                    <SPLIT distance="1350" swimtime="00:33:23.37" />
                    <SPLIT distance="1400" swimtime="00:34:39.49" />
                    <SPLIT distance="1450" swimtime="00:35:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="93" swimtime="00:04:56.16" resultid="2264" heatid="7327" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.90" />
                    <SPLIT distance="100" swimtime="00:02:18.01" />
                    <SPLIT distance="150" swimtime="00:03:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="78" swimtime="00:02:12.20" resultid="2265" heatid="7369" lane="9" entrytime="00:02:10.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="93" swimtime="00:02:17.36" resultid="2266" heatid="7407" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="78" swimtime="00:04:18.10" resultid="2267" heatid="7468" lane="4" entrytime="00:04:04.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.70" />
                    <SPLIT distance="100" swimtime="00:01:58.95" />
                    <SPLIT distance="150" swimtime="00:03:08.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="97" swimtime="00:01:02.02" resultid="2268" heatid="7537" lane="1" />
                <RESULT eventid="1721" points="76" swimtime="00:09:11.10" resultid="2269" heatid="7571" lane="2" entrytime="00:08:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.45" />
                    <SPLIT distance="100" swimtime="00:01:59.99" />
                    <SPLIT distance="150" swimtime="00:03:08.80" />
                    <SPLIT distance="200" swimtime="00:04:18.06" />
                    <SPLIT distance="250" swimtime="00:05:29.30" />
                    <SPLIT distance="300" swimtime="00:06:42.59" />
                    <SPLIT distance="350" swimtime="00:07:52.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" license="501806700050" athleteid="2248">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="2249" heatid="7334" lane="5" entrytime="00:03:35.00" entrycourse="SCM" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="2250" heatid="7420" lane="0" entrytime="00:01:28.71" entrycourse="SCM" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2251" heatid="7438" lane="6" entrytime="00:00:39.01" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2252" heatid="7554" lane="1" entrytime="00:00:38.41" entrycourse="SCM" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2253" heatid="7581" lane="8" entrytime="00:06:31.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="2254">
              <RESULTS>
                <RESULT eventid="1224" points="74" reactiontime="+89" swimtime="00:00:52.85" resultid="2255" heatid="7317" lane="7" entrytime="00:00:56.00" entrycourse="SCM" />
                <RESULT eventid="1320" points="89" reactiontime="+98" swimtime="00:01:52.35" resultid="2256" heatid="7378" lane="0" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="64" reactiontime="+93" swimtime="00:00:54.20" resultid="2257" heatid="7437" lane="8" entrytime="00:00:51.00" entrycourse="SCM" />
                <RESULT eventid="1481" points="65" swimtime="00:02:01.33" resultid="2258" heatid="7460" lane="2" entrytime="00:02:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="58" reactiontime="+59" swimtime="00:02:03.58" resultid="2259" heatid="7513" lane="7" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="95" reactiontime="+89" swimtime="00:00:55.31" resultid="2260" heatid="7547" lane="5" entrytime="00:00:58.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-27" firstname="Michał" gender="M" lastname="Klupa" nation="POL" athleteid="2280">
              <RESULTS>
                <RESULT eventid="1108" points="463" reactiontime="+77" swimtime="00:02:21.64" resultid="2281" heatid="7284" lane="2" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="478" reactiontime="+59" swimtime="00:00:28.40" resultid="2282" heatid="7326" lane="7" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1320" points="465" reactiontime="+72" swimtime="00:01:04.87" resultid="2283" heatid="7389" lane="3" entrytime="00:01:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="479" reactiontime="+63" swimtime="00:01:02.44" resultid="2284" heatid="7467" lane="1" entrytime="00:01:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="411" reactiontime="+74" swimtime="00:05:16.60" resultid="2285" heatid="8153" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                    <SPLIT distance="200" swimtime="00:02:28.64" />
                    <SPLIT distance="250" swimtime="00:03:15.44" />
                    <SPLIT distance="300" swimtime="00:04:04.01" />
                    <SPLIT distance="350" swimtime="00:04:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="448" reactiontime="+60" swimtime="00:02:17.98" resultid="2286" heatid="7536" lane="6" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="150" swimtime="00:01:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2287" heatid="7575" lane="5" entrytime="00:04:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="2288">
              <RESULTS>
                <RESULT eventid="1076" points="402" reactiontime="+82" swimtime="00:00:27.44" resultid="2289" heatid="7262" lane="4" entrytime="00:00:27.60" entrycourse="SCM" />
                <RESULT eventid="1156" points="383" swimtime="00:10:10.19" resultid="2290" heatid="7295" lane="0" entrytime="00:11:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:46.16" />
                    <SPLIT distance="200" swimtime="00:02:24.83" />
                    <SPLIT distance="250" swimtime="00:03:03.55" />
                    <SPLIT distance="350" swimtime="00:04:20.96" />
                    <SPLIT distance="400" swimtime="00:05:00.19" />
                    <SPLIT distance="450" swimtime="00:05:39.40" />
                    <SPLIT distance="500" swimtime="00:06:18.34" />
                    <SPLIT distance="550" swimtime="00:06:57.87" />
                    <SPLIT distance="650" swimtime="00:08:15.73" />
                    <SPLIT distance="700" swimtime="00:08:54.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="333" reactiontime="+85" swimtime="00:02:53.26" resultid="2291" heatid="7332" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                    <SPLIT distance="150" swimtime="00:02:08.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2292" heatid="7361" lane="2" entrytime="00:01:02.00" entrycourse="SCM" />
                <RESULT eventid="1417" points="360" reactiontime="+96" swimtime="00:01:18.13" resultid="2293" heatid="7423" lane="8" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2294" heatid="7484" lane="9" entrytime="00:02:18.00" entrycourse="SCM" />
                <RESULT eventid="1689" points="399" reactiontime="+79" swimtime="00:00:34.29" resultid="2295" heatid="7557" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2296" heatid="7576" lane="8" entrytime="00:05:05.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="2241">
              <RESULTS>
                <RESULT eventid="1076" points="70" swimtime="00:00:48.99" resultid="2242" heatid="7247" lane="3" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1224" points="41" reactiontime="+75" swimtime="00:01:04.43" resultid="2243" heatid="7317" lane="9" entrytime="00:01:05.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="66" swimtime="00:01:50.93" resultid="2244" heatid="7350" lane="2" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="51" swimtime="00:02:29.05" resultid="2245" heatid="7418" lane="6" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="60" swimtime="00:04:13.28" resultid="2246" heatid="7475" lane="5" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.82" />
                    <SPLIT distance="100" swimtime="00:02:00.55" />
                    <SPLIT distance="150" swimtime="00:03:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="57" swimtime="00:01:05.55" resultid="2247" heatid="7546" lane="5" entrytime="00:01:10.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-08-12" firstname="Konrad" gender="M" lastname="Plutecki" nation="POL" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1076" points="489" reactiontime="+66" swimtime="00:00:25.71" resultid="2316" heatid="7266" lane="3" entrytime="00:00:26.26" entrycourse="SCM" />
                <RESULT eventid="1156" points="305" reactiontime="+72" swimtime="00:10:58.03" resultid="2317" heatid="7295" lane="5" entrytime="00:10:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.54" />
                    <SPLIT distance="200" swimtime="00:02:28.67" />
                    <SPLIT distance="250" swimtime="00:03:08.92" />
                    <SPLIT distance="300" swimtime="00:03:48.81" />
                    <SPLIT distance="350" swimtime="00:04:29.63" />
                    <SPLIT distance="400" swimtime="00:05:11.15" />
                    <SPLIT distance="450" swimtime="00:05:53.51" />
                    <SPLIT distance="500" swimtime="00:06:36.41" />
                    <SPLIT distance="550" swimtime="00:07:19.41" />
                    <SPLIT distance="600" swimtime="00:08:02.90" />
                    <SPLIT distance="650" swimtime="00:08:46.67" />
                    <SPLIT distance="700" swimtime="00:09:31.13" />
                    <SPLIT distance="750" swimtime="00:10:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="310" reactiontime="+72" swimtime="00:00:32.80" resultid="2318" heatid="7322" lane="4" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="1288" points="495" reactiontime="+70" swimtime="00:00:56.78" resultid="2319" heatid="7364" lane="8" entrytime="00:00:58.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="2320" heatid="7423" lane="0" entrytime="00:01:18.18" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2321" heatid="7484" lane="6" entrytime="00:02:15.15" entrycourse="SCM" />
                <RESULT eventid="1657" points="335" reactiontime="+78" swimtime="00:02:32.02" resultid="2322" heatid="7535" lane="9" entrytime="00:02:33.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:13.85" />
                    <SPLIT distance="150" swimtime="00:01:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2323" heatid="7555" lane="9" entrytime="00:00:37.37" entrycourse="SCM" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2324" heatid="7576" lane="6" entrytime="00:04:59.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="2306">
              <RESULTS>
                <RESULT eventid="1059" points="105" swimtime="00:00:48.52" resultid="2307" heatid="7236" lane="7" entrytime="00:00:46.94" entrycourse="SCM" />
                <RESULT eventid="1092" points="83" swimtime="00:04:39.09" resultid="2308" heatid="7271" lane="8" entrytime="00:04:41.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.21" />
                    <SPLIT distance="100" swimtime="00:02:14.61" />
                    <SPLIT distance="150" swimtime="00:03:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="84" reactiontime="+98" swimtime="00:00:58.49" resultid="2309" heatid="7308" lane="8" entrytime="00:00:57.18" entrycourse="SCM" />
                <RESULT eventid="1336" points="38" swimtime="00:05:54.41" resultid="2310" heatid="7391" lane="3" entrytime="00:05:42.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.42" />
                    <SPLIT distance="100" swimtime="00:02:35.47" />
                    <SPLIT distance="150" swimtime="00:04:18.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="2311" heatid="7427" lane="9" entrytime="00:01:01.00" entrycourse="SCM" />
                <RESULT eventid="1465" points="84" reactiontime="+73" swimtime="00:02:05.35" resultid="2312" heatid="7453" lane="7" entrytime="00:02:07.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="2313" heatid="7507" lane="6" entrytime="00:02:21.30" entrycourse="SCM" />
                <RESULT eventid="1721" points="88" swimtime="00:08:44.15" resultid="2314" heatid="7571" lane="1" entrytime="00:08:40.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                    <SPLIT distance="100" swimtime="00:02:00.20" />
                    <SPLIT distance="150" swimtime="00:03:06.86" />
                    <SPLIT distance="200" swimtime="00:04:12.58" />
                    <SPLIT distance="250" swimtime="00:05:20.61" />
                    <SPLIT distance="300" swimtime="00:06:27.39" />
                    <SPLIT distance="350" swimtime="00:07:35.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="2297">
              <RESULTS>
                <RESULT eventid="1076" points="70" swimtime="00:00:48.93" resultid="2298" heatid="7248" lane="0" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="46" swimtime="00:05:04.81" resultid="2299" heatid="7277" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.67" />
                    <SPLIT distance="100" swimtime="00:02:26.40" />
                    <SPLIT distance="150" swimtime="00:03:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="68" reactiontime="+64" swimtime="00:00:54.28" resultid="2300" heatid="7317" lane="1" entrytime="00:00:58.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="58" reactiontime="+92" swimtime="00:01:55.66" resultid="2301" heatid="7350" lane="6" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="66" reactiontime="+75" swimtime="00:02:00.66" resultid="2302" heatid="7460" lane="3" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="52" swimtime="00:04:26.20" resultid="2303" heatid="7476" lane="9" entrytime="00:04:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="100" swimtime="00:02:02.62" />
                    <SPLIT distance="150" swimtime="00:03:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="67" reactiontime="+71" swimtime="00:04:19.12" resultid="2304" heatid="7530" lane="7" entrytime="00:04:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.62" />
                    <SPLIT distance="100" swimtime="00:02:08.26" />
                    <SPLIT distance="150" swimtime="00:03:15.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2305" heatid="7583" lane="4" entrytime="00:09:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="2528">
              <RESULTS>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="2529" heatid="7304" lane="4" entrytime="00:24:00.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="311" reactiontime="+80" swimtime="00:01:06.28" resultid="2530" heatid="7358" lane="0" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="292" reactiontime="+79" swimtime="00:00:32.76" resultid="2531" heatid="7442" lane="8" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="239" reactiontime="+81" swimtime="00:02:40.07" resultid="2532" heatid="7480" lane="0" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="197" reactiontime="+83" swimtime="00:01:22.55" resultid="2533" heatid="7516" lane="2" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" license="501806600051" athleteid="2270">
              <RESULTS>
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="2271" heatid="7328" lane="8" entrytime="00:04:23.00" entrycourse="SCM" />
                <RESULT eventid="1400" points="120" swimtime="00:02:06.21" resultid="2272" heatid="7408" lane="8" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="107" reactiontime="+67" swimtime="00:01:55.57" resultid="2273" heatid="7453" lane="6" entrytime="00:02:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="103" reactiontime="+85" swimtime="00:04:14.08" resultid="2274" heatid="7525" lane="0" entrytime="00:04:02.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.92" />
                    <SPLIT distance="100" swimtime="00:02:04.48" />
                    <SPLIT distance="150" swimtime="00:03:09.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="125" swimtime="00:00:57.09" resultid="2275" heatid="7538" lane="3" entrytime="00:00:56.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" license="501806700053" athleteid="2276">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2277" heatid="7276" lane="3" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2278" heatid="7377" lane="8" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="2279" heatid="7459" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Wisła 2" number="2">
              <RESULTS>
                <RESULT eventid="1391" points="135" reactiontime="+92" swimtime="00:02:55.97" resultid="2326" heatid="7403" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.94" />
                    <SPLIT distance="100" swimtime="00:01:57.41" />
                    <SPLIT distance="150" swimtime="00:02:26.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2241" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="2254" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="2280" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2288" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Wisła 3" number="3">
              <RESULTS>
                <RESULT eventid="1545" points="116" swimtime="00:02:47.30" resultid="2327" heatid="7493" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                    <SPLIT distance="100" swimtime="00:01:28.44" />
                    <SPLIT distance="150" swimtime="00:02:19.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2241" number="1" />
                    <RELAYPOSITION athleteid="2254" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2297" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2528" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" name="Wisła 1" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="82" swimtime="00:03:21.95" resultid="2325" heatid="7286" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                    <SPLIT distance="150" swimtime="00:02:32.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2241" number="1" />
                    <RELAYPOSITION athleteid="2261" number="2" reactiontime="+95" />
                    <RELAYPOSITION athleteid="2306" number="3" />
                    <RELAYPOSITION athleteid="2297" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Wisła 4" number="4">
              <RESULTS>
                <RESULT eventid="1705" status="DNS" swimtime="00:00:00.00" resultid="2328" heatid="7562" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2270" number="1" />
                    <RELAYPOSITION athleteid="2276" number="2" />
                    <RELAYPOSITION athleteid="2280" number="3" />
                    <RELAYPOSITION athleteid="2261" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAWRO" nation="POL" region="01" clubid="2062" name="Masters Wrocław">
          <CONTACT name="Krzekotowski" phone="693395453" />
          <ATHLETES>
            <ATHLETE birthdate="1976-05-09" firstname="Łukasz" gender="M" lastname="Amanowicz" nation="POL" athleteid="2489">
              <RESULTS>
                <RESULT eventid="1076" points="243" swimtime="00:00:32.45" resultid="2490" heatid="7251" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1288" points="167" reactiontime="+87" swimtime="00:01:21.48" resultid="2491" heatid="7351" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="139" reactiontime="+97" swimtime="00:01:47.25" resultid="2492" heatid="7416" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="161" reactiontime="+87" swimtime="00:00:46.34" resultid="2493" heatid="7548" lane="0" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="2394">
              <RESULTS>
                <RESULT eventid="1172" points="281" swimtime="00:23:22.81" resultid="2395" heatid="7300" lane="7" entrytime="00:23:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:28.31" />
                    <SPLIT distance="150" swimtime="00:02:14.93" />
                    <SPLIT distance="200" swimtime="00:03:01.39" />
                    <SPLIT distance="250" swimtime="00:03:47.98" />
                    <SPLIT distance="300" swimtime="00:04:35.25" />
                    <SPLIT distance="350" swimtime="00:05:22.12" />
                    <SPLIT distance="400" swimtime="00:06:09.19" />
                    <SPLIT distance="450" swimtime="00:06:55.81" />
                    <SPLIT distance="500" swimtime="00:07:42.87" />
                    <SPLIT distance="550" swimtime="00:08:29.87" />
                    <SPLIT distance="600" swimtime="00:09:17.05" />
                    <SPLIT distance="650" swimtime="00:10:03.91" />
                    <SPLIT distance="700" swimtime="00:10:50.91" />
                    <SPLIT distance="750" swimtime="00:11:38.42" />
                    <SPLIT distance="800" swimtime="00:12:25.44" />
                    <SPLIT distance="850" swimtime="00:13:13.16" />
                    <SPLIT distance="900" swimtime="00:14:01.01" />
                    <SPLIT distance="950" swimtime="00:14:48.05" />
                    <SPLIT distance="1000" swimtime="00:15:35.02" />
                    <SPLIT distance="1050" swimtime="00:16:21.93" />
                    <SPLIT distance="1100" swimtime="00:17:08.76" />
                    <SPLIT distance="1150" swimtime="00:17:55.53" />
                    <SPLIT distance="1200" swimtime="00:18:43.04" />
                    <SPLIT distance="1250" swimtime="00:19:30.81" />
                    <SPLIT distance="1300" swimtime="00:20:17.62" />
                    <SPLIT distance="1350" swimtime="00:21:04.26" />
                    <SPLIT distance="1400" swimtime="00:21:51.15" />
                    <SPLIT distance="1450" swimtime="00:22:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="191" swimtime="00:01:38.12" resultid="2396" heatid="7371" lane="9" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="200" swimtime="00:01:33.98" resultid="2397" heatid="7454" lane="5" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="245" swimtime="00:02:56.36" resultid="2398" heatid="7470" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:13.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="221" swimtime="00:03:17.20" resultid="2399" heatid="7526" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                    <SPLIT distance="150" swimtime="00:02:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="261" swimtime="00:06:05.80" resultid="2400" heatid="7569" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:28.23" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                    <SPLIT distance="200" swimtime="00:03:01.22" />
                    <SPLIT distance="250" swimtime="00:03:47.85" />
                    <SPLIT distance="300" swimtime="00:04:34.91" />
                    <SPLIT distance="350" swimtime="00:05:21.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="2078">
              <RESULTS>
                <RESULT eventid="1059" points="354" reactiontime="+74" swimtime="00:00:32.39" resultid="2079" heatid="7240" lane="5" entrytime="00:00:33.17" />
                <RESULT eventid="1092" points="270" reactiontime="+80" swimtime="00:03:08.33" resultid="2080" heatid="7273" lane="4" entrytime="00:03:04.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:02:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="272" reactiontime="+85" swimtime="00:00:39.61" resultid="2081" heatid="7311" lane="0" entrytime="00:00:39.50" />
                <RESULT eventid="1304" points="308" reactiontime="+78" swimtime="00:01:23.64" resultid="2082" heatid="7373" lane="9" entrytime="00:01:24.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="306" reactiontime="+80" swimtime="00:01:32.52" resultid="2083" heatid="7412" lane="9" entrytime="00:01:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="251" reactiontime="+87" swimtime="00:01:27.15" resultid="2084" heatid="7456" lane="2" entrytime="00:01:24.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="334" reactiontime="+72" swimtime="00:00:41.15" resultid="2085" heatid="7543" lane="8" entrytime="00:00:40.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="5886">
              <RESULTS>
                <RESULT eventid="1092" points="177" reactiontime="+85" swimtime="00:03:36.71" resultid="5887" heatid="7271" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="100" swimtime="00:01:47.09" />
                    <SPLIT distance="150" swimtime="00:02:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="189" swimtime="00:13:53.94" resultid="5888" heatid="7293" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:35.28" />
                    <SPLIT distance="150" swimtime="00:02:27.28" />
                    <SPLIT distance="200" swimtime="00:03:20.59" />
                    <SPLIT distance="250" swimtime="00:04:13.60" />
                    <SPLIT distance="300" swimtime="00:05:08.05" />
                    <SPLIT distance="350" swimtime="00:06:02.78" />
                    <SPLIT distance="400" swimtime="00:06:55.99" />
                    <SPLIT distance="450" swimtime="00:07:48.84" />
                    <SPLIT distance="500" swimtime="00:08:42.52" />
                    <SPLIT distance="550" swimtime="00:09:33.91" />
                    <SPLIT distance="600" swimtime="00:10:26.83" />
                    <SPLIT distance="650" swimtime="00:11:19.22" />
                    <SPLIT distance="700" swimtime="00:12:11.27" />
                    <SPLIT distance="750" swimtime="00:13:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="198" reactiontime="+67" swimtime="00:01:26.14" resultid="5889" heatid="7340" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="167" swimtime="00:01:42.49" resultid="5890" heatid="7368" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="143" reactiontime="+97" swimtime="00:01:45.10" resultid="5891" heatid="7452" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="182" swimtime="00:03:14.56" resultid="5892" heatid="7468" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                    <SPLIT distance="150" swimtime="00:02:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="153" reactiontime="+62" swimtime="00:03:42.68" resultid="5893" heatid="7523" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.15" />
                    <SPLIT distance="100" swimtime="00:01:50.07" />
                    <SPLIT distance="150" swimtime="00:02:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="199" swimtime="00:06:40.61" resultid="5894" heatid="7572" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:32.99" />
                    <SPLIT distance="150" swimtime="00:02:23.79" />
                    <SPLIT distance="200" swimtime="00:03:16.22" />
                    <SPLIT distance="250" swimtime="00:04:08.10" />
                    <SPLIT distance="300" swimtime="00:05:00.06" />
                    <SPLIT distance="350" swimtime="00:05:52.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-29" firstname="Piotr" gender="M" lastname="Krzekotowski" nation="POL" athleteid="2229">
              <RESULTS>
                <RESULT eventid="1076" points="148" reactiontime="+95" swimtime="00:00:38.23" resultid="2230" heatid="7251" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="1108" points="99" reactiontime="+96" swimtime="00:03:56.36" resultid="2231" heatid="7278" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.47" />
                    <SPLIT distance="100" swimtime="00:02:04.00" />
                    <SPLIT distance="150" swimtime="00:03:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="117" reactiontime="+93" swimtime="00:01:31.83" resultid="2232" heatid="7352" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="95" reactiontime="+89" swimtime="00:01:49.80" resultid="2233" heatid="7378" lane="6" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="118" reactiontime="+85" swimtime="00:01:53.09" resultid="2234" heatid="7417" lane="7" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="98" reactiontime="+94" swimtime="00:08:29.34" resultid="2235" heatid="8154" lane="4" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.82" />
                    <SPLIT distance="100" swimtime="00:02:08.38" />
                    <SPLIT distance="150" swimtime="00:03:25.69" />
                    <SPLIT distance="200" swimtime="00:04:38.22" />
                    <SPLIT distance="250" swimtime="00:05:40.67" />
                    <SPLIT distance="300" swimtime="00:06:43.19" />
                    <SPLIT distance="350" swimtime="00:07:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="114" reactiontime="+85" swimtime="00:00:51.94" resultid="2236" heatid="7549" lane="0" entrytime="00:00:48.00" />
                <RESULT eventid="1737" points="130" reactiontime="+87" swimtime="00:06:58.81" resultid="2237" heatid="7583" lane="5" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:41.31" />
                    <SPLIT distance="150" swimtime="00:02:35.23" />
                    <SPLIT distance="200" swimtime="00:03:28.52" />
                    <SPLIT distance="250" swimtime="00:04:21.33" />
                    <SPLIT distance="300" swimtime="00:05:14.69" />
                    <SPLIT distance="350" swimtime="00:06:07.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-10-24" firstname="Andrzej" gender="M" lastname="Marszałek" nation="POL" athleteid="2101">
              <RESULTS>
                <RESULT eventid="1076" points="107" reactiontime="+93" swimtime="00:00:42.64" resultid="2102" heatid="7249" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1156" points="108" reactiontime="+94" swimtime="00:15:29.01" resultid="2103" heatid="7299" lane="7" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:42.97" />
                    <SPLIT distance="150" swimtime="00:02:39.34" />
                    <SPLIT distance="200" swimtime="00:03:36.05" />
                    <SPLIT distance="250" swimtime="00:04:32.02" />
                    <SPLIT distance="300" swimtime="00:05:28.72" />
                    <SPLIT distance="350" swimtime="00:06:25.88" />
                    <SPLIT distance="400" swimtime="00:07:23.90" />
                    <SPLIT distance="450" swimtime="00:08:22.94" />
                    <SPLIT distance="500" swimtime="00:09:21.84" />
                    <SPLIT distance="550" swimtime="00:10:20.96" />
                    <SPLIT distance="600" swimtime="00:11:21.50" />
                    <SPLIT distance="650" swimtime="00:12:22.71" />
                    <SPLIT distance="700" swimtime="00:13:25.29" />
                    <SPLIT distance="750" swimtime="00:14:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="107" reactiontime="+94" swimtime="00:01:34.61" resultid="2104" heatid="7351" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="79" reactiontime="+92" swimtime="00:00:50.65" resultid="2105" heatid="7437" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1513" points="105" reactiontime="+92" swimtime="00:03:30.17" resultid="2106" heatid="7476" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                    <SPLIT distance="150" swimtime="00:02:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="104" reactiontime="+82" swimtime="00:07:29.93" resultid="2107" heatid="7583" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                    <SPLIT distance="100" swimtime="00:01:46.21" />
                    <SPLIT distance="150" swimtime="00:02:41.08" />
                    <SPLIT distance="200" swimtime="00:03:37.11" />
                    <SPLIT distance="250" swimtime="00:04:33.96" />
                    <SPLIT distance="300" swimtime="00:05:31.99" />
                    <SPLIT distance="350" swimtime="00:06:30.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-07-15" firstname="Alina" gender="F" lastname="Piekarska" nation="POL" athleteid="2061">
              <RESULTS>
                <RESULT eventid="1673" points="8" swimtime="00:02:17.95" resultid="2063" heatid="7537" lane="2" entrytime="00:02:09.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-04-26" firstname="Mateusz" gender="M" lastname="Pinkosz" nation="POL" athleteid="3820">
              <RESULTS>
                <RESULT eventid="1076" points="524" reactiontime="+70" swimtime="00:00:25.13" resultid="3821" heatid="7266" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="1156" points="467" reactiontime="+70" swimtime="00:09:31.51" resultid="3822" heatid="7294" lane="4" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:40.12" />
                    <SPLIT distance="200" swimtime="00:02:15.84" />
                    <SPLIT distance="250" swimtime="00:02:52.20" />
                    <SPLIT distance="300" swimtime="00:03:28.90" />
                    <SPLIT distance="350" swimtime="00:04:05.90" />
                    <SPLIT distance="400" swimtime="00:04:42.85" />
                    <SPLIT distance="450" swimtime="00:05:19.63" />
                    <SPLIT distance="500" swimtime="00:05:56.67" />
                    <SPLIT distance="550" swimtime="00:06:33.09" />
                    <SPLIT distance="600" swimtime="00:07:09.75" />
                    <SPLIT distance="650" swimtime="00:07:46.60" />
                    <SPLIT distance="700" swimtime="00:08:23.07" />
                    <SPLIT distance="750" swimtime="00:08:59.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="537" reactiontime="+65" swimtime="00:00:55.26" resultid="3823" heatid="7367" lane="6" entrytime="00:00:51.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="3824" heatid="7398" lane="0" entrytime="00:02:30.00" />
                <RESULT eventid="1449" points="492" reactiontime="+66" swimtime="00:00:27.55" resultid="3825" heatid="7451" lane="1" entrytime="00:00:25.82" />
                <RESULT eventid="1513" points="519" reactiontime="+66" swimtime="00:02:03.62" resultid="3826" heatid="7488" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="100" swimtime="00:00:58.30" />
                    <SPLIT distance="150" swimtime="00:01:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="3827" heatid="7517" lane="2" entrytime="00:01:02.00" />
                <RESULT eventid="1737" points="482" reactiontime="+64" swimtime="00:04:30.63" resultid="3828" heatid="7573" lane="4" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:01:02.15" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                    <SPLIT distance="200" swimtime="00:02:11.80" />
                    <SPLIT distance="250" swimtime="00:02:47.54" />
                    <SPLIT distance="300" swimtime="00:03:23.48" />
                    <SPLIT distance="350" swimtime="00:03:57.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAZDZ" nation="POL" region="11" clubid="5482" name="Masters Zdzieszowice">
          <CONTACT fax="masters.zdzieszowice" name="Jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-03" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="5507">
              <RESULTS>
                <RESULT eventid="1059" points="264" reactiontime="+72" swimtime="00:00:35.70" resultid="5508" heatid="7240" lane="9" entrytime="00:00:34.21" />
                <RESULT eventid="1092" points="255" reactiontime="+90" swimtime="00:03:12.11" resultid="5509" heatid="7273" lane="2" entrytime="00:03:10.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:34.64" />
                    <SPLIT distance="150" swimtime="00:02:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="285" reactiontime="+96" swimtime="00:03:24.41" resultid="5510" heatid="7329" lane="6" entrytime="00:03:42.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:40.75" />
                    <SPLIT distance="150" swimtime="00:02:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M3 - Pływak obrócił się na plecy w czasie wyścigu (z wyjątkiem wykonywania nawrotu, po dotknięciu dłońmi, a przed opuszczeniem ściany)." eventid="1336" reactiontime="+99" status="DSQ" swimtime="00:00:00.00" resultid="5511" heatid="7392" lane="5" entrytime="00:03:20.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="308" reactiontime="+87" swimtime="00:00:36.09" resultid="5512" heatid="7429" lane="4" entrytime="00:00:37.65" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="5513" heatid="7471" lane="8" entrytime="00:02:55.43" />
                <RESULT eventid="1608" points="238" reactiontime="+74" swimtime="00:01:28.04" resultid="5514" heatid="7510" lane="9" entrytime="00:01:25.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="286" reactiontime="+61" swimtime="00:00:43.30" resultid="5515" heatid="7541" lane="8" entrytime="00:00:45.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="5483">
              <RESULTS>
                <RESULT eventid="1256" points="411" reactiontime="+81" swimtime="00:02:41.59" resultid="5484" heatid="7332" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:01:59.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="368" reactiontime="+83" swimtime="00:02:30.91" resultid="5485" heatid="7394" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="5486" heatid="7459" lane="0" />
                <RESULT eventid="1577" status="WDR" swimtime="00:00:00.00" resultid="5487" heatid="8152" lane="3" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="5488" heatid="7512" lane="7" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5489" heatid="7529" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-06" firstname="Paulina" gender="F" lastname="Kawecka" nation="POL" athleteid="5495">
              <RESULTS>
                <RESULT eventid="1433" points="270" swimtime="00:00:37.69" resultid="5496" heatid="7429" lane="5" entrytime="00:00:37.85" />
                <RESULT eventid="1465" points="261" swimtime="00:01:26.05" resultid="5497" heatid="7456" lane="0" entrytime="00:01:26.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="214" swimtime="00:01:31.25" resultid="5498" heatid="7509" lane="2" entrytime="00:01:30.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="269" swimtime="00:03:04.58" resultid="5499" heatid="7526" lane="7" entrytime="00:03:15.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-09" firstname="Daria" gender="F" lastname="Szydłowska - Smętek" nation="POL" athleteid="5500">
              <RESULTS>
                <RESULT eventid="1092" points="370" reactiontime="+85" swimtime="00:02:49.60" resultid="5501" heatid="7274" lane="7" entrytime="00:02:55.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:10.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="396" reactiontime="+97" swimtime="00:10:52.44" resultid="5502" heatid="7291" lane="1" entrytime="00:12:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:02:36.55" />
                    <SPLIT distance="250" swimtime="00:03:17.97" />
                    <SPLIT distance="300" swimtime="00:03:59.44" />
                    <SPLIT distance="350" swimtime="00:04:41.35" />
                    <SPLIT distance="400" swimtime="00:05:23.00" />
                    <SPLIT distance="450" swimtime="00:06:04.58" />
                    <SPLIT distance="500" swimtime="00:06:46.25" />
                    <SPLIT distance="550" swimtime="00:07:28.03" />
                    <SPLIT distance="600" swimtime="00:08:10.05" />
                    <SPLIT distance="650" swimtime="00:08:51.55" />
                    <SPLIT distance="700" swimtime="00:09:32.69" />
                    <SPLIT distance="750" swimtime="00:10:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="308" reactiontime="+74" swimtime="00:00:37.99" resultid="5503" heatid="7311" lane="1" entrytime="00:00:39.25" />
                <RESULT eventid="1272" points="392" reactiontime="+80" swimtime="00:01:08.61" resultid="5504" heatid="7346" lane="9" entrytime="00:01:10.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="373" reactiontime="+85" swimtime="00:02:33.34" resultid="5505" heatid="7473" lane="0" entrytime="00:02:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="318" reactiontime="+96" swimtime="00:06:18.97" resultid="5506" heatid="8149" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:02:20.20" />
                    <SPLIT distance="200" swimtime="00:03:09.29" />
                    <SPLIT distance="250" swimtime="00:04:02.38" />
                    <SPLIT distance="300" swimtime="00:04:55.21" />
                    <SPLIT distance="350" swimtime="00:05:37.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-03" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="5490">
              <RESULTS>
                <RESULT eventid="1304" points="300" swimtime="00:01:24.41" resultid="5491" heatid="7373" lane="0" entrytime="00:01:24.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="224" reactiontime="+99" swimtime="00:03:16.85" resultid="5492" heatid="7393" lane="0" entrytime="00:03:14.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:34.98" />
                    <SPLIT distance="150" swimtime="00:02:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="282" reactiontime="+97" swimtime="00:00:37.17" resultid="5493" heatid="7429" lane="6" entrytime="00:00:38.75" />
                <RESULT eventid="1561" points="271" swimtime="00:06:39.96" resultid="5494" heatid="8151" lane="0" entrytime="00:06:29.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="150" swimtime="00:02:27.99" />
                    <SPLIT distance="200" swimtime="00:03:18.00" />
                    <SPLIT distance="250" swimtime="00:04:15.36" />
                    <SPLIT distance="300" swimtime="00:05:12.02" />
                    <SPLIT distance="350" swimtime="00:05:57.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" status="WDR" swimtime="00:00:00.00" resultid="5516" heatid="7490" lane="2" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5490" number="1" />
                    <RELAYPOSITION athleteid="5507" number="2" />
                    <RELAYPOSITION athleteid="5495" number="3" />
                    <RELAYPOSITION athleteid="5500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" status="WDR" swimtime="00:00:00.00" resultid="5517" heatid="7399" lane="6" entrytime="00:02:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5490" number="1" />
                    <RELAYPOSITION athleteid="5507" number="2" />
                    <RELAYPOSITION athleteid="5495" number="3" />
                    <RELAYPOSITION athleteid="5500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03605" nation="POL" region="05" clubid="4926" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1982-01-01" firstname="Łukasz" gender="M" lastname="Bogusiak" nation="POL" athleteid="6862">
              <RESULTS>
                <RESULT eventid="1076" points="189" swimtime="00:00:35.26" resultid="6863" heatid="7251" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1288" points="164" reactiontime="+85" swimtime="00:01:22.08" resultid="6864" heatid="7352" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach. (Time: 12:19)" eventid="1320" status="DSQ" swimtime="00:01:39.18" resultid="6865" heatid="7379" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6866" heatid="7436" lane="9" />
                <RESULT eventid="1513" points="127" reactiontime="+88" swimtime="00:03:17.28" resultid="6867" heatid="7477" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:24.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" license="503605700020" athleteid="4958">
              <RESULTS>
                <RESULT eventid="1076" points="426" reactiontime="+72" swimtime="00:00:26.91" resultid="4959" heatid="7261" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4960" heatid="7362" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1320" points="395" reactiontime="+81" swimtime="00:01:08.49" resultid="4961" heatid="7386" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="386" reactiontime="+82" swimtime="00:00:29.87" resultid="4962" heatid="7445" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1689" points="362" reactiontime="+78" swimtime="00:00:35.41" resultid="4963" heatid="7554" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-10-05" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" license="503605700014" athleteid="5022">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5023" heatid="7281" lane="2" entrytime="00:02:47.17" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5025" heatid="7357" lane="5" entrytime="00:01:07.17" />
                <RESULT eventid="1320" points="289" reactiontime="+88" swimtime="00:01:15.99" resultid="5026" heatid="7383" lane="1" entrytime="00:01:17.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="309" reactiontime="+82" swimtime="00:00:32.14" resultid="5027" heatid="7441" lane="7" entrytime="00:00:33.77" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5028" heatid="7482" lane="3" entrytime="00:02:27.17" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="5029" heatid="7517" lane="0" entrytime="00:01:17.17" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5030" heatid="7579" lane="8" entrytime="00:05:47.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-14" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" license="503605700017" athleteid="5050">
              <RESULTS>
                <RESULT eventid="1076" points="259" swimtime="00:00:31.77" resultid="5051" heatid="7257" lane="0" entrytime="00:00:30.90" />
                <RESULT eventid="1417" points="241" reactiontime="+87" swimtime="00:01:29.24" resultid="5052" heatid="7418" lane="4" entrytime="00:01:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="273" reactiontime="+84" swimtime="00:00:38.89" resultid="5053" heatid="7552" lane="1" entrytime="00:00:40.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-01" firstname="Marek" gender="M" lastname="Gurbski" nation="POL" license="503605700019" athleteid="5012">
              <RESULTS>
                <RESULT eventid="1076" points="347" swimtime="00:00:28.83" resultid="5013" heatid="7257" lane="8" entrytime="00:00:30.36" />
                <RESULT eventid="1224" points="276" reactiontime="+68" swimtime="00:00:34.10" resultid="5014" heatid="7321" lane="5" entrytime="00:00:36.02" />
                <RESULT eventid="1320" points="324" swimtime="00:01:13.17" resultid="5015" heatid="7382" lane="2" entrytime="00:01:19.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="327" reactiontime="+72" swimtime="00:00:31.54" resultid="5016" heatid="7441" lane="6" entrytime="00:00:33.34" />
                <RESULT eventid="1689" points="308" reactiontime="+86" swimtime="00:00:37.37" resultid="5017" heatid="7552" lane="7" entrytime="00:00:40.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-06-09" firstname="Michał" gender="M" lastname="Gurbski" nation="POL" license="503605700026" athleteid="5037">
              <RESULTS>
                <RESULT eventid="1076" points="306" reactiontime="+94" swimtime="00:00:30.06" resultid="5038" heatid="7256" lane="2" entrytime="00:00:31.36" />
                <RESULT eventid="1224" points="236" reactiontime="+89" swimtime="00:00:35.92" resultid="5039" heatid="7321" lane="1" entrytime="00:00:37.02" />
                <RESULT eventid="1320" points="246" reactiontime="+93" swimtime="00:01:20.14" resultid="5040" heatid="7381" lane="3" entrytime="00:01:20.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="241" reactiontime="+91" swimtime="00:00:34.93" resultid="5041" heatid="7440" lane="4" entrytime="00:00:34.34" />
                <RESULT eventid="1689" points="245" reactiontime="+88" swimtime="00:00:40.32" resultid="5042" heatid="7551" lane="5" entrytime="00:00:41.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-01" firstname="Paulina" gender="F" lastname="Kaczmarek" nation="POL" license="503605600032" athleteid="5000">
              <RESULTS>
                <RESULT eventid="1207" points="337" reactiontime="+71" swimtime="00:00:36.88" resultid="5001" heatid="7313" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1465" points="291" reactiontime="+77" swimtime="00:01:22.95" resultid="5002" heatid="7457" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" license="103605700004" athleteid="4964">
              <RESULTS>
                <RESULT eventid="1076" points="320" swimtime="00:00:29.61" resultid="4965" heatid="7249" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1108" points="225" swimtime="00:03:00.24" resultid="4966" heatid="7279" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="217" reactiontime="+62" swimtime="00:03:19.94" resultid="4967" heatid="7335" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:34.78" />
                    <SPLIT distance="150" swimtime="00:02:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="256" swimtime="00:01:19.14" resultid="4968" heatid="7380" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="251" reactiontime="+99" swimtime="00:01:28.08" resultid="4969" heatid="7417" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="161" swimtime="00:07:12.12" resultid="4971" heatid="8153" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:27.61" />
                    <SPLIT distance="200" swimtime="00:03:23.84" />
                    <SPLIT distance="250" swimtime="00:04:27.64" />
                    <SPLIT distance="300" swimtime="00:05:32.47" />
                    <SPLIT distance="350" swimtime="00:06:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="200" reactiontime="+78" swimtime="00:03:00.40" resultid="4972" heatid="7531" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:24.31" />
                    <SPLIT distance="150" swimtime="00:02:12.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="286" reactiontime="+99" swimtime="00:00:38.32" resultid="4973" heatid="7551" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-14" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" license="503605700018" athleteid="5003">
              <RESULTS>
                <RESULT eventid="1224" points="231" reactiontime="+68" swimtime="00:00:36.17" resultid="5004" heatid="7322" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-03-07" firstname="Julia" gender="F" lastname="Kałczak" nation="POL" license="503605600021" athleteid="4950">
              <RESULTS>
                <RESULT eventid="1092" points="399" reactiontime="+90" swimtime="00:02:45.47" resultid="4951" heatid="7274" lane="2" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:02:05.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="384" reactiontime="+66" swimtime="00:00:35.29" resultid="4952" heatid="7312" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1304" points="409" reactiontime="+85" swimtime="00:01:16.09" resultid="4953" heatid="7374" lane="8" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="4954" heatid="7433" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1465" points="362" reactiontime="+73" swimtime="00:01:17.21" resultid="4955" heatid="7457" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="419" reactiontime="+82" swimtime="00:01:12.96" resultid="4956" heatid="7510" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="326" reactiontime="+90" swimtime="00:00:41.47" resultid="4957" heatid="7543" lane="0" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-06" firstname="Monika" gender="F" lastname="Klarecka" nation="POL" license="503605600029" athleteid="4974">
              <RESULTS>
                <RESULT eventid="1092" points="151" reactiontime="+77" swimtime="00:03:48.82" resultid="4975" heatid="7271" lane="4" entrytime="00:03:55.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:54.77" />
                    <SPLIT distance="150" swimtime="00:02:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="153" reactiontime="+75" swimtime="00:14:55.67" resultid="4976" heatid="7292" lane="5" entrytime="00:13:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:41.20" />
                    <SPLIT distance="150" swimtime="00:02:37.30" />
                    <SPLIT distance="200" swimtime="00:03:34.59" />
                    <SPLIT distance="250" swimtime="00:04:30.92" />
                    <SPLIT distance="300" swimtime="00:05:27.73" />
                    <SPLIT distance="350" swimtime="00:06:24.88" />
                    <SPLIT distance="400" swimtime="00:07:22.62" />
                    <SPLIT distance="450" swimtime="00:08:20.67" />
                    <SPLIT distance="500" swimtime="00:09:18.67" />
                    <SPLIT distance="550" swimtime="00:10:16.84" />
                    <SPLIT distance="600" swimtime="00:11:13.89" />
                    <SPLIT distance="650" swimtime="00:12:10.70" />
                    <SPLIT distance="700" swimtime="00:13:07.56" />
                    <SPLIT distance="750" swimtime="00:14:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="189" reactiontime="+83" swimtime="00:03:54.35" resultid="4977" heatid="7328" lane="6" entrytime="00:04:03.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.32" />
                    <SPLIT distance="100" swimtime="00:01:55.89" />
                    <SPLIT distance="150" swimtime="00:02:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="122" reactiontime="+85" swimtime="00:04:00.52" resultid="4978" heatid="7392" lane="0" entrytime="00:04:14.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="100" swimtime="00:01:53.83" />
                    <SPLIT distance="150" swimtime="00:02:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="144" reactiontime="+93" swimtime="00:00:46.42" resultid="4979" heatid="7427" lane="5" entrytime="00:00:49.87" />
                <RESULT eventid="1561" points="143" reactiontime="+83" swimtime="00:08:14.68" resultid="4980" heatid="8149" lane="2" entrytime="00:08:20.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                    <SPLIT distance="100" swimtime="00:01:55.26" />
                    <SPLIT distance="150" swimtime="00:03:06.71" />
                    <SPLIT distance="200" swimtime="00:04:18.35" />
                    <SPLIT distance="250" swimtime="00:05:23.77" />
                    <SPLIT distance="300" swimtime="00:06:26.26" />
                    <SPLIT distance="350" swimtime="00:07:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="88" swimtime="00:04:27.35" resultid="4981" heatid="7525" lane="9" entrytime="00:04:27.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.58" />
                    <SPLIT distance="100" swimtime="00:02:15.94" />
                    <SPLIT distance="150" swimtime="00:03:22.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="164" reactiontime="+89" swimtime="00:07:07.23" resultid="4982" heatid="7570" lane="8" entrytime="00:07:25.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:42.82" />
                    <SPLIT distance="150" swimtime="00:02:37.59" />
                    <SPLIT distance="200" swimtime="00:03:32.88" />
                    <SPLIT distance="250" swimtime="00:04:26.59" />
                    <SPLIT distance="300" swimtime="00:05:22.28" />
                    <SPLIT distance="350" swimtime="00:06:16.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-01" firstname="Mateusz" gender="M" lastname="Klonowski" nation="POL" license="503605700033" athleteid="5054">
              <RESULTS>
                <RESULT eventid="1417" points="338" reactiontime="+84" swimtime="00:01:19.76" resultid="5055" heatid="7419" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="372" reactiontime="+75" swimtime="00:00:35.08" resultid="5056" heatid="7555" lane="4" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-30" firstname="Monika" gender="F" lastname="Kurstak-Jagiełło" nation="POL" license="503605600022" athleteid="4945">
              <RESULTS>
                <RESULT eventid="1059" points="411" reactiontime="+89" swimtime="00:00:30.84" resultid="4946" heatid="7243" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1207" points="280" reactiontime="+76" swimtime="00:00:39.21" resultid="4947" heatid="7311" lane="2" entrytime="00:00:38.50" />
                <RESULT eventid="1272" points="392" reactiontime="+87" swimtime="00:01:08.64" resultid="4948" heatid="7345" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="283" reactiontime="+76" swimtime="00:00:43.46" resultid="4949" heatid="7541" lane="5" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-18" firstname="Paweł" gender="M" lastname="Lipka" nation="POL" license="503605700025" athleteid="4941">
              <RESULTS>
                <RESULT eventid="1320" points="197" reactiontime="+88" swimtime="00:01:26.37" resultid="4942" heatid="7380" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="201" reactiontime="+85" swimtime="00:00:37.07" resultid="4943" heatid="7438" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1625" points="117" reactiontime="+89" swimtime="00:01:38.14" resultid="4944" heatid="7515" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-03-04" firstname="Maciej" gender="M" lastname="Machnicki" nation="POL" license="503605700030" athleteid="4998">
              <RESULTS>
                <RESULT eventid="1076" points="254" reactiontime="+90" swimtime="00:00:31.97" resultid="4999" heatid="7254" lane="9" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-12" firstname="Magdalena" gender="F" lastname="Maciąg" nation="POL" license="503605600031" athleteid="5018">
              <RESULTS>
                <RESULT eventid="1059" points="344" swimtime="00:00:32.71" resultid="5019" heatid="7239" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1272" points="333" reactiontime="+92" swimtime="00:01:12.47" resultid="5020" heatid="7343" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="305" reactiontime="+85" swimtime="00:01:23.86" resultid="5021" heatid="7370" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-11" firstname="Przemysław" gender="M" lastname="Michniewski" nation="POL" license="503605700012" athleteid="5043">
              <RESULTS>
                <RESULT eventid="1076" points="486" swimtime="00:00:25.76" resultid="5044" heatid="7266" lane="0" entrytime="00:00:26.50" />
                <RESULT eventid="1256" points="419" reactiontime="+79" swimtime="00:02:40.50" resultid="5045" heatid="7338" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                    <SPLIT distance="150" swimtime="00:01:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="468" reactiontime="+84" swimtime="00:01:04.70" resultid="5046" heatid="7388" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="478" reactiontime="+84" swimtime="00:01:11.08" resultid="5047" heatid="7424" lane="2" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="425" reactiontime="+77" swimtime="00:00:28.91" resultid="5048" heatid="7448" lane="9" entrytime="00:00:28.80" />
                <RESULT eventid="1689" points="469" reactiontime="+78" swimtime="00:00:32.48" resultid="5049" heatid="7560" lane="7" entrytime="00:00:32.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" license="503605700007" athleteid="4927">
              <RESULTS>
                <RESULT eventid="1076" points="508" reactiontime="+72" swimtime="00:00:25.38" resultid="4928" heatid="7266" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1288" points="508" reactiontime="+79" swimtime="00:00:56.29" resultid="4929" heatid="7363" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="344" reactiontime="+88" swimtime="00:02:34.44" resultid="4930" heatid="7397" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="480" reactiontime="+70" swimtime="00:00:27.77" resultid="4931" heatid="7447" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1513" points="408" reactiontime="+73" swimtime="00:02:13.90" resultid="4932" heatid="7483" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="458" reactiontime="+69" swimtime="00:01:02.33" resultid="4933" heatid="7519" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" license="503605700011" athleteid="5005">
              <RESULTS>
                <RESULT eventid="1188" points="316" reactiontime="+92" swimtime="00:20:43.84" resultid="5006" heatid="7303" lane="2" entrytime="00:21:57.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:50.02" />
                    <SPLIT distance="200" swimtime="00:02:29.73" />
                    <SPLIT distance="250" swimtime="00:03:10.34" />
                    <SPLIT distance="300" swimtime="00:03:51.48" />
                    <SPLIT distance="350" swimtime="00:04:33.09" />
                    <SPLIT distance="400" swimtime="00:05:15.03" />
                    <SPLIT distance="450" swimtime="00:05:57.10" />
                    <SPLIT distance="500" swimtime="00:06:39.71" />
                    <SPLIT distance="550" swimtime="00:07:22.28" />
                    <SPLIT distance="600" swimtime="00:08:04.79" />
                    <SPLIT distance="650" swimtime="00:08:48.16" />
                    <SPLIT distance="700" swimtime="00:09:31.60" />
                    <SPLIT distance="750" swimtime="00:10:14.01" />
                    <SPLIT distance="800" swimtime="00:10:56.43" />
                    <SPLIT distance="850" swimtime="00:11:38.48" />
                    <SPLIT distance="900" swimtime="00:12:21.11" />
                    <SPLIT distance="950" swimtime="00:13:04.06" />
                    <SPLIT distance="1000" swimtime="00:13:46.64" />
                    <SPLIT distance="1050" swimtime="00:14:29.14" />
                    <SPLIT distance="1100" swimtime="00:15:11.61" />
                    <SPLIT distance="1150" swimtime="00:15:53.31" />
                    <SPLIT distance="1200" swimtime="00:16:34.31" />
                    <SPLIT distance="1250" swimtime="00:17:16.75" />
                    <SPLIT distance="1300" swimtime="00:17:58.80" />
                    <SPLIT distance="1350" swimtime="00:18:41.34" />
                    <SPLIT distance="1400" swimtime="00:19:23.81" />
                    <SPLIT distance="1450" swimtime="00:20:06.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="5007" heatid="7322" lane="5" entrytime="00:00:34.44" />
                <RESULT eventid="1288" points="398" reactiontime="+81" swimtime="00:01:01.08" resultid="5008" heatid="7357" lane="3" entrytime="00:01:07.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="351" reactiontime="+79" swimtime="00:00:30.82" resultid="5009" heatid="7445" lane="5" entrytime="00:00:29.99" />
                <RESULT eventid="1513" points="363" reactiontime="+92" swimtime="00:02:19.24" resultid="5010" heatid="7482" lane="6" entrytime="00:02:27.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="306" reactiontime="+95" swimtime="00:05:14.79" resultid="5011" heatid="7577" lane="1" entrytime="00:05:17.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:49.18" />
                    <SPLIT distance="200" swimtime="00:02:27.75" />
                    <SPLIT distance="250" swimtime="00:03:07.20" />
                    <SPLIT distance="300" swimtime="00:03:48.79" />
                    <SPLIT distance="350" swimtime="00:04:32.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-14" firstname="Anna" gender="F" lastname="Ostrowska" nation="POL" license="103605600003" athleteid="4986">
              <RESULTS>
                <RESULT eventid="1059" points="386" reactiontime="+96" swimtime="00:00:31.49" resultid="4987" heatid="7241" lane="6" entrytime="00:00:32.20" />
                <RESULT eventid="1433" points="313" reactiontime="+91" swimtime="00:00:35.88" resultid="4988" heatid="7430" lane="0" entrytime="00:00:37.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" license="503605700016" athleteid="4983">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4984" heatid="7253" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1689" points="232" reactiontime="+87" swimtime="00:00:41.06" resultid="4985" heatid="7551" lane="9" entrytime="00:00:42.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-04" firstname="Jakub" gender="M" lastname="Sidorowicz" nation="POL" license="503605700023" athleteid="5031">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5032" heatid="7280" lane="1" entrytime="00:03:09.99" />
                <RESULT eventid="1256" points="195" reactiontime="+94" swimtime="00:03:27.10" resultid="5033" heatid="7336" lane="8" entrytime="00:03:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:36.17" />
                    <SPLIT distance="150" swimtime="00:02:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="173" reactiontime="+97" swimtime="00:01:30.14" resultid="5034" heatid="7383" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="209" reactiontime="+84" swimtime="00:01:33.70" resultid="5035" heatid="7419" lane="4" entrytime="00:01:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="222" reactiontime="+92" swimtime="00:00:41.67" resultid="5036" heatid="7553" lane="0" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" license="503605700001" athleteid="4934">
              <RESULTS>
                <RESULT eventid="1320" points="329" reactiontime="+82" swimtime="00:01:12.80" resultid="4935" heatid="7385" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="348" reactiontime="+80" swimtime="00:01:19.04" resultid="4936" heatid="7423" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="384" reactiontime="+83" swimtime="00:00:34.71" resultid="4937" heatid="7558" lane="0" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-02" firstname="Ksawery" gender="M" lastname="Wiaderek" nation="POL" license="103605700005" athleteid="4993">
              <RESULTS>
                <RESULT eventid="1076" points="410" swimtime="00:00:27.26" resultid="4994" heatid="7263" lane="0" entrytime="00:00:27.50" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="4995" heatid="7322" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4996" heatid="7362" lane="8" entrytime="00:01:01.00" />
                <RESULT eventid="1449" points="383" reactiontime="+77" swimtime="00:00:29.94" resultid="4997" heatid="7448" lane="8" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Joanna" gender="F" lastname="Wilińska-Nowak" nation="POL" license="103605600002" athleteid="4938">
              <RESULTS>
                <RESULT eventid="1336" points="373" reactiontime="+98" swimtime="00:02:46.07" resultid="4939" heatid="7393" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="441" reactiontime="+91" swimtime="00:01:11.73" resultid="4940" heatid="7511" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" license="503605700010" athleteid="4989">
              <RESULTS>
                <RESULT eventid="1076" points="402" reactiontime="+81" swimtime="00:00:27.43" resultid="4990" heatid="7259" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1449" points="329" reactiontime="+78" swimtime="00:00:31.49" resultid="4991" heatid="7442" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1689" points="371" reactiontime="+81" swimtime="00:00:35.14" resultid="4992" heatid="7557" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1545" points="314" reactiontime="+83" swimtime="00:02:00.31" resultid="5063" heatid="7494" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                    <SPLIT distance="150" swimtime="00:01:27.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5005" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="5050" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4998" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4941" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1545" points="368" reactiontime="+89" swimtime="00:01:54.13" resultid="5064" heatid="7494" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                    <SPLIT distance="150" swimtime="00:01:26.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5037" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="5003" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4983" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="5012" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="1545" points="457" reactiontime="+82" swimtime="00:01:46.17" resultid="5065" heatid="7495" lane="5" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                    <SPLIT distance="100" swimtime="00:00:53.57" />
                    <SPLIT distance="150" swimtime="00:01:19.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4958" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5022" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4927" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="4989" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="1545" status="WDR" swimtime="00:00:00.00" resultid="5066" heatid="7495" lane="7" entrytime="00:01:49.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5043" number="1" />
                    <RELAYPOSITION athleteid="4964" number="2" />
                    <RELAYPOSITION athleteid="4934" number="3" />
                    <RELAYPOSITION athleteid="4993" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="11">
              <RESULTS>
                <RESULT eventid="1391" points="388" reactiontime="+75" swimtime="00:02:03.99" resultid="5067" heatid="7406" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:37.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5022" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4934" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4927" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4958" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="12">
              <RESULTS>
                <RESULT eventid="1391" points="301" swimtime="00:02:14.83" resultid="5068" heatid="7405" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:47.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4964" number="1" />
                    <RELAYPOSITION athleteid="5050" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="4989" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="5005" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="13">
              <RESULTS>
                <RESULT eventid="1391" points="362" reactiontime="+70" swimtime="00:02:06.89" resultid="5069" heatid="7405" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:38.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5003" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5043" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4993" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5012" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="14">
              <RESULTS>
                <RESULT eventid="1391" points="252" reactiontime="+87" swimtime="00:02:23.05" resultid="5070" heatid="7404" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:01:53.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5037" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="4983" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4941" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4998" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="1368" points="301" reactiontime="+73" swimtime="00:02:32.75" resultid="5061" heatid="7401" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="150" swimtime="00:02:01.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5000" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4974" number="2" />
                    <RELAYPOSITION athleteid="4950" number="3" />
                    <RELAYPOSITION athleteid="4986" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="6">
              <RESULTS>
                <RESULT eventid="1529" points="374" swimtime="00:02:10.34" resultid="5062" heatid="7491" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:38.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5000" number="1" />
                    <RELAYPOSITION athleteid="4950" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5018" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4986" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="467" reactiontime="+84" swimtime="00:01:53.28" resultid="5059" heatid="7289" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:00:57.03" />
                    <SPLIT distance="150" swimtime="00:01:27.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4986" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="5005" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4945" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4927" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="329" swimtime="00:02:07.23" resultid="5058" heatid="7289" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:36.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4958" number="1" />
                    <RELAYPOSITION athleteid="4974" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="5012" number="3" />
                    <RELAYPOSITION athleteid="4950" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1124" points="404" swimtime="00:01:58.84" resultid="5057" heatid="7288" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                    <SPLIT distance="150" swimtime="00:01:31.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5000" number="1" />
                    <RELAYPOSITION athleteid="4993" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="5018" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4989" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1705" points="361" reactiontime="+84" swimtime="00:02:15.34" resultid="5060" heatid="7564" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:20.94" />
                    <SPLIT distance="150" swimtime="00:01:48.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4986" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4950" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4927" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="4958" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="15">
              <RESULTS>
                <RESULT eventid="1705" points="275" reactiontime="+65" swimtime="00:02:28.17" resultid="5071" heatid="7564" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:55.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5003" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4934" number="2" reactiontime="+10" />
                    <RELAYPOSITION athleteid="4974" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5018" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00116" nation="POL" region="16" clubid="2552" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="4459">
              <RESULTS>
                <RESULT eventid="1076" points="188" reactiontime="+94" swimtime="00:00:35.35" resultid="4460" heatid="7251" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="2559">
              <RESULTS>
                <RESULT eventid="1108" points="156" reactiontime="+83" swimtime="00:03:23.47" resultid="2560" heatid="7279" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                    <SPLIT distance="150" swimtime="00:02:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="173" reactiontime="+83" swimtime="00:03:35.26" resultid="2561" heatid="7334" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:43.45" />
                    <SPLIT distance="150" swimtime="00:02:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="198" reactiontime="+81" swimtime="00:01:35.35" resultid="2562" heatid="7415" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="176" reactiontime="+80" swimtime="00:00:38.75" resultid="2563" heatid="7439" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1689" points="227" reactiontime="+76" swimtime="00:00:41.39" resultid="2564" heatid="7550" lane="5" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="2583">
              <RESULTS>
                <RESULT eventid="1156" points="356" swimtime="00:10:25.10" resultid="2584" heatid="7294" lane="3" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:46.82" />
                    <SPLIT distance="200" swimtime="00:02:24.65" />
                    <SPLIT distance="250" swimtime="00:03:03.09" />
                    <SPLIT distance="300" swimtime="00:03:41.92" />
                    <SPLIT distance="350" swimtime="00:04:21.39" />
                    <SPLIT distance="400" swimtime="00:05:01.06" />
                    <SPLIT distance="450" swimtime="00:05:41.18" />
                    <SPLIT distance="500" swimtime="00:06:21.31" />
                    <SPLIT distance="550" swimtime="00:07:01.55" />
                    <SPLIT distance="600" swimtime="00:07:42.12" />
                    <SPLIT distance="650" swimtime="00:08:23.45" />
                    <SPLIT distance="700" swimtime="00:09:04.31" />
                    <SPLIT distance="750" swimtime="00:09:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="247" reactiontime="+95" swimtime="00:02:52.29" resultid="2585" heatid="7397" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:07.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="352" reactiontime="+93" swimtime="00:05:33.36" resultid="2586" heatid="8157" lane="4" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:01:58.13" />
                    <SPLIT distance="200" swimtime="00:02:41.42" />
                    <SPLIT distance="250" swimtime="00:03:29.47" />
                    <SPLIT distance="300" swimtime="00:04:18.42" />
                    <SPLIT distance="350" swimtime="00:04:56.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="353" swimtime="00:05:00.18" resultid="2587" heatid="7574" lane="0" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:44.70" />
                    <SPLIT distance="200" swimtime="00:02:22.92" />
                    <SPLIT distance="250" swimtime="00:03:02.13" />
                    <SPLIT distance="300" swimtime="00:03:41.63" />
                    <SPLIT distance="350" swimtime="00:04:21.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="2574">
              <RESULTS>
                <RESULT eventid="1240" points="48" swimtime="00:06:08.53" resultid="2575" heatid="7327" lane="3" entrytime="00:05:04.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.50" />
                    <SPLIT distance="100" swimtime="00:02:59.23" />
                    <SPLIT distance="150" swimtime="00:04:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="47" swimtime="00:02:52.21" resultid="2576" heatid="7408" lane="9" entrytime="00:02:27.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="44" swimtime="00:01:20.62" resultid="2577" heatid="7537" lane="5" entrytime="00:01:07.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Piotr" gender="M" lastname="Orłowski" nation="POL" athleteid="2578">
              <RESULTS>
                <RESULT eventid="1076" points="574" reactiontime="+74" swimtime="00:00:24.37" resultid="2579" heatid="7270" lane="2" entrytime="00:00:23.50" />
                <RESULT eventid="1288" points="583" reactiontime="+76" swimtime="00:00:53.78" resultid="2580" heatid="7367" lane="7" entrytime="00:00:53.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="555" reactiontime="+79" swimtime="00:00:26.46" resultid="2581" heatid="7451" lane="8" entrytime="00:00:25.84" />
                <RESULT eventid="1625" points="562" reactiontime="+76" swimtime="00:00:58.25" resultid="2582" heatid="7522" lane="7" entrytime="00:00:56.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="2553">
              <RESULTS>
                <RESULT eventid="1140" points="419" reactiontime="+72" swimtime="00:10:40.11" resultid="2554" heatid="7290" lane="2" entrytime="00:10:32.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:54.25" />
                    <SPLIT distance="200" swimtime="00:02:34.53" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:55.27" />
                    <SPLIT distance="350" swimtime="00:04:35.53" />
                    <SPLIT distance="400" swimtime="00:05:15.93" />
                    <SPLIT distance="450" swimtime="00:05:56.40" />
                    <SPLIT distance="500" swimtime="00:06:36.72" />
                    <SPLIT distance="550" swimtime="00:07:17.30" />
                    <SPLIT distance="600" swimtime="00:07:57.81" />
                    <SPLIT distance="650" swimtime="00:08:38.71" />
                    <SPLIT distance="700" swimtime="00:09:19.59" />
                    <SPLIT distance="750" swimtime="00:10:00.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="393" reactiontime="+71" swimtime="00:01:08.60" resultid="2555" heatid="7346" lane="7" entrytime="00:01:09.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="422" reactiontime="+73" swimtime="00:02:27.14" resultid="2556" heatid="7473" lane="3" entrytime="00:02:27.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="303" reactiontime="+87" swimtime="00:02:57.51" resultid="2557" heatid="7527" lane="2" entrytime="00:02:55.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:13.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="422" reactiontime="+75" swimtime="00:05:11.65" resultid="2558" heatid="7566" lane="0" entrytime="00:05:09.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:14.17" />
                    <SPLIT distance="150" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:32.59" />
                    <SPLIT distance="250" swimtime="00:03:12.26" />
                    <SPLIT distance="300" swimtime="00:03:52.33" />
                    <SPLIT distance="350" swimtime="00:04:32.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="2565">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2566" heatid="7280" lane="9" entrytime="00:03:10.00" />
                <RESULT eventid="1156" points="170" swimtime="00:13:19.95" resultid="2567" heatid="7298" lane="1" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                    <SPLIT distance="150" swimtime="00:02:14.41" />
                    <SPLIT distance="200" swimtime="00:03:02.85" />
                    <SPLIT distance="250" swimtime="00:03:51.92" />
                    <SPLIT distance="300" swimtime="00:04:41.36" />
                    <SPLIT distance="350" swimtime="00:05:31.48" />
                    <SPLIT distance="400" swimtime="00:06:21.57" />
                    <SPLIT distance="450" swimtime="00:07:13.05" />
                    <SPLIT distance="500" swimtime="00:08:04.99" />
                    <SPLIT distance="550" swimtime="00:08:56.98" />
                    <SPLIT distance="600" swimtime="00:09:49.66" />
                    <SPLIT distance="650" swimtime="00:10:42.62" />
                    <SPLIT distance="700" swimtime="00:11:34.96" />
                    <SPLIT distance="750" swimtime="00:12:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="200" swimtime="00:03:25.19" resultid="2568" heatid="7336" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:36.39" />
                    <SPLIT distance="150" swimtime="00:02:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="229" swimtime="00:01:22.07" resultid="2569" heatid="7382" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="237" reactiontime="+99" swimtime="00:01:29.75" resultid="2570" heatid="7419" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="2571" heatid="7463" lane="6" entrytime="00:01:22.00" />
                <RESULT eventid="1625" points="184" reactiontime="+96" swimtime="00:01:24.46" resultid="2572" heatid="7516" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="248" reactiontime="+96" swimtime="00:00:40.14" resultid="2573" heatid="7551" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00709" nation="POL" region="09" clubid="5919" name="MKS Barracuda Białystok" shortname="Barracuda Białystok">
          <ATHLETES>
            <ATHLETE birthdate="1953-10-13" firstname="Mirosław" gender="M" lastname="Gawryluk" nation="POL" athleteid="5932">
              <RESULTS>
                <RESULT eventid="1076" points="129" swimtime="00:00:40.06" resultid="5933" heatid="7250" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1288" points="109" swimtime="00:01:33.89" resultid="5934" heatid="7351" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="129" swimtime="00:01:50.04" resultid="5935" heatid="7416" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="127" swimtime="00:00:50.12" resultid="5936" heatid="7548" lane="7" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-10-29" firstname="Jacek" gender="M" lastname="Gregorczuk" nation="POL" athleteid="5926">
              <RESULTS>
                <RESULT eventid="1076" points="287" swimtime="00:00:30.71" resultid="5927" heatid="7246" lane="3" />
                <RESULT eventid="1288" points="203" swimtime="00:01:16.44" resultid="5928" heatid="7350" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="5929" heatid="7435" lane="4" />
                <RESULT eventid="1513" points="138" swimtime="00:03:11.87" resultid="5930" heatid="7475" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:34.30" />
                    <SPLIT distance="150" swimtime="00:02:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="5931" heatid="7512" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-19" firstname="Hubert" gender="M" lastname="Milewski" nation="POL" athleteid="5918">
              <RESULTS>
                <RESULT eventid="1156" points="241" swimtime="00:11:52.22" resultid="5920" heatid="7297" lane="3" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                    <SPLIT distance="200" swimtime="00:02:41.54" />
                    <SPLIT distance="250" swimtime="00:03:26.20" />
                    <SPLIT distance="300" swimtime="00:04:12.08" />
                    <SPLIT distance="350" swimtime="00:04:58.12" />
                    <SPLIT distance="400" swimtime="00:05:44.90" />
                    <SPLIT distance="450" swimtime="00:06:31.58" />
                    <SPLIT distance="500" swimtime="00:07:18.17" />
                    <SPLIT distance="550" swimtime="00:08:04.65" />
                    <SPLIT distance="600" swimtime="00:08:50.77" />
                    <SPLIT distance="650" swimtime="00:09:37.89" />
                    <SPLIT distance="700" swimtime="00:10:24.03" />
                    <SPLIT distance="750" swimtime="00:11:09.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="318" reactiontime="+96" swimtime="00:02:55.90" resultid="5921" heatid="7338" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                    <SPLIT distance="150" swimtime="00:02:10.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="324" reactiontime="+98" swimtime="00:01:20.89" resultid="5922" heatid="7423" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="251" swimtime="00:06:13.28" resultid="5923" heatid="8153" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                    <SPLIT distance="200" swimtime="00:03:05.83" />
                    <SPLIT distance="250" swimtime="00:03:54.00" />
                    <SPLIT distance="300" swimtime="00:04:43.54" />
                    <SPLIT distance="350" swimtime="00:05:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="231" reactiontime="+93" swimtime="00:02:52.04" resultid="5924" heatid="7532" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:21.24" />
                    <SPLIT distance="150" swimtime="00:02:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="331" reactiontime="+90" swimtime="00:00:36.47" resultid="5925" heatid="7557" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00701" nation="POL" region="01" clubid="3377" name="MKS Dziewiątka Dzierżoniów" shortname="Dziewiątka Dzierżoniów">
          <CONTACT city="Dzierżoniów" email="ewajuraszek99@op.pl" name="Wojtal Andrzej" phone="508 509 429" state="DOLNO" street="Sienkiewicza 13" zip="58-200" />
          <ATHLETES>
            <ATHLETE birthdate="1986-11-23" firstname="Monika" gender="F" lastname="Babicka" nation="POL" athleteid="3390">
              <RESULTS>
                <RESULT eventid="1059" points="328" reactiontime="+79" swimtime="00:00:33.24" resultid="3391" heatid="7239" lane="7" entrytime="00:00:35.36" entrycourse="SCM" />
                <RESULT eventid="1304" points="269" reactiontime="+75" swimtime="00:01:27.52" resultid="3392" heatid="7372" lane="2" entrytime="00:01:27.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="310" reactiontime="+73" swimtime="00:00:35.99" resultid="3393" heatid="7429" lane="8" entrytime="00:00:39.36" entrycourse="SCM" />
                <RESULT eventid="1673" points="287" reactiontime="+71" swimtime="00:00:43.29" resultid="3394" heatid="7541" lane="1" entrytime="00:00:45.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-21" firstname="Edyta" gender="F" lastname="Bejster" nation="POL" athleteid="3385">
              <RESULTS>
                <RESULT eventid="1059" points="188" reactiontime="+62" swimtime="00:00:40.02" resultid="3386" heatid="7238" lane="9" entrytime="00:00:39.68" entrycourse="SCM" />
                <RESULT eventid="1304" points="148" reactiontime="+99" swimtime="00:01:46.72" resultid="3387" heatid="7370" lane="7" entrytime="00:01:44.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="76" reactiontime="+95" swimtime="00:00:57.50" resultid="3388" heatid="7427" lane="1" entrytime="00:00:52.85" entrycourse="SCM" />
                <RESULT eventid="1673" points="158" reactiontime="+81" swimtime="00:00:52.80" resultid="3389" heatid="7539" lane="0" entrytime="00:00:53.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-11-06" firstname="Zuzanna" gender="F" lastname="Pisarska" nation="POL" athleteid="3378">
              <RESULTS>
                <RESULT eventid="1059" points="617" reactiontime="+76" swimtime="00:00:26.93" resultid="3379" heatid="7245" lane="5" entrytime="00:00:27.33" entrycourse="SCM" />
                <RESULT eventid="1207" points="552" reactiontime="+59" swimtime="00:00:31.28" resultid="3380" heatid="7314" lane="6" entrytime="00:00:31.67" entrycourse="SCM" />
                <RESULT eventid="1304" points="576" reactiontime="+71" swimtime="00:01:07.89" resultid="3381" heatid="7376" lane="8" entrytime="00:01:10.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="591" reactiontime="+66" swimtime="00:00:29.05" resultid="3382" heatid="7434" lane="5" entrytime="00:00:29.43" entrycourse="SCM" />
                <RESULT eventid="1465" points="506" reactiontime="+60" swimtime="00:01:09.02" resultid="3383" heatid="7457" lane="5" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="547" reactiontime="+66" swimtime="00:01:06.77" resultid="3384" heatid="7511" lane="2" entrytime="00:01:09.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="16" clubid="3738" name="MKS Neptun Stargard" shortname="Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1973-02-20" firstname="Mariusz" gender="M" lastname="Chrzan" nation="POL" athleteid="3739">
              <RESULTS>
                <RESULT eventid="1076" points="446" swimtime="00:00:26.51" resultid="3740" heatid="7267" lane="0" entrytime="00:00:26.10" />
                <RESULT eventid="1108" points="434" reactiontime="+71" swimtime="00:02:24.77" resultid="3741" heatid="7285" lane="8" entrytime="00:02:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="390" reactiontime="+76" swimtime="00:00:30.40" resultid="3742" heatid="7325" lane="5" entrytime="00:00:30.10" />
                <RESULT eventid="1320" points="442" reactiontime="+71" swimtime="00:01:05.98" resultid="3743" heatid="7389" lane="0" entrytime="00:01:04.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="417" reactiontime="+79" swimtime="00:00:29.11" resultid="3744" heatid="7449" lane="0" entrytime="00:00:27.70" />
                <RESULT eventid="1481" points="434" reactiontime="+78" swimtime="00:01:04.52" resultid="3745" heatid="7467" lane="8" entrytime="00:01:04.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="438" reactiontime="+63" swimtime="00:02:19.07" resultid="3746" heatid="7536" lane="2" entrytime="00:02:21.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01201" nation="POL" region="01" clubid="1995" name="MKS Piast Głogów" shortname="Piast Głogów">
          <CONTACT email="skib0303@wp.pl" name="Skiba" phone="667122270" />
          <ATHLETES>
            <ATHLETE birthdate="1977-01-12" firstname="Przemysław" gender="M" lastname="Sosiński" nation="POL" athleteid="1996">
              <RESULTS>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="1997" heatid="7423" lane="9" entrytime="00:01:19.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="1998" heatid="7558" lane="7" entrytime="00:00:34.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04501" nation="POL" region="DOL" clubid="2595" name="MKS Swim Academy Termy Jakuba Oława" shortname="Swim Academy Termy Jakuba Oław">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOL" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-27" firstname="Magdalena" gender="F" lastname="Mruk" nation="POL" license="104501600044" athleteid="2596">
              <RESULTS>
                <RESULT eventid="1304" points="411" reactiontime="+88" swimtime="00:01:15.99" resultid="2597" heatid="7373" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="427" reactiontime="+90" swimtime="00:01:22.76" resultid="2598" heatid="7412" lane="6" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="417" reactiontime="+85" swimtime="00:00:32.61" resultid="2599" heatid="7432" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="1673" points="455" reactiontime="+88" swimtime="00:00:37.12" resultid="2600" heatid="7543" lane="6" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" nation="POL" region="12" clubid="2197" name="MOSiR Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Żak Marek" phone="780063689" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-01" firstname="Zbigniew" gender="M" lastname="Broda" nation="POL" athleteid="5765" />
            <ATHLETE birthdate="1967-11-05" firstname="Krzysztof" gender="M" lastname="Dudek" nation="POL" athleteid="5762" />
            <ATHLETE birthdate="1960-07-13" firstname="Włodzimierz" gender="M" lastname="Mitoraj" nation="POL" athleteid="4358">
              <RESULTS>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="4359" heatid="7417" lane="8" entrytime="00:01:40.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4360" heatid="7550" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="501012700001" athleteid="2198">
              <RESULTS>
                <RESULT eventid="1076" points="207" reactiontime="+98" swimtime="00:00:34.23" resultid="2199" heatid="7253" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1108" points="123" reactiontime="+94" swimtime="00:03:40.37" resultid="2200" heatid="7278" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="107" reactiontime="+94" swimtime="00:04:12.97" resultid="2201" heatid="7333" lane="3" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.97" />
                    <SPLIT distance="100" swimtime="00:02:00.85" />
                    <SPLIT distance="150" swimtime="00:03:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="152" reactiontime="+95" swimtime="00:01:34.05" resultid="2202" heatid="7379" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="185" reactiontime="+91" swimtime="00:00:38.11" resultid="2203" heatid="7439" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1577" points="107" reactiontime="+98" swimtime="00:08:15.18" resultid="2204" heatid="8154" lane="7" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.34" />
                    <SPLIT distance="100" swimtime="00:02:03.04" />
                    <SPLIT distance="150" swimtime="00:03:09.80" />
                    <SPLIT distance="200" swimtime="00:04:16.27" />
                    <SPLIT distance="250" swimtime="00:05:21.77" />
                    <SPLIT distance="300" swimtime="00:06:27.54" />
                    <SPLIT distance="350" swimtime="00:07:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="107" swimtime="00:01:41.08" resultid="2205" heatid="7514" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="173" reactiontime="+89" swimtime="00:00:45.28" resultid="2206" heatid="7550" lane="9" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-05-04" firstname="Stanisław" gender="M" lastname="Sejmicki" nation="POL" athleteid="5766" />
            <ATHLETE birthdate="1959-11-22" firstname="Marek" gender="M" lastname="Żak" nation="POL" athleteid="4355">
              <RESULTS>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="4356" heatid="7319" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="4357" heatid="7462" lane="0" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="172" reactiontime="+85" swimtime="00:02:42.48" resultid="5760" heatid="7404" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:02:13.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4355" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4358" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2198" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5762" number="4" reactiontime="+84" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="207" reactiontime="+56" swimtime="00:02:18.17" resultid="5763" heatid="7493" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:10.50" />
                    <SPLIT distance="150" swimtime="00:01:48.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5765" number="1" reactiontime="+56" />
                    <RELAYPOSITION athleteid="5766" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="2198" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5762" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00908" nation="POL" region="08" clubid="2357" name="Motyl MOSiR Stalowa Wola" shortname="Motyl MOSiR St. Wola">
          <CONTACT city="Stalowa Wola" email="petecka.m@gmail.com" name="Petecka" phone="602829589" street="Al.Jana Pawła II 13/59" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="2358">
              <RESULTS>
                <RESULT eventid="1076" points="473" reactiontime="+76" swimtime="00:00:25.99" resultid="2359" heatid="7253" lane="8" entrytime="00:00:34.99" />
                <RESULT eventid="1108" points="498" reactiontime="+76" swimtime="00:02:18.22" resultid="2360" heatid="7285" lane="2" entrytime="00:02:18.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="517" reactiontime="+72" swimtime="00:00:55.99" resultid="2361" heatid="7365" lane="4" entrytime="00:00:56.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="515" reactiontime="+72" swimtime="00:01:02.70" resultid="2362" heatid="7389" lane="4" entrytime="00:01:02.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="497" reactiontime="+66" swimtime="00:00:27.45" resultid="2363" heatid="7449" lane="6" entrytime="00:00:27.49" />
                <RESULT eventid="1513" points="529" reactiontime="+72" swimtime="00:02:02.86" resultid="2364" heatid="7488" lane="9" entrytime="00:02:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                    <SPLIT distance="150" swimtime="00:01:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="499" reactiontime="+69" swimtime="00:01:00.59" resultid="2365" heatid="7521" lane="3" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="391" reactiontime="+79" swimtime="00:02:24.42" resultid="2366" heatid="7536" lane="9" entrytime="00:02:24.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:47.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="2367">
              <RESULTS>
                <RESULT eventid="1059" points="262" reactiontime="+92" swimtime="00:00:35.81" resultid="2368" heatid="7238" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1092" points="249" reactiontime="+93" swimtime="00:03:13.61" resultid="2369" heatid="7273" lane="8" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:01:33.97" />
                    <SPLIT distance="150" swimtime="00:02:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="247" reactiontime="+87" swimtime="00:03:34.38" resultid="2370" heatid="7330" lane="8" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                    <SPLIT distance="100" swimtime="00:01:42.92" />
                    <SPLIT distance="150" swimtime="00:02:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="251" reactiontime="+88" swimtime="00:01:29.48" resultid="2371" heatid="7372" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="248" reactiontime="+96" swimtime="00:01:39.17" resultid="2372" heatid="7410" lane="0" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="243" reactiontime="+81" swimtime="00:00:39.04" resultid="2373" heatid="7428" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1608" points="188" reactiontime="+95" swimtime="00:01:35.16" resultid="2374" heatid="7508" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="228" reactiontime="+90" swimtime="00:00:46.72" resultid="2375" heatid="7540" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="02" clubid="3875" name="Multisport Team Toruń">
          <CONTACT city="Toruń" email="g.arentewicz@onet.pl" name="Arentewicz" phone="535-763-476" state="KUJ-P" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="3931">
              <RESULTS>
                <RESULT eventid="1108" points="53" reactiontime="+99" swimtime="00:04:50.12" resultid="3932" heatid="7277" lane="1" entrytime="00:05:09.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.57" />
                    <SPLIT distance="100" swimtime="00:02:29.13" />
                    <SPLIT distance="150" swimtime="00:03:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="27" reactiontime="+98" swimtime="00:01:13.97" resultid="3933" heatid="7316" lane="6" entrytime="00:01:15.78" />
                <RESULT eventid="1352" points="28" swimtime="00:05:54.91" resultid="3934" heatid="7394" lane="7" entrytime="00:05:58.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.21" />
                    <SPLIT distance="100" swimtime="00:02:55.46" />
                    <SPLIT distance="150" swimtime="00:04:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="51" swimtime="00:04:26.43" resultid="3935" heatid="7476" lane="0" entrytime="00:03:59.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.87" />
                    <SPLIT distance="100" swimtime="00:02:13.82" />
                    <SPLIT distance="150" swimtime="00:03:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="45" swimtime="00:10:58.34" resultid="3936" heatid="8153" lane="4" entrytime="00:10:31.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.71" />
                    <SPLIT distance="150" swimtime="00:04:20.13" />
                    <SPLIT distance="200" swimtime="00:05:49.78" />
                    <SPLIT distance="250" swimtime="00:07:20.99" />
                    <SPLIT distance="300" swimtime="00:08:49.65" />
                    <SPLIT distance="350" swimtime="00:09:51.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="34" swimtime="00:02:27.98" resultid="3937" heatid="7512" lane="5" entrytime="00:02:50.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="3938" heatid="7583" lane="9" entrytime="00:08:58.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="3885">
              <RESULTS>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="7324" lane="1" entrytime="00:00:32.41" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3887" heatid="7386" lane="9" entrytime="00:01:11.40" />
                <RESULT eventid="1481" points="325" reactiontime="+84" swimtime="00:01:11.09" resultid="3888" heatid="7465" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="311" reactiontime="+82" swimtime="00:05:47.34" resultid="3889" heatid="8157" lane="5" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                    <SPLIT distance="200" swimtime="00:02:42.84" />
                    <SPLIT distance="250" swimtime="00:03:33.59" />
                    <SPLIT distance="300" swimtime="00:04:24.16" />
                    <SPLIT distance="350" swimtime="00:05:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="321" reactiontime="+81" swimtime="00:02:34.17" resultid="3890" heatid="7535" lane="7" entrytime="00:02:29.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="150" swimtime="00:01:54.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="3891" heatid="7577" lane="6" entrytime="00:05:14.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-11" firstname="Kamil" gender="M" lastname="Kordowski" nation="POL" athleteid="3892">
              <RESULTS>
                <RESULT eventid="1076" points="433" reactiontime="+86" swimtime="00:00:26.77" resultid="3893" heatid="7266" lane="7" entrytime="00:00:26.45" />
                <RESULT eventid="1288" points="394" reactiontime="+79" swimtime="00:01:01.30" resultid="3894" heatid="7362" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="343" reactiontime="+73" swimtime="00:00:31.07" resultid="3895" heatid="7444" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1625" points="284" reactiontime="+82" swimtime="00:01:13.12" resultid="3896" heatid="7517" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="3939">
              <RESULTS>
                <RESULT eventid="1076" points="94" swimtime="00:00:44.46" resultid="3940" heatid="7249" lane="9" entrytime="00:00:43.20" />
                <RESULT eventid="1224" points="41" reactiontime="+91" swimtime="00:01:04.09" resultid="3941" heatid="7316" lane="5" entrytime="00:01:08.15" />
                <RESULT eventid="1288" points="79" swimtime="00:01:44.64" resultid="3942" heatid="7350" lane="5" entrytime="00:01:48.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="36" reactiontime="+79" swimtime="00:02:26.83" resultid="3943" heatid="7460" lane="8" entrytime="00:02:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="34" reactiontime="+77" swimtime="00:05:24.99" resultid="3944" heatid="7529" lane="4" entrytime="00:05:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.91" />
                    <SPLIT distance="100" swimtime="00:02:37.92" />
                    <SPLIT distance="150" swimtime="00:04:05.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="3923">
              <RESULTS>
                <RESULT eventid="1076" points="240" reactiontime="+94" swimtime="00:00:32.56" resultid="3924" heatid="7254" lane="2" entrytime="00:00:33.10" />
                <RESULT eventid="1156" points="178" reactiontime="+79" swimtime="00:13:06.92" resultid="3925" heatid="7298" lane="6" entrytime="00:13:08.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:18.23" />
                    <SPLIT distance="200" swimtime="00:03:06.55" />
                    <SPLIT distance="250" swimtime="00:03:56.92" />
                    <SPLIT distance="300" swimtime="00:04:47.66" />
                    <SPLIT distance="350" swimtime="00:05:39.38" />
                    <SPLIT distance="400" swimtime="00:06:30.49" />
                    <SPLIT distance="450" swimtime="00:07:21.55" />
                    <SPLIT distance="500" swimtime="00:08:11.57" />
                    <SPLIT distance="550" swimtime="00:09:02.25" />
                    <SPLIT distance="600" swimtime="00:09:52.63" />
                    <SPLIT distance="650" swimtime="00:10:42.79" />
                    <SPLIT distance="700" swimtime="00:11:32.34" />
                    <SPLIT distance="750" swimtime="00:12:21.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="222" reactiontime="+86" swimtime="00:01:14.15" resultid="3926" heatid="7355" lane="9" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="200" reactiontime="+80" swimtime="00:00:37.14" resultid="3927" heatid="7439" lane="2" entrytime="00:00:37.20" />
                <RESULT eventid="1513" points="181" reactiontime="+80" swimtime="00:02:55.59" resultid="3928" heatid="7478" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                    <SPLIT distance="150" swimtime="00:02:14.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="140" reactiontime="+81" swimtime="00:01:32.41" resultid="3929" heatid="7515" lane="8" entrytime="00:01:33.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="172" reactiontime="+82" swimtime="00:06:21.58" resultid="3930" heatid="7581" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:19.86" />
                    <SPLIT distance="200" swimtime="00:03:08.68" />
                    <SPLIT distance="250" swimtime="00:03:56.65" />
                    <SPLIT distance="300" swimtime="00:04:45.88" />
                    <SPLIT distance="350" swimtime="00:05:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="3906">
              <RESULTS>
                <RESULT eventid="1059" points="96" swimtime="00:00:49.93" resultid="3907" heatid="7235" lane="3" entrytime="00:00:52.08" />
                <RESULT eventid="1172" points="90" reactiontime="+99" swimtime="00:34:10.82" resultid="3908" heatid="7301" lane="1" entrytime="00:35:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.25" />
                    <SPLIT distance="100" swimtime="00:02:01.95" />
                    <SPLIT distance="150" swimtime="00:03:08.47" />
                    <SPLIT distance="200" swimtime="00:04:16.58" />
                    <SPLIT distance="400" swimtime="00:08:52.60" />
                    <SPLIT distance="500" swimtime="00:11:10.53" />
                    <SPLIT distance="750" swimtime="00:16:56.03" />
                    <SPLIT distance="800" swimtime="00:19:14.45" />
                    <SPLIT distance="900" swimtime="00:20:23.12" />
                    <SPLIT distance="950" swimtime="00:21:32.09" />
                    <SPLIT distance="1000" swimtime="00:22:40.92" />
                    <SPLIT distance="1100" swimtime="00:24:59.94" />
                    <SPLIT distance="1150" swimtime="00:26:08.77" />
                    <SPLIT distance="1200" swimtime="00:27:18.06" />
                    <SPLIT distance="1250" swimtime="00:28:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="77" reactiontime="+88" swimtime="00:01:00.09" resultid="3909" heatid="7307" lane="5" entrytime="00:01:01.00" />
                <RESULT eventid="1272" points="85" reactiontime="+94" swimtime="00:01:54.10" resultid="3910" heatid="7341" lane="0" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="81" reactiontime="+91" swimtime="00:02:06.82" resultid="3911" heatid="7453" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="91" swimtime="00:04:05.25" resultid="3912" heatid="7468" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.74" />
                    <SPLIT distance="100" swimtime="00:01:58.16" />
                    <SPLIT distance="150" swimtime="00:03:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="85" reactiontime="+85" swimtime="00:04:30.47" resultid="3913" heatid="7524" lane="4" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="82" swimtime="00:08:57.37" resultid="3914" heatid="7571" lane="0" entrytime="00:08:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                    <SPLIT distance="100" swimtime="00:02:02.11" />
                    <SPLIT distance="150" swimtime="00:03:08.78" />
                    <SPLIT distance="200" swimtime="00:04:16.89" />
                    <SPLIT distance="250" swimtime="00:05:27.14" />
                    <SPLIT distance="300" swimtime="00:06:37.25" />
                    <SPLIT distance="350" swimtime="00:07:49.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="3876">
              <RESULTS>
                <RESULT eventid="1059" points="424" reactiontime="+82" swimtime="00:00:30.51" resultid="3877" heatid="7243" lane="5" entrytime="00:00:30.90" />
                <RESULT eventid="1092" points="430" reactiontime="+79" swimtime="00:02:41.39" resultid="3878" heatid="7275" lane="2" entrytime="00:02:37.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:02.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="415" reactiontime="+75" swimtime="00:03:00.29" resultid="3879" heatid="7331" lane="5" entrytime="00:02:59.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                    <SPLIT distance="100" swimtime="00:01:26.20" />
                    <SPLIT distance="150" swimtime="00:02:12.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="423" reactiontime="+77" swimtime="00:01:15.26" resultid="3880" heatid="7375" lane="3" entrytime="00:01:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="407" reactiontime="+76" swimtime="00:01:24.12" resultid="3881" heatid="7413" lane="1" entrytime="00:01:21.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" status="DNS" swimtime="00:00:00.00" resultid="3882" heatid="8151" lane="6" entrytime="00:05:40.51" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="3883" heatid="7544" lane="0" entrytime="00:00:38.47" />
                <RESULT eventid="1721" status="WDR" swimtime="00:00:00.00" resultid="3884" heatid="7567" lane="4" entrytime="00:05:12.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="3945">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3946" heatid="7248" lane="6" entrytime="00:00:46.34" />
                <RESULT eventid="1224" points="69" reactiontime="+83" swimtime="00:00:54.14" resultid="3947" heatid="7317" lane="4" entrytime="00:00:52.05" />
                <RESULT eventid="1256" points="69" reactiontime="+98" swimtime="00:04:51.68" resultid="3948" heatid="7333" lane="2" entrytime="00:04:21.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.87" />
                    <SPLIT distance="100" swimtime="00:02:10.99" />
                    <SPLIT distance="150" swimtime="00:03:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="85" swimtime="00:02:06.24" resultid="3949" heatid="7416" lane="9" entrytime="00:02:05.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="3950" heatid="7460" lane="7" entrytime="00:02:11.56" />
                <RESULT eventid="1689" points="83" reactiontime="+89" swimtime="00:00:57.67" resultid="3951" heatid="7548" lane="8" entrytime="00:00:52.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-24" firstname="Anita" gender="F" lastname="Śliwa" nation="POL" athleteid="3915">
              <RESULTS>
                <RESULT eventid="1059" points="236" swimtime="00:00:37.07" resultid="3916" heatid="7238" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1172" points="215" swimtime="00:25:34.46" resultid="3917" heatid="7300" lane="9" entrytime="00:27:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:30.44" />
                    <SPLIT distance="150" swimtime="00:02:20.58" />
                    <SPLIT distance="200" swimtime="00:03:12.11" />
                    <SPLIT distance="250" swimtime="00:04:03.76" />
                    <SPLIT distance="300" swimtime="00:04:55.71" />
                    <SPLIT distance="350" swimtime="00:05:47.77" />
                    <SPLIT distance="400" swimtime="00:06:39.82" />
                    <SPLIT distance="450" swimtime="00:07:31.55" />
                    <SPLIT distance="500" swimtime="00:08:23.09" />
                    <SPLIT distance="550" swimtime="00:09:14.79" />
                    <SPLIT distance="600" swimtime="00:10:06.54" />
                    <SPLIT distance="650" swimtime="00:10:59.38" />
                    <SPLIT distance="700" swimtime="00:11:51.35" />
                    <SPLIT distance="750" swimtime="00:12:43.08" />
                    <SPLIT distance="800" swimtime="00:13:34.94" />
                    <SPLIT distance="850" swimtime="00:14:26.62" />
                    <SPLIT distance="900" swimtime="00:15:18.09" />
                    <SPLIT distance="950" swimtime="00:16:09.51" />
                    <SPLIT distance="1000" swimtime="00:17:02.16" />
                    <SPLIT distance="1050" swimtime="00:17:53.72" />
                    <SPLIT distance="1100" swimtime="00:18:45.12" />
                    <SPLIT distance="1150" swimtime="00:19:37.07" />
                    <SPLIT distance="1200" swimtime="00:20:28.62" />
                    <SPLIT distance="1250" swimtime="00:21:20.62" />
                    <SPLIT distance="1300" swimtime="00:22:12.12" />
                    <SPLIT distance="1350" swimtime="00:23:03.96" />
                    <SPLIT distance="1400" swimtime="00:23:55.27" />
                    <SPLIT distance="1450" swimtime="00:24:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="221" swimtime="00:01:23.08" resultid="3918" heatid="7342" lane="5" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="182" reactiontime="+90" swimtime="00:01:36.93" resultid="3919" heatid="7454" lane="6" entrytime="00:01:37.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="213" swimtime="00:03:04.80" resultid="3920" heatid="7470" lane="1" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="198" swimtime="00:03:24.37" resultid="3921" heatid="7525" lane="5" entrytime="00:03:32.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="150" swimtime="00:02:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="199" swimtime="00:06:40.52" resultid="3922" heatid="7570" lane="3" entrytime="00:06:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:32.23" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                    <SPLIT distance="200" swimtime="00:03:16.50" />
                    <SPLIT distance="250" swimtime="00:04:08.94" />
                    <SPLIT distance="300" swimtime="00:05:00.83" />
                    <SPLIT distance="350" swimtime="00:05:52.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Toruń Multisport Team1" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="86" reactiontime="+89" swimtime="00:03:24.11" resultid="3952" heatid="7403" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.99" />
                    <SPLIT distance="100" swimtime="00:01:57.40" />
                    <SPLIT distance="150" swimtime="00:02:36.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3939" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3945" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3923" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3931" number="4" reactiontime="+94" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Toruń Multisport Team2" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="98" swimtime="00:02:57.30" resultid="3953" heatid="7493" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:36.20" />
                    <SPLIT distance="150" swimtime="00:02:23.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3939" number="1" />
                    <RELAYPOSITION athleteid="3945" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3931" number="3" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3923" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NADECA" nation="POL" region="14" clubid="3462" name="Nabaiji Team Decathlon">
          <CONTACT city="Gdańsk" email="martyna.gorajewska@decathlon.com" name="Górajewska Martyna" phone="601990157" street="Szczęśliwa 1" zip="80-176" />
          <ATHLETES>
            <ATHLETE birthdate="1986-11-21" firstname="Laura" gender="F" lastname="Abucewicz" nation="POL" athleteid="3514">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3515" heatid="7236" lane="1" entrytime="00:00:47.59" />
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="3516" heatid="7308" lane="5" entrytime="00:00:54.02" />
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="3518" heatid="7524" lane="8" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="3519" heatid="7538" lane="2" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-06" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="3506">
              <RESULTS>
                <RESULT eventid="1076" points="538" reactiontime="+74" swimtime="00:00:24.90" resultid="3507" heatid="7269" lane="4" entrytime="00:00:24.50" />
                <RESULT eventid="1156" points="350" reactiontime="+99" swimtime="00:10:28.79" resultid="3508" heatid="7294" lane="7" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                    <SPLIT distance="200" swimtime="00:02:20.72" />
                    <SPLIT distance="250" swimtime="00:02:58.36" />
                    <SPLIT distance="300" swimtime="00:03:37.07" />
                    <SPLIT distance="350" swimtime="00:04:17.02" />
                    <SPLIT distance="400" swimtime="00:04:57.72" />
                    <SPLIT distance="450" swimtime="00:05:38.61" />
                    <SPLIT distance="500" swimtime="00:06:19.97" />
                    <SPLIT distance="550" swimtime="00:07:01.03" />
                    <SPLIT distance="600" swimtime="00:07:42.74" />
                    <SPLIT distance="650" swimtime="00:08:24.62" />
                    <SPLIT distance="700" swimtime="00:09:06.75" />
                    <SPLIT distance="750" swimtime="00:09:48.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="545" reactiontime="+75" swimtime="00:00:54.99" resultid="3509" heatid="7366" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="392" reactiontime="+82" swimtime="00:02:27.85" resultid="3510" heatid="7398" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                    <SPLIT distance="150" swimtime="00:01:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="419" reactiontime="+81" swimtime="00:05:14.49" resultid="3511" heatid="8158" lane="3" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                    <SPLIT distance="200" swimtime="00:02:27.37" />
                    <SPLIT distance="250" swimtime="00:03:11.93" />
                    <SPLIT distance="300" swimtime="00:03:57.44" />
                    <SPLIT distance="350" swimtime="00:04:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="465" reactiontime="+77" swimtime="00:01:02.02" resultid="3512" heatid="7521" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="414" reactiontime="+76" swimtime="00:04:44.61" resultid="3513" heatid="7575" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:40.90" />
                    <SPLIT distance="200" swimtime="00:02:17.01" />
                    <SPLIT distance="250" swimtime="00:02:53.39" />
                    <SPLIT distance="300" swimtime="00:03:30.95" />
                    <SPLIT distance="350" swimtime="00:04:07.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-07" firstname="Jan" gender="M" lastname="Dalke" nation="POL" athleteid="3534">
              <RESULTS>
                <RESULT eventid="1076" points="318" reactiontime="+97" swimtime="00:00:29.67" resultid="3535" heatid="7246" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-27" firstname="Michał" gender="M" lastname="Diakonow" nation="POL" athleteid="3588">
              <RESULTS>
                <RESULT eventid="1076" points="466" swimtime="00:00:26.12" resultid="3589" heatid="7265" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="1449" points="327" reactiontime="+86" swimtime="00:00:31.55" resultid="3590" heatid="7447" lane="7" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-31" firstname="Agnieszka" gender="F" lastname="Dusza-Sabadasz" nation="POL" athleteid="3524">
              <RESULTS>
                <RESULT eventid="1059" points="229" reactiontime="+85" swimtime="00:00:37.45" resultid="3525" heatid="7238" lane="3" entrytime="00:00:37.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-06" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="3463">
              <RESULTS>
                <RESULT eventid="1059" points="385" reactiontime="+81" swimtime="00:00:31.50" resultid="3464" heatid="7243" lane="4" entrytime="00:00:30.80" />
                <RESULT eventid="1304" points="348" reactiontime="+79" swimtime="00:01:20.28" resultid="3465" heatid="7373" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="366" reactiontime="+83" swimtime="00:01:27.16" resultid="3466" heatid="7412" lane="0" entrytime="00:01:30.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="371" reactiontime="+79" swimtime="00:00:39.73" resultid="3467" heatid="7543" lane="3" entrytime="00:00:39.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="3468">
              <RESULTS>
                <RESULT eventid="1059" points="397" reactiontime="+80" swimtime="00:00:31.18" resultid="3469" heatid="7243" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1272" points="383" reactiontime="+87" swimtime="00:01:09.17" resultid="3470" heatid="7345" lane="4" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="414" reactiontime="+78" swimtime="00:02:28.09" resultid="3471" heatid="7473" lane="9" entrytime="00:02:31.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:50.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-27" firstname="Aneta" gender="F" lastname="Konkel" nation="POL" athleteid="3569">
              <RESULTS>
                <RESULT eventid="1240" points="116" swimtime="00:04:35.22" resultid="3570" heatid="7327" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.83" />
                    <SPLIT distance="100" swimtime="00:02:06.44" />
                    <SPLIT distance="150" swimtime="00:03:22.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="129" swimtime="00:02:03.39" resultid="3571" heatid="7407" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="3572" heatid="7452" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-10-02" firstname="Agnieszka" gender="F" lastname="Kos" nation="POL" athleteid="3552">
              <RESULTS>
                <RESULT eventid="1272" points="193" reactiontime="+89" swimtime="00:01:26.83" resultid="3553" heatid="7342" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="3554" heatid="7469" lane="8" entrytime="00:03:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-17" firstname="Tomasz" gender="M" lastname="Kosmala" nation="POL" athleteid="3541">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3542" heatid="7249" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3543" heatid="7352" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3544" heatid="7476" lane="4" entrytime="00:03:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-18" firstname="Dawid" gender="M" lastname="Kułakowski" nation="POL" athleteid="3548">
              <RESULTS>
                <RESULT eventid="1288" points="185" reactiontime="+45" swimtime="00:01:18.83" resultid="3549" heatid="7354" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="152" swimtime="00:03:06.13" resultid="3550" heatid="7479" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:16.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="142" swimtime="00:06:46.50" resultid="3551" heatid="7580" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                    <SPLIT distance="200" swimtime="00:03:13.52" />
                    <SPLIT distance="250" swimtime="00:04:07.03" />
                    <SPLIT distance="300" swimtime="00:05:01.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-11-30" firstname="Andrei" gender="M" lastname="Lehatski" nation="POL" athleteid="3476">
              <RESULTS>
                <RESULT eventid="1076" points="468" reactiontime="+81" swimtime="00:00:26.09" resultid="3477" heatid="7265" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="1288" points="433" reactiontime="+80" swimtime="00:00:59.38" resultid="3478" heatid="7362" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="338" reactiontime="+81" swimtime="00:00:31.20" resultid="3479" heatid="7446" lane="4" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="3480">
              <RESULTS>
                <RESULT eventid="1689" points="488" reactiontime="+93" swimtime="00:00:32.05" resultid="3481" heatid="7558" lane="6" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-05-04" firstname="Anna" gender="F" lastname="Majewska" nation="POL" athleteid="3561">
              <RESULTS>
                <RESULT eventid="1304" points="217" reactiontime="+80" swimtime="00:01:33.98" resultid="3562" heatid="7370" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-02" firstname="Karolina" gender="F" lastname="Mazurek-Świstak" nation="POL" athleteid="3520">
              <RESULTS>
                <RESULT eventid="1207" points="513" reactiontime="+76" swimtime="00:00:32.06" resultid="3521" heatid="7314" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1304" points="542" reactiontime="+78" swimtime="00:01:09.30" resultid="3522" heatid="7375" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="495" reactiontime="+74" swimtime="00:00:36.10" resultid="3523" heatid="7544" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1465" points="504" reactiontime="+81" swimtime="00:01:09.12" resultid="8229" heatid="7452" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-30" firstname="Tomasz" gender="M" lastname="Mirek" nation="POL" athleteid="3545">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3546" heatid="7248" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3547" heatid="7351" lane="3" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-17" firstname="Urszula" gender="F" lastname="Moczulska" nation="POL" athleteid="3591">
              <RESULTS>
                <RESULT eventid="1059" points="149" swimtime="00:00:43.20" resultid="3592" heatid="7234" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-06-25" firstname="Rafał" gender="M" lastname="Młynek" nation="POL" athleteid="3563">
              <RESULTS>
                <RESULT eventid="1417" points="254" reactiontime="+79" swimtime="00:01:27.72" resultid="3564" heatid="7415" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-07" firstname="Marzena" gender="F" lastname="Piekarczyk" nation="POL" athleteid="3482">
              <RESULTS>
                <RESULT eventid="1059" points="294" swimtime="00:00:34.45" resultid="3483" heatid="7241" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1272" points="280" swimtime="00:01:16.74" resultid="3484" heatid="7343" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="204" swimtime="00:03:07.57" resultid="3485" heatid="7469" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:02:20.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Kamila" gender="F" lastname="Popielarz" nation="POL" athleteid="3503">
              <RESULTS>
                <RESULT eventid="1207" points="72" reactiontime="+86" swimtime="00:01:01.52" resultid="3504" heatid="7308" lane="6" entrytime="00:00:55.00" />
                <RESULT eventid="1272" points="88" swimtime="00:01:52.63" resultid="3505" heatid="7341" lane="9" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-17" firstname="Paweł" gender="M" lastname="Radziński" nation="POL" athleteid="3580">
              <RESULTS>
                <RESULT eventid="1076" points="393" reactiontime="+93" swimtime="00:00:27.64" resultid="3581" heatid="7265" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3582" heatid="7365" lane="9" entrytime="00:00:58.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3583" heatid="7485" lane="4" entrytime="00:02:11.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-04" firstname="Tomasz" gender="M" lastname="Sabadasz" nation="POL" athleteid="3526">
              <RESULTS>
                <RESULT eventid="1108" points="200" swimtime="00:03:07.41" resultid="3527" heatid="7280" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                    <SPLIT distance="150" swimtime="00:02:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="218" reactiontime="+74" swimtime="00:01:23.50" resultid="3528" heatid="7380" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="203" reactiontime="+75" swimtime="00:06:40.69" resultid="3529" heatid="8156" lane="8" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="100" swimtime="00:01:33.91" />
                    <SPLIT distance="150" swimtime="00:02:28.07" />
                    <SPLIT distance="200" swimtime="00:03:19.72" />
                    <SPLIT distance="250" swimtime="00:04:14.61" />
                    <SPLIT distance="300" swimtime="00:05:09.98" />
                    <SPLIT distance="350" swimtime="00:05:56.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-25" firstname="Kamil" gender="M" lastname="Siwik" nation="POL" athleteid="3530">
              <RESULTS>
                <RESULT eventid="1076" points="183" reactiontime="+98" swimtime="00:00:35.68" resultid="3531" heatid="7247" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-08-10" firstname="Robert" gender="M" lastname="Sowa" nation="POL" athleteid="3494">
              <RESULTS>
                <RESULT eventid="1108" points="420" reactiontime="+97" swimtime="00:02:26.31" resultid="3495" heatid="7284" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="417" swimtime="00:09:53.27" resultid="3496" heatid="7295" lane="4" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.45" />
                    <SPLIT distance="200" swimtime="00:02:24.50" />
                    <SPLIT distance="250" swimtime="00:03:02.61" />
                    <SPLIT distance="300" swimtime="00:03:41.22" />
                    <SPLIT distance="350" swimtime="00:04:20.55" />
                    <SPLIT distance="400" swimtime="00:04:59.57" />
                    <SPLIT distance="450" swimtime="00:05:37.80" />
                    <SPLIT distance="500" swimtime="00:06:15.92" />
                    <SPLIT distance="550" swimtime="00:06:53.42" />
                    <SPLIT distance="600" swimtime="00:07:30.57" />
                    <SPLIT distance="650" swimtime="00:08:07.51" />
                    <SPLIT distance="700" swimtime="00:08:44.15" />
                    <SPLIT distance="750" swimtime="00:09:20.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="396" reactiontime="+73" swimtime="00:00:30.25" resultid="3497" heatid="7325" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3498" heatid="7388" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1481" points="442" reactiontime="+71" swimtime="00:01:04.13" resultid="3499" heatid="7466" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="3500" heatid="8158" lane="2" entrytime="00:05:15.00" />
                <RESULT eventid="1657" points="419" reactiontime="+72" swimtime="00:02:21.06" resultid="3501" heatid="7535" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="433" reactiontime="+92" swimtime="00:04:40.39" resultid="3502" heatid="7575" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:41.06" />
                    <SPLIT distance="200" swimtime="00:02:16.96" />
                    <SPLIT distance="250" swimtime="00:02:53.47" />
                    <SPLIT distance="300" swimtime="00:03:30.60" />
                    <SPLIT distance="350" swimtime="00:04:07.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-18" firstname="Magdalena" gender="F" lastname="Sproska" nation="POL" athleteid="3555">
              <RESULTS>
                <RESULT eventid="1304" points="429" reactiontime="+82" swimtime="00:01:14.92" resultid="3556" heatid="7375" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="436" reactiontime="+78" swimtime="00:00:32.14" resultid="3557" heatid="7432" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-18" firstname="Emil" gender="M" lastname="Strumiński" nation="POL" athleteid="3486">
              <RESULTS>
                <RESULT eventid="1076" points="537" reactiontime="+74" swimtime="00:00:24.92" resultid="3487" heatid="7267" lane="3" entrytime="00:00:25.90" />
                <RESULT eventid="1108" points="384" reactiontime="+75" swimtime="00:02:30.75" resultid="3488" heatid="7284" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="562" reactiontime="+78" swimtime="00:00:54.43" resultid="3489" heatid="7366" lane="0" entrytime="00:00:56.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="381" reactiontime="+80" swimtime="00:02:29.30" resultid="3490" heatid="7398" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="517" reactiontime="+69" swimtime="00:00:27.09" resultid="3491" heatid="7449" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1513" points="505" reactiontime="+76" swimtime="00:02:04.73" resultid="3492" heatid="7486" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:01:00.62" />
                    <SPLIT distance="150" swimtime="00:01:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="490" reactiontime="+76" swimtime="00:01:00.96" resultid="3493" heatid="7521" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-19" firstname="Tomasz" gender="M" lastname="Sypuła" nation="POL" athleteid="3584">
              <RESULTS>
                <RESULT eventid="1076" points="350" reactiontime="+84" swimtime="00:00:28.74" resultid="3585" heatid="7265" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1288" points="286" reactiontime="+84" swimtime="00:01:08.15" resultid="3586" heatid="7364" lane="5" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="250" reactiontime="+86" swimtime="00:00:34.50" resultid="3587" heatid="7447" lane="2" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-09-22" firstname="Marta" gender="F" lastname="Szulżycka" nation="POL" athleteid="3558">
              <RESULTS>
                <RESULT eventid="1272" points="283" reactiontime="+98" swimtime="00:01:16.47" resultid="3559" heatid="7343" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="252" reactiontime="+95" swimtime="00:02:54.83" resultid="3560" heatid="7471" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-07-28" firstname="Julia" gender="F" lastname="Tomczak" nation="POL" athleteid="3536">
              <RESULTS>
                <RESULT eventid="1059" points="359" reactiontime="+98" swimtime="00:00:32.24" resultid="3537" heatid="7243" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1207" points="353" reactiontime="+63" swimtime="00:00:36.32" resultid="3538" heatid="7306" lane="6" />
                <RESULT eventid="1304" points="293" reactiontime="+90" swimtime="00:01:25.04" resultid="3539" heatid="7368" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="278" reactiontime="+71" swimtime="00:01:24.23" resultid="3540" heatid="7452" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-03" firstname="Mateusz" gender="M" lastname="Turowski" nation="POL" athleteid="3575">
              <RESULTS>
                <RESULT eventid="1076" points="301" reactiontime="+91" swimtime="00:00:30.23" resultid="3576" heatid="7259" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-25" firstname="Filip" gender="M" lastname="Wasielewski" nation="POL" athleteid="3472">
              <RESULTS>
                <RESULT eventid="1076" points="389" reactiontime="+71" swimtime="00:00:27.74" resultid="3473" heatid="7264" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1288" points="315" reactiontime="+77" swimtime="00:01:06.00" resultid="3474" heatid="7358" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="381" reactiontime="+71" swimtime="00:00:29.98" resultid="3475" heatid="7447" lane="9" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-25" firstname="Kamil" gender="M" lastname="Ziemianin" nation="POL" athleteid="3565">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3566" heatid="7338" lane="7" entrytime="00:02:49.00" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="3567" heatid="7424" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="3568" heatid="7560" lane="1" entrytime="00:00:32.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-13" firstname="Aleksander" gender="M" lastname="Ziemiński" nation="POL" athleteid="3532">
              <RESULTS>
                <RESULT eventid="1076" points="200" reactiontime="+97" swimtime="00:00:34.60" resultid="3533" heatid="7252" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Piotr" gender="M" lastname="Ławniczak" nation="POL" athleteid="3577">
              <RESULTS>
                <RESULT eventid="1076" points="354" reactiontime="+81" swimtime="00:00:28.63" resultid="3578" heatid="7265" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1449" points="308" reactiontime="+80" swimtime="00:00:32.20" resultid="3579" heatid="7447" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-18" firstname="Krystian" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1076" points="348" reactiontime="+91" swimtime="00:00:28.80" resultid="3574" heatid="7265" lane="2" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" status="DNS" swimtime="00:00:00.00" resultid="3598" heatid="7405" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3577" number="1" />
                    <RELAYPOSITION athleteid="3565" number="2" />
                    <RELAYPOSITION athleteid="3506" number="3" />
                    <RELAYPOSITION athleteid="3472" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" status="DNS" swimtime="00:00:00.00" resultid="3603" heatid="7493" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3506" number="1" />
                    <RELAYPOSITION athleteid="3472" number="2" />
                    <RELAYPOSITION athleteid="3565" number="3" />
                    <RELAYPOSITION athleteid="3486" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1391" points="353" reactiontime="+81" swimtime="00:02:07.86" resultid="3599" heatid="7403" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:39.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3573" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3575" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="3588" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3580" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="370" reactiontime="+78" swimtime="00:01:53.85" resultid="3604" heatid="7493" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                    <SPLIT distance="150" swimtime="00:01:27.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3577" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3575" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3573" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3494" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1545" status="DNS" swimtime="00:00:00.00" resultid="3605" heatid="7493" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3588" number="1" />
                    <RELAYPOSITION athleteid="3541" number="2" />
                    <RELAYPOSITION athleteid="3545" number="3" />
                    <RELAYPOSITION athleteid="3548" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="387" reactiontime="+84" swimtime="00:02:20.41" resultid="3596" heatid="7401" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:46.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3520" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3463" number="2" />
                    <RELAYPOSITION athleteid="3468" number="3" />
                    <RELAYPOSITION athleteid="3482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" points="417" reactiontime="+76" swimtime="00:02:05.63" resultid="3600" heatid="7489" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:03.08" />
                    <SPLIT distance="150" swimtime="00:01:34.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3520" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3482" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3463" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="3468" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1368" status="WDR" swimtime="00:00:00.00" resultid="3597" heatid="7399" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3514" number="1" />
                    <RELAYPOSITION athleteid="3503" number="2" />
                    <RELAYPOSITION athleteid="3552" number="3" />
                    <RELAYPOSITION athleteid="3482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1529" status="WDR" swimtime="00:00:00.00" resultid="3601" heatid="7489" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3591" number="1" />
                    <RELAYPOSITION athleteid="3503" number="2" />
                    <RELAYPOSITION athleteid="3514" number="3" />
                    <RELAYPOSITION athleteid="3524" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="3602" heatid="7489" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3555" number="1" />
                    <RELAYPOSITION athleteid="3552" number="2" />
                    <RELAYPOSITION athleteid="3558" number="3" />
                    <RELAYPOSITION athleteid="3561" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="494" reactiontime="+75" swimtime="00:01:51.13" resultid="3593" heatid="7286" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.80" />
                    <SPLIT distance="100" swimtime="00:00:50.94" />
                    <SPLIT distance="150" swimtime="00:01:22.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3506" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3486" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3463" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3520" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="465" reactiontime="+76" swimtime="00:02:04.37" resultid="3606" heatid="7562" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:40.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3520" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3463" number="2" />
                    <RELAYPOSITION athleteid="3486" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="3506" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="357" reactiontime="+94" swimtime="00:02:03.79" resultid="3594" heatid="7286" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:00:58.59" />
                    <SPLIT distance="150" swimtime="00:01:32.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3575" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="3573" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3482" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3468" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" status="DNS" swimtime="00:00:00.00" resultid="3607" heatid="7562" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3534" number="1" />
                    <RELAYPOSITION athleteid="3503" number="2" />
                    <RELAYPOSITION athleteid="3468" number="3" />
                    <RELAYPOSITION athleteid="3573" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1124" points="243" reactiontime="+90" swimtime="00:02:20.78" resultid="3595" heatid="7286" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                    <SPLIT distance="100" swimtime="00:00:56.10" />
                    <SPLIT distance="150" swimtime="00:01:36.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3588" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="3534" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3524" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3591" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1705" status="WDR" swimtime="00:00:00.00" resultid="3608" heatid="7562" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3536" number="1" />
                    <RELAYPOSITION athleteid="3555" number="2" />
                    <RELAYPOSITION athleteid="3476" number="3" />
                    <RELAYPOSITION athleteid="3575" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NAZIL" nation="SVK" region="SSO" clubid="2410" name="Nareus Žilina">
          <ATHLETES>
            <ATHLETE birthdate="1960-11-14" firstname="Ratislav" gender="M" lastname="Pavlik" nation="SVK" athleteid="2409">
              <RESULTS>
                <RESULT eventid="1076" points="433" reactiontime="+76" swimtime="00:00:26.77" resultid="2411" heatid="7263" lane="3" entrytime="00:00:27.23" />
                <RESULT eventid="1224" points="373" reactiontime="+77" swimtime="00:00:30.85" resultid="2412" heatid="7325" lane="1" entrytime="00:00:31.03" />
                <RESULT eventid="1320" points="425" reactiontime="+76" swimtime="00:01:06.83" resultid="2413" heatid="7387" lane="3" entrytime="00:01:07.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="384" reactiontime="+78" swimtime="00:01:07.20" resultid="2414" heatid="7466" lane="0" entrytime="00:01:07.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="438" reactiontime="+82" swimtime="00:00:33.23" resultid="2415" heatid="7559" lane="1" entrytime="00:00:33.54" />
                <RESULT eventid="1737" points="225" reactiontime="+78" swimtime="00:05:48.70" resultid="2416" heatid="7579" lane="4" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                    <SPLIT distance="200" swimtime="00:02:41.23" />
                    <SPLIT distance="250" swimtime="00:03:28.67" />
                    <SPLIT distance="300" swimtime="00:04:15.86" />
                    <SPLIT distance="350" swimtime="00:05:02.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NMPRA" nation="CZE" clubid="3078" name="Neptun Masters Praha">
          <ATHLETES>
            <ATHLETE birthdate="1968-06-15" firstname="Hana" gender="F" lastname="Bohuslávková" nation="CZE" athleteid="3080">
              <RESULTS>
                <RESULT eventid="1240" points="479" reactiontime="+86" swimtime="00:02:51.95" resultid="3090" heatid="7331" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:23.06" />
                    <SPLIT distance="150" swimtime="00:02:07.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="431" reactiontime="+84" swimtime="00:01:14.77" resultid="3091" heatid="7374" lane="3" entrytime="00:01:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="468" reactiontime="+81" swimtime="00:01:20.29" resultid="3092" heatid="7413" lane="7" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="467" reactiontime="+83" swimtime="00:00:36.79" resultid="3093" heatid="7545" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-06" firstname="Věra" gender="F" lastname="Civínová" nation="CZE" athleteid="3079">
              <RESULTS>
                <RESULT eventid="1272" points="276" reactiontime="+89" swimtime="00:01:17.13" resultid="3086" heatid="7344" lane="9" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="258" reactiontime="+94" swimtime="00:00:38.29" resultid="3087" heatid="7430" lane="8" entrytime="00:00:37.20" />
                <RESULT eventid="1497" points="281" reactiontime="+94" swimtime="00:02:48.47" resultid="3088" heatid="7471" lane="1" entrytime="00:02:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="225" reactiontime="+86" swimtime="00:01:29.67" resultid="3089" heatid="7510" lane="1" entrytime="00:01:24.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-04" firstname="Tomáš" gender="M" lastname="Vonšovský" nation="CZE" athleteid="3077">
              <RESULTS>
                <RESULT eventid="1224" points="328" reactiontime="+65" swimtime="00:00:32.20" resultid="3081" heatid="7323" lane="5" entrytime="00:00:33.20" />
                <RESULT eventid="1320" points="340" reactiontime="+78" swimtime="00:01:11.95" resultid="3082" heatid="7384" lane="5" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="356" reactiontime="+79" swimtime="00:00:30.66" resultid="3083" heatid="7444" lane="2" entrytime="00:00:30.90" />
                <RESULT eventid="1625" points="328" reactiontime="+79" swimtime="00:01:09.70" resultid="3084" heatid="7518" lane="9" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="299" reactiontime="+83" swimtime="00:00:37.76" resultid="3085" heatid="7554" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZJG" nation="POL" region="01" clubid="5861" name="Niezreszony Jelenia Góra">
          <ATHLETES>
            <ATHLETE birthdate="1985-06-16" firstname="Anna" gender="F" lastname="Lara" nation="POL" athleteid="5868">
              <RESULTS>
                <RESULT eventid="1140" points="281" swimtime="00:12:11.03" resultid="5869" heatid="7291" lane="0" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:19.39" />
                    <SPLIT distance="150" swimtime="00:02:02.69" />
                    <SPLIT distance="200" swimtime="00:02:47.75" />
                    <SPLIT distance="250" swimtime="00:03:33.97" />
                    <SPLIT distance="300" swimtime="00:04:20.57" />
                    <SPLIT distance="350" swimtime="00:05:07.10" />
                    <SPLIT distance="400" swimtime="00:05:53.39" />
                    <SPLIT distance="450" swimtime="00:06:39.71" />
                    <SPLIT distance="500" swimtime="00:07:26.76" />
                    <SPLIT distance="550" swimtime="00:08:14.13" />
                    <SPLIT distance="600" swimtime="00:09:01.96" />
                    <SPLIT distance="650" swimtime="00:09:49.61" />
                    <SPLIT distance="700" swimtime="00:10:37.45" />
                    <SPLIT distance="750" swimtime="00:11:24.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="272" reactiontime="+96" swimtime="00:01:17.47" resultid="5870" heatid="7342" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="172" reactiontime="+73" swimtime="00:03:34.82" resultid="5871" heatid="7392" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                    <SPLIT distance="150" swimtime="00:02:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="245" reactiontime="+94" swimtime="00:00:38.96" resultid="5872" heatid="7428" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1497" points="271" reactiontime="+99" swimtime="00:02:50.52" resultid="5873" heatid="7470" lane="7" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                    <SPLIT distance="150" swimtime="00:02:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="175" reactiontime="+71" swimtime="00:01:37.51" resultid="5874" heatid="7508" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="269" reactiontime="+51" swimtime="00:06:01.95" resultid="5875" heatid="7569" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                    <SPLIT distance="150" swimtime="00:02:12.58" />
                    <SPLIT distance="200" swimtime="00:02:58.83" />
                    <SPLIT distance="250" swimtime="00:03:44.76" />
                    <SPLIT distance="300" swimtime="00:04:30.83" />
                    <SPLIT distance="350" swimtime="00:05:16.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-05" firstname="Marek" gender="M" lastname="Lipka" nation="POL" athleteid="5860">
              <RESULTS>
                <RESULT eventid="1188" points="175" swimtime="00:25:15.85" resultid="5862" heatid="7304" lane="2" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:32.71" />
                    <SPLIT distance="150" swimtime="00:02:22.96" />
                    <SPLIT distance="200" swimtime="00:03:13.90" />
                    <SPLIT distance="250" swimtime="00:04:04.67" />
                    <SPLIT distance="300" swimtime="00:04:55.76" />
                    <SPLIT distance="350" swimtime="00:05:47.00" />
                    <SPLIT distance="400" swimtime="00:06:38.30" />
                    <SPLIT distance="450" swimtime="00:07:28.98" />
                    <SPLIT distance="500" swimtime="00:08:19.64" />
                    <SPLIT distance="550" swimtime="00:09:10.12" />
                    <SPLIT distance="600" swimtime="00:10:00.66" />
                    <SPLIT distance="650" swimtime="00:10:50.53" />
                    <SPLIT distance="700" swimtime="00:11:41.08" />
                    <SPLIT distance="750" swimtime="00:12:31.69" />
                    <SPLIT distance="800" swimtime="00:13:22.18" />
                    <SPLIT distance="850" swimtime="00:14:12.67" />
                    <SPLIT distance="900" swimtime="00:15:02.77" />
                    <SPLIT distance="950" swimtime="00:15:53.34" />
                    <SPLIT distance="1000" swimtime="00:16:44.61" />
                    <SPLIT distance="1050" swimtime="00:17:36.25" />
                    <SPLIT distance="1100" swimtime="00:18:28.07" />
                    <SPLIT distance="1150" swimtime="00:19:20.32" />
                    <SPLIT distance="1200" swimtime="00:20:11.01" />
                    <SPLIT distance="1250" swimtime="00:21:01.95" />
                    <SPLIT distance="1300" swimtime="00:21:54.43" />
                    <SPLIT distance="1350" swimtime="00:22:45.45" />
                    <SPLIT distance="1400" swimtime="00:23:36.75" />
                    <SPLIT distance="1450" swimtime="00:24:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="180" reactiontime="+97" swimtime="00:01:19.57" resultid="5863" heatid="7355" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="113" reactiontime="+56" swimtime="00:03:43.76" resultid="5864" heatid="7396" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.09" />
                    <SPLIT distance="100" swimtime="00:01:51.24" />
                    <SPLIT distance="150" swimtime="00:02:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="179" reactiontime="+94" swimtime="00:02:56.29" resultid="5865" heatid="7477" lane="4" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="150" swimtime="00:02:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="129" swimtime="00:01:35.14" resultid="5866" heatid="7514" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="171" swimtime="00:06:22.28" resultid="5867" heatid="7580" lane="0" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:30.68" />
                    <SPLIT distance="150" swimtime="00:02:19.10" />
                    <SPLIT distance="200" swimtime="00:03:08.94" />
                    <SPLIT distance="250" swimtime="00:03:58.82" />
                    <SPLIT distance="300" swimtime="00:04:47.25" />
                    <SPLIT distance="350" swimtime="00:05:35.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZKAC" nation="POL" region="15" clubid="2539" name="Niezrzeszeni Kaczory">
          <ATHLETES>
            <ATHLETE birthdate="1982-01-28" firstname="Paweł" gender="M" lastname="Lisiecki" nation="POL" athleteid="2538">
              <RESULTS>
                <RESULT eventid="1076" points="261" swimtime="00:00:31.69" resultid="2540" heatid="7256" lane="0" entrytime="00:00:31.57" />
                <RESULT eventid="1156" points="282" swimtime="00:11:15.92" resultid="2541" heatid="7296" lane="4" entrytime="00:11:03.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:56.55" />
                    <SPLIT distance="200" swimtime="00:02:38.18" />
                    <SPLIT distance="250" swimtime="00:03:20.30" />
                    <SPLIT distance="300" swimtime="00:04:02.96" />
                    <SPLIT distance="350" swimtime="00:04:45.85" />
                    <SPLIT distance="400" swimtime="00:05:28.79" />
                    <SPLIT distance="450" swimtime="00:06:11.96" />
                    <SPLIT distance="500" swimtime="00:06:55.28" />
                    <SPLIT distance="550" swimtime="00:07:38.62" />
                    <SPLIT distance="600" swimtime="00:08:21.81" />
                    <SPLIT distance="650" swimtime="00:09:05.52" />
                    <SPLIT distance="700" swimtime="00:09:49.44" />
                    <SPLIT distance="750" swimtime="00:10:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="190" reactiontime="+93" swimtime="00:00:38.62" resultid="2542" heatid="7321" lane="0" entrytime="00:00:37.72" />
                <RESULT eventid="1288" points="261" swimtime="00:01:10.30" resultid="2543" heatid="7356" lane="3" entrytime="00:01:09.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="240" reactiontime="+87" swimtime="00:01:18.58" resultid="2544" heatid="7459" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="270" reactiontime="+98" swimtime="00:02:33.72" resultid="2545" heatid="7481" lane="9" entrytime="00:02:35.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                    <SPLIT distance="150" swimtime="00:01:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="253" reactiontime="+93" swimtime="00:02:46.94" resultid="2546" heatid="7533" lane="6" entrytime="00:02:47.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:03.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="277" reactiontime="+87" swimtime="00:05:25.47" resultid="2547" heatid="7578" lane="6" entrytime="00:05:27.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:01:56.87" />
                    <SPLIT distance="200" swimtime="00:02:38.92" />
                    <SPLIT distance="250" swimtime="00:03:20.95" />
                    <SPLIT distance="300" swimtime="00:04:03.20" />
                    <SPLIT distance="350" swimtime="00:04:44.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZBIA" nation="POL" region="09" clubid="6868" name="Niezrzeszony Białystok">
          <ATHLETES>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="2427">
              <RESULTS>
                <RESULT eventid="1076" points="389" reactiontime="+79" swimtime="00:00:27.75" resultid="2429" heatid="7261" lane="9" entrytime="00:00:28.25" />
                <RESULT eventid="1108" points="345" reactiontime="+87" swimtime="00:02:36.29" resultid="2430" heatid="7282" lane="3" entrytime="00:02:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="383" reactiontime="+80" swimtime="00:01:01.86" resultid="2431" heatid="7360" lane="5" entrytime="00:01:02.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="353" reactiontime="+81" swimtime="00:01:11.11" resultid="2432" heatid="7385" lane="4" entrytime="00:01:11.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="386" reactiontime="+80" swimtime="00:00:29.87" resultid="2433" heatid="7444" lane="7" entrytime="00:00:30.95" />
                <RESULT eventid="1481" points="294" reactiontime="+72" swimtime="00:01:13.46" resultid="2434" heatid="7464" lane="6" entrytime="00:01:16.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="337" reactiontime="+81" swimtime="00:01:09.09" resultid="2435" heatid="7518" lane="4" entrytime="00:01:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="356" reactiontime="+76" swimtime="00:00:35.61" resultid="2436" heatid="7554" lane="4" entrytime="00:00:37.55" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZGDA" nation="POL" region="10" clubid="5747" name="Niezrzeszony Gdańsk">
          <ATHLETES>
            <ATHLETE birthdate="1961-01-18" firstname="Wojciech" gender="M" lastname="Warchoł" nation="POL" athleteid="5746">
              <RESULTS>
                <RESULT eventid="1320" points="320" reactiontime="+93" swimtime="00:01:13.47" resultid="5748" heatid="7383" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="287" reactiontime="+87" swimtime="00:05:56.69" resultid="5749" heatid="8156" lane="4" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="150" swimtime="00:02:06.52" />
                    <SPLIT distance="200" swimtime="00:02:53.17" />
                    <SPLIT distance="250" swimtime="00:03:44.62" />
                    <SPLIT distance="300" swimtime="00:04:36.15" />
                    <SPLIT distance="350" swimtime="00:05:16.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="289" reactiontime="+84" swimtime="00:05:20.78" resultid="5750" heatid="7578" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:55.38" />
                    <SPLIT distance="200" swimtime="00:02:36.23" />
                    <SPLIT distance="250" swimtime="00:03:17.09" />
                    <SPLIT distance="300" swimtime="00:03:58.82" />
                    <SPLIT distance="350" swimtime="00:04:40.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZGDY" nation="POL" region="10" clubid="2727" name="Niezrzeszony Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1992-08-06" firstname="Kamil" gender="M" lastname="Lubiński" nation="POL" athleteid="3451">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3452" heatid="7262" lane="6" entrytime="00:00:27.90" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="3453" heatid="7282" lane="0" entrytime="00:02:40.00" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3454" heatid="7324" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3455" heatid="7338" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3456" heatid="7387" lane="8" entrytime="00:01:10.00" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="3457" heatid="7422" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="3458" heatid="7465" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="3459" heatid="8157" lane="2" entrytime="00:05:45.00" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="3460" heatid="7534" lane="1" entrytime="00:02:40.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="3461" heatid="7558" lane="2" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka " nation="POL" athleteid="2726">
              <RESULTS>
                <RESULT eventid="1108" points="48" swimtime="00:05:01.59" resultid="2728" heatid="7277" lane="7" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.20" />
                    <SPLIT distance="100" swimtime="00:02:28.80" />
                    <SPLIT distance="150" swimtime="00:03:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="62" swimtime="00:05:02.79" resultid="2729" heatid="7332" lane="3" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.34" />
                    <SPLIT distance="100" swimtime="00:02:25.94" />
                    <SPLIT distance="150" swimtime="00:03:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="36" swimtime="00:05:27.03" resultid="2730" heatid="7394" lane="2" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.10" />
                    <SPLIT distance="100" swimtime="00:02:36.44" />
                    <SPLIT distance="150" swimtime="00:04:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="53" swimtime="00:00:57.70" resultid="2731" heatid="7436" lane="4" entrytime="00:00:56.00" />
                <RESULT eventid="1577" points="51" swimtime="00:10:33.56" resultid="2732" heatid="8153" lane="3" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.97" />
                    <SPLIT distance="100" swimtime="00:02:33.58" />
                    <SPLIT distance="150" swimtime="00:04:00.62" />
                    <SPLIT distance="200" swimtime="00:05:23.89" />
                    <SPLIT distance="250" swimtime="00:06:48.17" />
                    <SPLIT distance="300" swimtime="00:08:10.24" />
                    <SPLIT distance="350" swimtime="00:09:23.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="36" swimtime="00:02:24.48" resultid="2733" heatid="7513" lane="9" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="46" swimtime="00:09:48.61" resultid="2734" heatid="7583" lane="2" entrytime="00:10:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.28" />
                    <SPLIT distance="100" swimtime="00:02:19.94" />
                    <SPLIT distance="150" swimtime="00:03:36.18" />
                    <SPLIT distance="200" swimtime="00:04:52.37" />
                    <SPLIT distance="250" swimtime="00:06:09.62" />
                    <SPLIT distance="300" swimtime="00:07:25.81" />
                    <SPLIT distance="350" swimtime="00:08:39.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZGLI" nation="POL" region="11" clubid="5785" name="Niezrzeszony Gliwice">
          <ATHLETES>
            <ATHLETE birthdate="1983-08-29" firstname="Leszek" gender="M" lastname="Zawadzki" nation="POL" athleteid="5784">
              <RESULTS>
                <RESULT eventid="1076" points="316" swimtime="00:00:29.72" resultid="5786" heatid="7252" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1156" points="278" swimtime="00:11:19.04" resultid="5787" heatid="7297" lane="4" entrytime="00:11:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:52.70" />
                    <SPLIT distance="200" swimtime="00:02:34.05" />
                    <SPLIT distance="250" swimtime="00:03:16.62" />
                    <SPLIT distance="300" swimtime="00:04:00.02" />
                    <SPLIT distance="350" swimtime="00:04:43.48" />
                    <SPLIT distance="400" swimtime="00:05:27.25" />
                    <SPLIT distance="450" swimtime="00:06:11.40" />
                    <SPLIT distance="500" swimtime="00:06:55.59" />
                    <SPLIT distance="550" swimtime="00:07:39.89" />
                    <SPLIT distance="600" swimtime="00:08:24.14" />
                    <SPLIT distance="650" swimtime="00:09:08.48" />
                    <SPLIT distance="700" swimtime="00:09:53.22" />
                    <SPLIT distance="750" swimtime="00:10:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="299" swimtime="00:01:07.16" resultid="5788" heatid="7354" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="291" swimtime="00:02:29.89" resultid="5789" heatid="7476" lane="8" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5790" heatid="7583" lane="8" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZKAL" nation="POL" region="15" clubid="6481" name="Niezrzeszony Kalisz">
          <ATHLETES>
            <ATHLETE birthdate="1964-05-29" firstname="Andrzej" gender="M" lastname="Wiśniewski" nation="POL" athleteid="6480">
              <RESULTS>
                <RESULT eventid="1076" points="142" swimtime="00:00:38.79" resultid="6482" heatid="7251" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZKNU" nation="POL" region="11" clubid="2919" name="Niezrzeszony Knurów">
          <ATHLETES>
            <ATHLETE birthdate="1990-03-14" firstname="Sylwia" gender="F" lastname="Kuśpiet" nation="POL" athleteid="2911">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="2912" heatid="7275" lane="3" entrytime="00:02:36.00" />
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="2913" heatid="7314" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="2914" heatid="7376" lane="9" entrytime="00:01:11.00" />
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="2915" heatid="7413" lane="3" entrytime="00:01:17.00" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="2916" heatid="7432" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="2917" heatid="7511" lane="6" entrytime="00:01:08.00" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="2918" heatid="7545" lane="6" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZLEG" nation="POL" region="14" clubid="5768" name="Niezrzeszony Legionowo">
          <ATHLETES>
            <ATHLETE birthdate="1973-01-14" firstname="Andrzej" gender="M" lastname="Fajdasz" nation="POL" athleteid="5767">
              <RESULTS>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="5769" heatid="7320" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5770" heatid="7361" lane="5" entrytime="00:01:01.50" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="5771" heatid="7382" lane="3" entrytime="00:01:19.00" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="5772" heatid="7464" lane="1" entrytime="00:01:18.50" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5773" heatid="7481" lane="6" entrytime="00:02:30.50" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5774" heatid="7533" lane="4" entrytime="00:02:43.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZLES" nation="POL" region="15" clubid="6870" name="Niezrzeszony Leszno">
          <ATHLETES>
            <ATHLETE birthdate="1985-01-11" firstname="Tomasz" gender="M" lastname="Grzelczak" nation="POL" athleteid="2015">
              <RESULTS>
                <RESULT eventid="1256" points="181" swimtime="00:03:32.31" resultid="2017" heatid="7334" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="116" swimtime="00:01:42.94" resultid="2018" heatid="7378" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="206" swimtime="00:01:34.02" resultid="2019" heatid="7418" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="126" swimtime="00:00:43.35" resultid="2020" heatid="7437" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2021" heatid="7552" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2022" heatid="7581" lane="1" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZLVI" nation="UKR" clubid="5877" name="Niezrzeszony Lviv">
          <ATHLETES>
            <ATHLETE birthdate="1968-05-23" firstname="Igor" gender="M" lastname="Karpenko" nation="UKR" athleteid="5876">
              <RESULTS>
                <RESULT eventid="1417" points="281" reactiontime="+83" swimtime="00:01:24.85" resultid="5878" heatid="7421" lane="9" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="298" reactiontime="+90" swimtime="00:00:37.80" resultid="5879" heatid="7556" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZPIO" nation="POL" region="14" clubid="2377" name="Niezrzeszony Pionki">
          <ATHLETES>
            <ATHLETE birthdate="1981-03-09" firstname="Krystian" gender="M" lastname="Bator" nation="POL" athleteid="2376">
              <RESULTS>
                <RESULT eventid="1076" points="438" reactiontime="+67" swimtime="00:00:26.66" resultid="2378" heatid="7263" lane="9" entrytime="00:00:27.53" />
                <RESULT eventid="1288" points="422" reactiontime="+69" swimtime="00:00:59.89" resultid="2379" heatid="7360" lane="7" entrytime="00:01:03.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="370" reactiontime="+70" swimtime="00:00:30.28" resultid="2380" heatid="7444" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1513" points="323" reactiontime="+70" swimtime="00:02:24.81" resultid="2381" heatid="7482" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                    <SPLIT distance="150" swimtime="00:01:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2382" heatid="7555" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZPIO" nation="POL" region="05" clubid="2523" name="Niezrzeszony Piotrków Tryb.">
          <ATHLETES>
            <ATHLETE birthdate="1966-03-05" firstname="Jarosław" gender="M" lastname="Guziński" nation="POL" athleteid="2522">
              <RESULTS>
                <RESULT eventid="1076" points="228" reactiontime="+84" swimtime="00:00:33.16" resultid="2524" heatid="7252" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2525" heatid="7351" lane="1" entrytime="00:01:40.00" />
                <RESULT eventid="1449" points="165" reactiontime="+99" swimtime="00:00:39.65" resultid="2526" heatid="7437" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="2527" heatid="7514" lane="8" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZPIL" nation="POL" region="15" clubid="2634" name="Niezrzeszony Piła">
          <ATHLETES>
            <ATHLETE birthdate="1944-06-14" firstname="Andrzej" gender="M" lastname="Rusinowicz" nation="POL" athleteid="2633">
              <RESULTS>
                <RESULT eventid="1108" points="63" swimtime="00:04:35.51" resultid="2635" heatid="7277" lane="5" entrytime="00:04:32.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                    <SPLIT distance="100" swimtime="00:02:13.64" />
                    <SPLIT distance="150" swimtime="00:03:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="74" swimtime="00:33:31.47" resultid="2636" heatid="7305" lane="4" entrytime="00:35:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                    <SPLIT distance="100" swimtime="00:02:02.22" />
                    <SPLIT distance="150" swimtime="00:03:09.61" />
                    <SPLIT distance="200" swimtime="00:04:17.13" />
                    <SPLIT distance="250" swimtime="00:05:25.22" />
                    <SPLIT distance="300" swimtime="00:06:36.30" />
                    <SPLIT distance="350" swimtime="00:07:44.70" />
                    <SPLIT distance="400" swimtime="00:08:53.37" />
                    <SPLIT distance="450" swimtime="00:10:02.01" />
                    <SPLIT distance="500" swimtime="00:11:10.19" />
                    <SPLIT distance="550" swimtime="00:12:16.17" />
                    <SPLIT distance="600" swimtime="00:13:24.66" />
                    <SPLIT distance="650" swimtime="00:14:31.70" />
                    <SPLIT distance="700" swimtime="00:15:38.30" />
                    <SPLIT distance="750" swimtime="00:16:46.16" />
                    <SPLIT distance="800" swimtime="00:17:53.31" />
                    <SPLIT distance="850" swimtime="00:19:00.59" />
                    <SPLIT distance="900" swimtime="00:20:07.90" />
                    <SPLIT distance="950" swimtime="00:21:15.45" />
                    <SPLIT distance="1000" swimtime="00:22:22.61" />
                    <SPLIT distance="1050" swimtime="00:23:29.47" />
                    <SPLIT distance="1150" swimtime="00:25:43.24" />
                    <SPLIT distance="1200" swimtime="00:26:50.55" />
                    <SPLIT distance="1250" swimtime="00:27:57.97" />
                    <SPLIT distance="1300" swimtime="00:29:05.20" />
                    <SPLIT distance="1350" swimtime="00:30:11.90" />
                    <SPLIT distance="1400" swimtime="00:31:18.64" />
                    <SPLIT distance="1450" swimtime="00:32:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="66" swimtime="00:04:56.13" resultid="2637" heatid="7333" lane="9" entrytime="00:04:49.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.90" />
                    <SPLIT distance="100" swimtime="00:02:18.77" />
                    <SPLIT distance="150" swimtime="00:03:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="64" swimtime="00:02:05.07" resultid="2638" heatid="7377" lane="5" entrytime="00:01:59.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="66" swimtime="00:02:17.46" resultid="2639" heatid="7415" lane="3" entrytime="00:02:12.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="56" swimtime="00:10:14.48" resultid="2640" heatid="8153" lane="5" entrytime="00:10:31.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.00" />
                    <SPLIT distance="100" swimtime="00:02:33.77" />
                    <SPLIT distance="150" swimtime="00:03:53.79" />
                    <SPLIT distance="200" swimtime="00:05:14.77" />
                    <SPLIT distance="250" swimtime="00:06:38.09" />
                    <SPLIT distance="300" swimtime="00:08:00.64" />
                    <SPLIT distance="350" swimtime="00:09:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="36" swimtime="00:02:24.71" resultid="2641" heatid="7512" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="77" swimtime="00:00:59.20" resultid="2642" heatid="7547" lane="4" entrytime="00:00:57.44" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZPOR" nation="POL" region="01" clubid="3647" name="Niezrzeszony Porajów">
          <ATHLETES>
            <ATHLETE birthdate="1950-05-17" firstname="Tadeusz" gender="M" lastname="Okorski" nation="POL" athleteid="3646">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3648" heatid="7247" lane="8" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="3649" heatid="7299" lane="9" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3650" heatid="7315" lane="3" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3651" heatid="7332" lane="2" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="3652" heatid="7414" lane="3" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="3653" heatid="7459" lane="1" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="3654" heatid="7529" lane="7" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="3655" heatid="7546" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZSOS" nation="POL" region="11" clubid="2052" name="Niezrzeszony Sosnowiec">
          <ATHLETES>
            <ATHLETE birthdate="1977-11-05" firstname="Sebastian" gender="M" lastname="Kapka" nation="POL" athleteid="2051">
              <RESULTS>
                <RESULT eventid="1076" points="338" reactiontime="+76" swimtime="00:00:29.06" resultid="2053" heatid="7256" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1108" points="280" reactiontime="+82" swimtime="00:02:47.43" resultid="2054" heatid="7280" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:02:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="296" reactiontime="+82" swimtime="00:00:33.31" resultid="2055" heatid="7323" lane="7" entrytime="00:00:33.92" />
                <RESULT eventid="1320" points="308" reactiontime="+78" swimtime="00:01:14.35" resultid="2056" heatid="7383" lane="6" entrytime="00:01:16.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="315" reactiontime="+80" swimtime="00:00:31.94" resultid="2057" heatid="7443" lane="7" entrytime="00:00:31.52" />
                <RESULT eventid="1481" points="250" reactiontime="+82" swimtime="00:01:17.59" resultid="2058" heatid="7464" lane="0" entrytime="00:01:19.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="234" reactiontime="+76" swimtime="00:02:51.29" resultid="2059" heatid="7533" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:09.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="290" reactiontime="+77" swimtime="00:00:38.13" resultid="2060" heatid="7550" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWRO" nation="POL" region="01" clubid="5944" name="Niezrzeszony Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1995-04-25" firstname="Adriana" gender="F" lastname="Hofman" nation="POL" athleteid="2224">
              <RESULTS>
                <RESULT eventid="1400" points="417" reactiontime="+73" swimtime="00:01:23.41" resultid="2225" heatid="7413" lane="6" entrytime="00:01:18.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="451" reactiontime="+75" swimtime="00:00:37.23" resultid="2226" heatid="7545" lane="7" entrytime="00:00:35.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-07-12" firstname="Sara" gender="F" lastname="Skrzydłoo" nation="POL" athleteid="6334">
              <RESULTS>
                <RESULT eventid="1059" points="597" reactiontime="+76" swimtime="00:00:27.23" resultid="6335" heatid="7245" lane="6" entrytime="00:00:27.48" />
                <RESULT eventid="1272" points="506" reactiontime="+64" swimtime="00:01:03.03" resultid="6336" heatid="7348" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="471" reactiontime="+63" swimtime="00:01:12.62" resultid="6337" heatid="7376" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="600" reactiontime="+59" swimtime="00:00:28.90" resultid="6338" heatid="7434" lane="4" entrytime="00:00:28.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZZG" nation="POL" region="04" clubid="3322" name="Niezrzeszony Zielona Góra">
          <ATHLETES>
            <ATHLETE birthdate="1974-06-11" firstname="Tomasz" gender="M" lastname="Karczewski" nation="POL" athleteid="3321">
              <RESULTS>
                <RESULT eventid="1076" points="361" reactiontime="+89" swimtime="00:00:28.44" resultid="3323" heatid="7258" lane="3" entrytime="00:00:29.88" />
                <RESULT eventid="1156" points="296" reactiontime="+90" swimtime="00:11:04.65" resultid="3324" heatid="7297" lane="5" entrytime="00:11:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                    <SPLIT distance="200" swimtime="00:02:42.63" />
                    <SPLIT distance="250" swimtime="00:03:26.43" />
                    <SPLIT distance="300" swimtime="00:04:09.69" />
                    <SPLIT distance="350" swimtime="00:04:52.60" />
                    <SPLIT distance="400" swimtime="00:05:35.35" />
                    <SPLIT distance="450" swimtime="00:06:17.66" />
                    <SPLIT distance="500" swimtime="00:07:00.28" />
                    <SPLIT distance="550" swimtime="00:07:42.55" />
                    <SPLIT distance="600" swimtime="00:08:25.12" />
                    <SPLIT distance="650" swimtime="00:09:08.08" />
                    <SPLIT distance="700" swimtime="00:09:49.77" />
                    <SPLIT distance="750" swimtime="00:10:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="353" reactiontime="+86" swimtime="00:01:03.57" resultid="3325" heatid="7358" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="338" reactiontime="+86" swimtime="00:00:31.22" resultid="3326" heatid="7442" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZSWI" nation="POL" region="03" clubid="5881" name="Niezrzeszony Świdnik">
          <ATHLETES>
            <ATHLETE birthdate="1974-10-05" firstname="Tomasz" gender="M" lastname="Sitkowski" nation="POL" athleteid="5880">
              <RESULTS>
                <RESULT eventid="1224" points="287" reactiontime="+94" swimtime="00:00:33.67" resultid="5882" heatid="7322" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="347" reactiontime="+80" swimtime="00:01:11.50" resultid="5883" heatid="7384" lane="3" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="321" reactiontime="+83" swimtime="00:00:31.76" resultid="5884" heatid="7442" lane="7" entrytime="00:00:32.80" />
                <RESULT eventid="1481" points="282" reactiontime="+78" swimtime="00:01:14.49" resultid="5885" heatid="7464" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZLOD" nation="POL" region="05" clubid="2028" name="Niezrzezony Łódź">
          <ATHLETES>
            <ATHLETE birthdate="1979-08-13" firstname="Tomasz" gender="M" lastname="Dębecki" nation="POL" athleteid="2027">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2029" heatid="7264" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2030" heatid="7359" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2031" heatid="7447" lane="6" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-07" firstname="Jacek" gender="M" lastname="Kaczmarski" nation="POL" athleteid="2404">
              <RESULTS>
                <RESULT eventid="1076" points="334" reactiontime="+99" swimtime="00:00:29.20" resultid="2405" heatid="7261" lane="2" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-12-22" firstname="Maciej" gender="M" lastname="Kaczmarski" nation="POL" athleteid="2406">
              <RESULTS>
                <RESULT eventid="1320" points="419" reactiontime="+76" swimtime="00:01:07.13" resultid="2407" heatid="7387" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="475" reactiontime="+72" swimtime="00:00:32.34" resultid="2408" heatid="7558" lane="4" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-12-22" firstname="Przemysław" gender="M" lastname="Kaczmarski" nation="POL" athleteid="2401">
              <RESULTS>
                <RESULT eventid="1076" points="539" reactiontime="+79" swimtime="00:00:24.89" resultid="2402" heatid="7267" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1449" points="497" reactiontime="+72" swimtime="00:00:27.44" resultid="2403" heatid="7450" lane="0" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLBYS" nation="POL" region="01" clubid="2736" name="Olimpijczyk Bystre">
          <ATHLETES>
            <ATHLETE birthdate="1975-12-16" firstname="Piotr" gender="M" lastname="Kielesiński" nation="POL" athleteid="2735">
              <RESULTS>
                <RESULT eventid="1076" points="119" reactiontime="+75" swimtime="00:00:41.17" resultid="2737" heatid="7248" lane="4" entrytime="00:00:44.04" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2738" heatid="7315" lane="4" />
                <RESULT eventid="1288" points="87" swimtime="00:01:41.24" resultid="2739" heatid="7351" lane="9" entrytime="00:01:43.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="117" swimtime="00:01:53.50" resultid="2740" heatid="7416" lane="8" entrytime="00:02:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="2741" heatid="7459" lane="2" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2742" heatid="7548" lane="9" entrytime="00:00:56.65" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAUST" nation="CZE" clubid="5279" name="PK Masters Ústí nad Labem" shortname="Masters Ústí nad Labem">
          <CONTACT email="benova.dana@seznam.cz" name="PK Masters Ústí nad Labem" phone="+420728212656" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Beňová" nation="CZE" swrid="4223032" athleteid="5289">
              <RESULTS>
                <RESULT eventid="1092" points="78" swimtime="00:04:44.35" resultid="5290" heatid="7271" lane="0" entrytime="00:04:48.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.69" />
                    <SPLIT distance="100" swimtime="00:02:23.35" />
                    <SPLIT distance="150" swimtime="00:03:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="84" reactiontime="+86" swimtime="00:34:57.84" resultid="5291" heatid="7301" lane="7" entrytime="00:35:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.77" />
                    <SPLIT distance="100" swimtime="00:02:06.50" />
                    <SPLIT distance="150" swimtime="00:03:14.35" />
                    <SPLIT distance="200" swimtime="00:04:21.34" />
                    <SPLIT distance="250" swimtime="00:05:29.77" />
                    <SPLIT distance="300" swimtime="00:06:38.52" />
                    <SPLIT distance="350" swimtime="00:07:47.74" />
                    <SPLIT distance="400" swimtime="00:08:57.33" />
                    <SPLIT distance="450" swimtime="00:10:06.47" />
                    <SPLIT distance="500" swimtime="00:11:15.95" />
                    <SPLIT distance="550" swimtime="00:12:26.60" />
                    <SPLIT distance="600" swimtime="00:13:36.91" />
                    <SPLIT distance="650" swimtime="00:14:47.36" />
                    <SPLIT distance="700" swimtime="00:15:58.02" />
                    <SPLIT distance="750" swimtime="00:17:07.91" />
                    <SPLIT distance="800" swimtime="00:18:17.98" />
                    <SPLIT distance="850" swimtime="00:19:27.82" />
                    <SPLIT distance="900" swimtime="00:20:37.76" />
                    <SPLIT distance="950" swimtime="00:21:48.76" />
                    <SPLIT distance="1000" swimtime="00:23:00.06" />
                    <SPLIT distance="1050" swimtime="00:24:11.09" />
                    <SPLIT distance="1100" swimtime="00:25:23.15" />
                    <SPLIT distance="1150" swimtime="00:26:35.26" />
                    <SPLIT distance="1200" swimtime="00:27:47.34" />
                    <SPLIT distance="1250" swimtime="00:28:59.99" />
                    <SPLIT distance="1300" swimtime="00:30:11.73" />
                    <SPLIT distance="1350" swimtime="00:31:24.24" />
                    <SPLIT distance="1400" swimtime="00:32:37.20" />
                    <SPLIT distance="1450" swimtime="00:33:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="82" reactiontime="+89" swimtime="00:05:09.23" resultid="5292" heatid="7327" lane="5" entrytime="00:04:56.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.40" />
                    <SPLIT distance="100" swimtime="00:02:27.87" />
                    <SPLIT distance="150" swimtime="00:03:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="45" reactiontime="+90" swimtime="00:05:35.47" resultid="5293" heatid="7391" lane="5" entrytime="00:05:37.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.53" />
                    <SPLIT distance="100" swimtime="00:02:49.46" />
                    <SPLIT distance="150" swimtime="00:04:18.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="77" reactiontime="+72" swimtime="00:04:18.91" resultid="5294" heatid="7468" lane="2" entrytime="00:04:19.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.56" />
                    <SPLIT distance="100" swimtime="00:02:07.22" />
                    <SPLIT distance="150" swimtime="00:03:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="75" reactiontime="+94" swimtime="00:10:12.88" resultid="5295" heatid="8149" lane="8" entrytime="00:10:03.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.41" />
                    <SPLIT distance="100" swimtime="00:02:46.88" />
                    <SPLIT distance="150" swimtime="00:04:06.68" />
                    <SPLIT distance="200" swimtime="00:05:22.97" />
                    <SPLIT distance="250" swimtime="00:06:40.72" />
                    <SPLIT distance="300" swimtime="00:07:56.74" />
                    <SPLIT distance="350" swimtime="00:09:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="77" reactiontime="+84" swimtime="00:04:39.82" resultid="5296" heatid="7524" lane="5" entrytime="00:04:38.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.66" />
                    <SPLIT distance="100" swimtime="00:02:22.00" />
                    <SPLIT distance="150" swimtime="00:03:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="86" reactiontime="+89" swimtime="00:08:47.97" resultid="5297" heatid="7571" lane="9" entrytime="00:08:59.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.69" />
                    <SPLIT distance="100" swimtime="00:02:06.22" />
                    <SPLIT distance="150" swimtime="00:03:13.91" />
                    <SPLIT distance="200" swimtime="00:04:21.72" />
                    <SPLIT distance="250" swimtime="00:05:28.36" />
                    <SPLIT distance="300" swimtime="00:06:35.18" />
                    <SPLIT distance="350" swimtime="00:07:42.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-10" firstname="Václav" gender="M" lastname="Valtr" nation="CZE" swrid="4182881" athleteid="5280">
              <RESULTS>
                <RESULT eventid="1108" points="253" reactiontime="+97" swimtime="00:02:53.25" resultid="5281" heatid="7281" lane="9" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:02:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="236" reactiontime="+97" swimtime="00:22:52.06" resultid="5282" heatid="7303" lane="9" entrytime="00:23:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:24.91" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                    <SPLIT distance="200" swimtime="00:02:55.28" />
                    <SPLIT distance="250" swimtime="00:03:41.03" />
                    <SPLIT distance="300" swimtime="00:04:26.68" />
                    <SPLIT distance="350" swimtime="00:05:12.37" />
                    <SPLIT distance="400" swimtime="00:05:58.20" />
                    <SPLIT distance="450" swimtime="00:06:43.82" />
                    <SPLIT distance="500" swimtime="00:07:29.73" />
                    <SPLIT distance="550" swimtime="00:08:15.64" />
                    <SPLIT distance="600" swimtime="00:09:01.04" />
                    <SPLIT distance="650" swimtime="00:09:46.67" />
                    <SPLIT distance="700" swimtime="00:10:32.19" />
                    <SPLIT distance="750" swimtime="00:11:18.02" />
                    <SPLIT distance="800" swimtime="00:12:03.96" />
                    <SPLIT distance="850" swimtime="00:12:49.56" />
                    <SPLIT distance="900" swimtime="00:13:35.90" />
                    <SPLIT distance="950" swimtime="00:14:22.55" />
                    <SPLIT distance="1000" swimtime="00:15:08.37" />
                    <SPLIT distance="1050" swimtime="00:15:54.80" />
                    <SPLIT distance="1100" swimtime="00:16:43.23" />
                    <SPLIT distance="1150" swimtime="00:17:29.64" />
                    <SPLIT distance="1200" swimtime="00:18:16.39" />
                    <SPLIT distance="1250" swimtime="00:19:02.62" />
                    <SPLIT distance="1300" swimtime="00:19:49.17" />
                    <SPLIT distance="1350" swimtime="00:20:35.58" />
                    <SPLIT distance="1400" swimtime="00:21:21.50" />
                    <SPLIT distance="1450" swimtime="00:22:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="233" reactiontime="+93" swimtime="00:03:15.01" resultid="5283" heatid="7335" lane="7" entrytime="00:03:25.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:33.26" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="302" reactiontime="+91" swimtime="00:01:14.86" resultid="5284" heatid="7383" lane="2" entrytime="00:01:16.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="279" swimtime="00:00:33.25" resultid="5285" heatid="7442" lane="1" entrytime="00:00:32.90" />
                <RESULT eventid="1577" points="212" reactiontime="+97" swimtime="00:06:34.79" resultid="5286" heatid="8156" lane="3" entrytime="00:06:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:02:23.27" />
                    <SPLIT distance="200" swimtime="00:03:13.20" />
                    <SPLIT distance="250" swimtime="00:04:09.75" />
                    <SPLIT distance="300" swimtime="00:05:06.10" />
                    <SPLIT distance="350" swimtime="00:05:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="215" reactiontime="+84" swimtime="00:02:56.19" resultid="5287" heatid="7533" lane="9" entrytime="00:03:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:12.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="256" reactiontime="+92" swimtime="00:05:34.19" resultid="5288" heatid="7579" lane="0" entrytime="00:05:54.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                    <SPLIT distance="150" swimtime="00:02:02.90" />
                    <SPLIT distance="200" swimtime="00:02:45.21" />
                    <SPLIT distance="250" swimtime="00:03:28.15" />
                    <SPLIT distance="300" swimtime="00:04:10.56" />
                    <SPLIT distance="350" swimtime="00:04:52.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PKZÁ" nation="CZE" clubid="2658" name="Plavecký klub Zábřeh">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-26" firstname="David" gender="M" lastname="Kochwasser" nation="CZE" athleteid="2657">
              <RESULTS>
                <RESULT eventid="1076" points="382" swimtime="00:00:27.91" resultid="2659" heatid="7260" lane="0" entrytime="00:00:28.77" />
                <RESULT eventid="1288" points="373" reactiontime="+73" swimtime="00:01:02.41" resultid="2660" heatid="7360" lane="1" entrytime="00:01:03.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="387" reactiontime="+72" swimtime="00:01:16.25" resultid="2661" heatid="7423" lane="5" entrytime="00:01:17.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="345" reactiontime="+72" swimtime="00:00:30.99" resultid="2662" heatid="7443" lane="3" entrytime="00:00:31.29" />
                <RESULT eventid="1625" points="256" reactiontime="+73" swimtime="00:01:15.67" resultid="2663" heatid="7518" lane="1" entrytime="00:01:14.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="402" reactiontime="+70" swimtime="00:00:34.21" resultid="2664" heatid="7559" lane="2" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-19" firstname="Jiri" gender="M" lastname="Sip" nation="CZE" athleteid="2665">
              <RESULTS>
                <RESULT eventid="1076" points="444" reactiontime="+87" swimtime="00:00:26.55" resultid="2666" heatid="7265" lane="4" entrytime="00:00:26.75" />
                <RESULT eventid="1108" points="429" reactiontime="+89" swimtime="00:02:25.31" resultid="2667" heatid="7283" lane="4" entrytime="00:02:26.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="373" reactiontime="+71" swimtime="00:00:30.86" resultid="2668" heatid="7325" lane="0" entrytime="00:00:31.17" />
                <RESULT eventid="1320" points="449" reactiontime="+85" swimtime="00:01:05.60" resultid="2669" heatid="7388" lane="2" entrytime="00:01:06.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="394" reactiontime="+68" swimtime="00:01:06.65" resultid="2670" heatid="7466" lane="1" entrytime="00:01:07.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="391" reactiontime="+93" swimtime="00:05:22.02" resultid="2671" heatid="8158" lane="8" entrytime="00:05:21.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="200" swimtime="00:02:37.57" />
                    <SPLIT distance="250" swimtime="00:03:24.51" />
                    <SPLIT distance="300" swimtime="00:04:10.93" />
                    <SPLIT distance="350" swimtime="00:04:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="367" reactiontime="+71" swimtime="00:02:27.43" resultid="2672" heatid="7535" lane="1" entrytime="00:02:29.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-04-23" firstname="Pavlína" gender="F" lastname="Troblová" nation="CZE" athleteid="2673">
              <RESULTS>
                <RESULT eventid="1059" points="351" reactiontime="+91" swimtime="00:00:32.49" resultid="2674" heatid="7240" lane="4" entrytime="00:00:33.11" />
                <RESULT eventid="1272" points="332" reactiontime="+77" swimtime="00:01:12.54" resultid="2675" heatid="7345" lane="2" entrytime="00:01:12.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="321" reactiontime="+92" swimtime="00:01:22.47" resultid="2676" heatid="7373" lane="8" entrytime="00:01:24.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="265" reactiontime="+83" swimtime="00:01:37.02" resultid="2677" heatid="7411" lane="2" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="283" reactiontime="+83" swimtime="00:01:23.81" resultid="2678" heatid="7456" lane="7" entrytime="00:01:24.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="291" reactiontime="+74" swimtime="00:00:43.08" resultid="2679" heatid="7541" lane="0" entrytime="00:00:45.60" />
                <RESULT eventid="1721" points="315" reactiontime="+79" swimtime="00:05:43.55" resultid="2680" heatid="7568" lane="4" entrytime="00:05:45.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                    <SPLIT distance="200" swimtime="00:02:45.86" />
                    <SPLIT distance="250" swimtime="00:03:30.71" />
                    <SPLIT distance="300" swimtime="00:04:16.17" />
                    <SPLIT distance="350" swimtime="00:05:00.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PSWRO" nation="POL" region="01" clubid="3726" name="Power Swimming Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1991-02-10" firstname="Jacek" gender="M" lastname="Sokulski" nation="POL" athleteid="3725">
              <RESULTS>
                <RESULT eventid="1076" points="665" reactiontime="+77" swimtime="00:00:23.21" resultid="3727" heatid="7270" lane="1" entrytime="00:00:24.00" />
                <RESULT eventid="1288" points="685" reactiontime="+65" swimtime="00:00:50.97" resultid="3728" heatid="7349" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="581" reactiontime="+68" swimtime="00:01:00.23" resultid="3729" heatid="7389" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="695" reactiontime="+67" swimtime="00:00:24.55" resultid="3730" heatid="7451" lane="3" entrytime="00:00:24.80" />
                <RESULT eventid="1513" points="610" reactiontime="+72" swimtime="00:01:57.11" resultid="3731" heatid="7488" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="100" swimtime="00:00:57.39" />
                    <SPLIT distance="150" swimtime="00:01:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="605" reactiontime="+71" swimtime="00:00:56.84" resultid="3732" heatid="7522" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="497" reactiontime="+61" swimtime="00:04:27.80" resultid="3733" heatid="7573" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="150" swimtime="00:01:36.61" />
                    <SPLIT distance="200" swimtime="00:02:11.73" />
                    <SPLIT distance="250" swimtime="00:02:47.48" />
                    <SPLIT distance="300" swimtime="00:03:22.72" />
                    <SPLIT distance="350" swimtime="00:03:55.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-12-04" firstname="Angelika" gender="F" lastname="Wróbel" nation="POL" athleteid="3734">
              <RESULTS>
                <RESULT eventid="1059" points="574" reactiontime="+86" swimtime="00:00:27.58" resultid="3735" heatid="7245" lane="3" entrytime="00:00:27.43" />
                <RESULT eventid="1272" points="565" reactiontime="+87" swimtime="00:01:00.75" resultid="3736" heatid="7348" lane="0" entrytime="00:01:00.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="536" reactiontime="+86" swimtime="00:02:15.89" resultid="3737" heatid="7474" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PRKAL" nation="RUS" clubid="5796" name="Pregel Kaliningrad">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Elena" gender="F" lastname="Dautova" nation="RUS" athleteid="5802">
              <RESULTS>
                <RESULT eventid="1059" points="378" reactiontime="+87" swimtime="00:00:31.71" resultid="5803" heatid="7242" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1207" points="329" reactiontime="+70" swimtime="00:00:37.15" resultid="5804" heatid="7311" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1272" points="343" reactiontime="+82" swimtime="00:01:11.73" resultid="5805" heatid="7345" lane="3" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="263" reactiontime="+83" swimtime="00:01:25.83" resultid="5806" heatid="7455" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="5816">
              <RESULTS>
                <RESULT eventid="1108" points="253" reactiontime="+65" swimtime="00:02:53.21" resultid="5817" heatid="7281" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="294" reactiontime="+81" swimtime="00:21:15.11" resultid="5818" heatid="7303" lane="6" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:05.06" />
                    <SPLIT distance="200" swimtime="00:02:48.53" />
                    <SPLIT distance="250" swimtime="00:03:32.18" />
                    <SPLIT distance="300" swimtime="00:04:15.67" />
                    <SPLIT distance="350" swimtime="00:04:59.74" />
                    <SPLIT distance="400" swimtime="00:05:42.87" />
                    <SPLIT distance="450" swimtime="00:06:26.13" />
                    <SPLIT distance="500" swimtime="00:07:09.78" />
                    <SPLIT distance="550" swimtime="00:07:52.45" />
                    <SPLIT distance="600" swimtime="00:08:35.26" />
                    <SPLIT distance="650" swimtime="00:09:18.28" />
                    <SPLIT distance="700" swimtime="00:10:01.30" />
                    <SPLIT distance="750" swimtime="00:10:44.66" />
                    <SPLIT distance="800" swimtime="00:11:27.44" />
                    <SPLIT distance="850" swimtime="00:12:09.99" />
                    <SPLIT distance="900" swimtime="00:12:52.44" />
                    <SPLIT distance="950" swimtime="00:13:34.91" />
                    <SPLIT distance="1000" swimtime="00:14:17.37" />
                    <SPLIT distance="1050" swimtime="00:14:59.18" />
                    <SPLIT distance="1100" swimtime="00:15:41.17" />
                    <SPLIT distance="1150" swimtime="00:16:23.21" />
                    <SPLIT distance="1200" swimtime="00:17:05.86" />
                    <SPLIT distance="1250" swimtime="00:17:48.09" />
                    <SPLIT distance="1300" swimtime="00:18:31.09" />
                    <SPLIT distance="1350" swimtime="00:19:13.11" />
                    <SPLIT distance="1400" swimtime="00:19:55.15" />
                    <SPLIT distance="1450" swimtime="00:20:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="284" reactiontime="+68" swimtime="00:01:08.36" resultid="5819" heatid="7357" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="265" reactiontime="+70" swimtime="00:01:18.24" resultid="5820" heatid="7383" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="292" reactiontime="+67" swimtime="00:01:23.79" resultid="5821" heatid="7420" lane="4" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="288" reactiontime="+66" swimtime="00:02:30.43" resultid="5822" heatid="7481" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5823" heatid="7555" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5824" heatid="7577" lane="8" entrytime="00:05:19.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="5807">
              <RESULTS>
                <RESULT eventid="1059" points="639" reactiontime="+83" swimtime="00:00:26.61" resultid="5808" heatid="7245" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="1272" points="632" reactiontime="+81" swimtime="00:00:58.53" resultid="5809" heatid="7348" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="525" reactiontime="+85" swimtime="00:00:30.21" resultid="5810" heatid="7433" lane="5" entrytime="00:00:30.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="5811">
              <RESULTS>
                <RESULT eventid="1076" points="198" swimtime="00:00:34.74" resultid="5812" heatid="7252" lane="8" entrytime="00:00:35.80" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="5813" heatid="7319" lane="9" entrytime="00:00:44.80" />
                <RESULT eventid="1417" points="181" reactiontime="+94" swimtime="00:01:38.14" resultid="5814" heatid="7417" lane="3" entrytime="00:01:42.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5815" heatid="7550" lane="7" entrytime="00:00:43.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="5795">
              <RESULTS>
                <RESULT eventid="1059" points="285" reactiontime="+92" swimtime="00:00:34.84" resultid="5797" heatid="7239" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1207" points="203" reactiontime="+80" swimtime="00:00:43.61" resultid="5798" heatid="7309" lane="5" entrytime="00:00:44.50" />
                <RESULT eventid="1272" points="295" reactiontime="+91" swimtime="00:01:15.46" resultid="5799" heatid="7344" lane="0" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="315" reactiontime="+71" swimtime="00:02:42.15" resultid="5800" heatid="7471" lane="3" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:19.04" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="308" reactiontime="+77" swimtime="00:05:46.33" resultid="5801" heatid="7568" lane="5" entrytime="00:05:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:06.48" />
                    <SPLIT distance="200" swimtime="00:02:51.18" />
                    <SPLIT distance="250" swimtime="00:03:35.78" />
                    <SPLIT distance="300" swimtime="00:04:20.22" />
                    <SPLIT distance="350" swimtime="00:05:04.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="328" reactiontime="+90" swimtime="00:02:07.35" resultid="6869" heatid="7287" lane="4" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:34.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5795" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="5816" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5807" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="5811" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="PLOLE" nation="POL" region="01" clubid="2444" name="Pływak Oleśnica">
          <ATHLETES>
            <ATHLETE birthdate="1980-02-06" firstname="Marcin" gender="M" lastname="Hejninger" nation="POL" athleteid="2443">
              <RESULTS>
                <RESULT eventid="1076" points="205" reactiontime="+90" swimtime="00:00:34.33" resultid="2445" heatid="7251" lane="3" entrytime="00:00:36.82" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2446" heatid="7276" lane="5" />
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu. (Time: 10:36)" eventid="1256" reactiontime="+87" status="DSQ" swimtime="00:03:33.19" resultid="2447" heatid="7334" lane="0" entrytime="00:03:58.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="194" reactiontime="+97" swimtime="00:01:17.62" resultid="2448" heatid="7351" lane="6" entrytime="00:01:35.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="208" reactiontime="+77" swimtime="00:01:33.76" resultid="2449" heatid="7417" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2450" heatid="7435" lane="5" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="2451" heatid="7512" lane="1" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2452" heatid="7549" lane="7" entrytime="00:00:47.11" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01911" nation="POL" region="11" clubid="2437" name="RMKS Rybnik">
          <CONTACT city="Rybnik" email="piotrandrosz992@gmail.com" name="Androsz" phone="504013886" state="SLA" street="Powstańców Sl. 40/42" zip="44-200" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" license="101911600104" athleteid="2438">
              <RESULTS>
                <RESULT eventid="1059" points="551" reactiontime="+71" swimtime="00:00:27.96" resultid="2439" heatid="7245" lane="8" entrytime="00:00:27.70" />
                <RESULT eventid="1092" points="433" swimtime="00:02:41.00" resultid="2440" heatid="7275" lane="0" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="498" reactiontime="+74" swimtime="00:01:03.37" resultid="2441" heatid="7347" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="544" reactiontime="+71" swimtime="00:00:29.85" resultid="2442" heatid="7434" lane="6" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-01" firstname="Szymon" gender="M" lastname="Lindner" nation="POL" license="501911700158" athleteid="4394">
              <RESULTS>
                <RESULT eventid="1076" points="566" reactiontime="+78" swimtime="00:00:24.49" resultid="4395" heatid="7246" lane="4" />
                <RESULT eventid="1108" points="494" reactiontime="+73" swimtime="00:02:18.67" resultid="4396" heatid="7277" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="547" reactiontime="+72" swimtime="00:00:54.95" resultid="4397" heatid="7365" lane="6" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="491" reactiontime="+73" swimtime="00:01:03.70" resultid="4398" heatid="7377" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="533" reactiontime="+72" swimtime="00:02:02.50" resultid="4399" heatid="7486" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="150" swimtime="00:01:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="476" reactiontime="+82" swimtime="00:05:01.48" resultid="4400" heatid="8153" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                    <SPLIT distance="200" swimtime="00:02:28.25" />
                    <SPLIT distance="250" swimtime="00:03:11.69" />
                    <SPLIT distance="300" swimtime="00:03:54.51" />
                    <SPLIT distance="350" swimtime="00:04:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="376" reactiontime="+79" swimtime="00:02:26.31" resultid="4401" heatid="7529" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="499" reactiontime="+78" swimtime="00:04:27.59" resultid="4402" heatid="7574" lane="6" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="150" swimtime="00:01:36.82" />
                    <SPLIT distance="200" swimtime="00:02:11.38" />
                    <SPLIT distance="250" swimtime="00:02:46.12" />
                    <SPLIT distance="300" swimtime="00:03:20.82" />
                    <SPLIT distance="350" swimtime="00:03:55.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ROYAL" nation="SVK" region="BAO" clubid="2905" name="Royal plavecký klub Bratislava" shortname="Royal Bratislava">
          <CONTACT city="Bratislava" email="schild@royalclub.sk" name="Schild Igor" phone="0911175865" street="Iľjušinová 6" zip="85101" />
          <ATHLETES>
            <ATHLETE birthdate="1991-03-13" firstname="Peter" gender="M" lastname="Hrinda" nation="SVK" license="SVK11097" athleteid="2906">
              <RESULTS>
                <RESULT eventid="1076" points="526" reactiontime="+68" swimtime="00:00:25.09" resultid="2907" heatid="7269" lane="2" entrytime="00:00:24.98" entrycourse="SCM" />
                <RESULT eventid="1288" points="495" reactiontime="+72" swimtime="00:00:56.80" resultid="2908" heatid="7366" lane="3" entrytime="00:00:55.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="521" reactiontime="+65" swimtime="00:00:27.03" resultid="2909" heatid="7450" lane="7" entrytime="00:00:26.67" entrycourse="SCM" />
                <RESULT eventid="1689" points="638" reactiontime="+63" swimtime="00:00:29.33" resultid="2910" heatid="7561" lane="7" entrytime="00:00:29.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03706" nation="POL" region="06" clubid="2650" name="Siemacha Kraków">
          <CONTACT name="Joanna Kwatera" phone="790611187" />
          <ATHLETES>
            <ATHLETE birthdate="1980-01-08" firstname="Karolina" gender="F" lastname="Spuła" nation="POL" athleteid="2651">
              <RESULTS>
                <RESULT eventid="1059" points="139" swimtime="00:00:44.24" resultid="2652" heatid="7236" lane="0" entrytime="00:00:49.00" />
                <RESULT eventid="1272" points="105" reactiontime="+91" swimtime="00:01:46.22" resultid="2653" heatid="7341" lane="3" entrytime="00:01:48.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03111" nation="POL" region="11" clubid="4144" name="Sikret Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@tlen.pl" internet="https://www.facebook.com/joanna.sikret" name="Joanna Zagała" phone="693651233" state="ŚLĄSK" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="4145">
              <RESULTS>
                <RESULT eventid="1059" points="158" swimtime="00:00:42.37" resultid="4146" heatid="7237" lane="0" entrytime="00:00:43.00" />
                <RESULT eventid="1140" points="135" swimtime="00:15:33.91" resultid="4147" heatid="7292" lane="0" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:45.28" />
                    <SPLIT distance="150" swimtime="00:02:44.77" />
                    <SPLIT distance="200" swimtime="00:03:43.32" />
                    <SPLIT distance="250" swimtime="00:04:41.90" />
                    <SPLIT distance="300" swimtime="00:05:41.15" />
                    <SPLIT distance="350" swimtime="00:06:40.17" />
                    <SPLIT distance="400" swimtime="00:07:39.40" />
                    <SPLIT distance="450" swimtime="00:08:38.37" />
                    <SPLIT distance="500" swimtime="00:09:37.69" />
                    <SPLIT distance="550" swimtime="00:10:38.02" />
                    <SPLIT distance="600" swimtime="00:11:37.21" />
                    <SPLIT distance="650" swimtime="00:12:36.00" />
                    <SPLIT distance="700" swimtime="00:13:36.09" />
                    <SPLIT distance="750" swimtime="00:14:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="141" reactiontime="+90" swimtime="00:04:18.15" resultid="4148" heatid="7328" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.12" />
                    <SPLIT distance="100" swimtime="00:02:06.12" />
                    <SPLIT distance="150" swimtime="00:03:13.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="116" reactiontime="+87" swimtime="00:01:55.55" resultid="4149" heatid="7369" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="135" reactiontime="+88" swimtime="00:02:01.42" resultid="4150" heatid="7409" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="99" reactiontime="+97" swimtime="00:09:18.26" resultid="4151" heatid="8149" lane="7" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.74" />
                    <SPLIT distance="100" swimtime="00:02:20.53" />
                    <SPLIT distance="150" swimtime="00:03:41.24" />
                    <SPLIT distance="200" swimtime="00:04:56.63" />
                    <SPLIT distance="250" swimtime="00:06:09.84" />
                    <SPLIT distance="300" swimtime="00:07:21.86" />
                    <SPLIT distance="350" swimtime="00:08:21.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="72" reactiontime="+82" swimtime="00:02:10.93" resultid="4152" heatid="7507" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="179" reactiontime="+86" swimtime="00:00:50.64" resultid="4153" heatid="7538" lane="6" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-04-20" firstname="Wojciech" gender="M" lastname="Kosiak" nation="POL" athleteid="4169">
              <RESULTS>
                <RESULT eventid="1076" points="110" swimtime="00:00:42.27" resultid="4170" heatid="7249" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1288" points="93" swimtime="00:01:38.89" resultid="4171" heatid="7351" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="68" swimtime="00:00:53.28" resultid="4172" heatid="7437" lane="0" entrytime="00:00:52.00" />
                <RESULT eventid="1513" points="80" swimtime="00:03:49.91" resultid="4173" heatid="7476" lane="2" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:54.43" />
                    <SPLIT distance="150" swimtime="00:02:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="81" swimtime="00:08:10.50" resultid="4174" heatid="7583" lane="3" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.54" />
                    <SPLIT distance="100" swimtime="00:02:00.28" />
                    <SPLIT distance="150" swimtime="00:03:04.87" />
                    <SPLIT distance="200" swimtime="00:04:07.31" />
                    <SPLIT distance="250" swimtime="00:05:10.65" />
                    <SPLIT distance="300" swimtime="00:06:12.96" />
                    <SPLIT distance="350" swimtime="00:07:16.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="4154">
              <RESULTS>
                <RESULT eventid="1076" points="178" reactiontime="+94" swimtime="00:00:36.00" resultid="4155" heatid="7252" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1108" points="144" swimtime="00:03:28.93" resultid="4156" heatid="7279" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:02:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="137" reactiontime="+77" swimtime="00:00:43.02" resultid="4157" heatid="7319" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1288" points="191" swimtime="00:01:17.97" resultid="4158" heatid="7353" lane="8" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="142" reactiontime="+77" swimtime="00:01:33.49" resultid="4159" heatid="7461" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="178" reactiontime="+98" swimtime="00:02:56.54" resultid="4160" heatid="7477" lane="3" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:22.14" />
                    <SPLIT distance="150" swimtime="00:02:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="126" reactiontime="+76" swimtime="00:03:30.69" resultid="4161" heatid="7531" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="100" swimtime="00:01:41.33" />
                    <SPLIT distance="150" swimtime="00:02:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="170" reactiontime="+98" swimtime="00:06:22.79" resultid="4162" heatid="7582" lane="3" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:02:14.59" />
                    <SPLIT distance="200" swimtime="00:03:04.56" />
                    <SPLIT distance="250" swimtime="00:03:55.01" />
                    <SPLIT distance="300" swimtime="00:04:45.39" />
                    <SPLIT distance="350" swimtime="00:05:35.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="4175">
              <RESULTS>
                <RESULT eventid="1108" points="268" reactiontime="+84" swimtime="00:02:50.04" resultid="4176" heatid="7281" lane="8" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:02:08.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="282" reactiontime="+73" swimtime="00:00:33.88" resultid="4177" heatid="7323" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1449" points="378" reactiontime="+82" swimtime="00:00:30.06" resultid="4178" heatid="7443" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1481" points="278" reactiontime="+75" swimtime="00:01:14.86" resultid="4179" heatid="7463" lane="5" entrytime="00:01:20.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="324" reactiontime="+78" swimtime="00:01:09.99" resultid="4180" heatid="7516" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="274" reactiontime="+76" swimtime="00:05:26.66" resultid="4181" heatid="7579" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.62" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                    <SPLIT distance="200" swimtime="00:02:37.32" />
                    <SPLIT distance="250" swimtime="00:03:19.54" />
                    <SPLIT distance="300" swimtime="00:04:02.34" />
                    <SPLIT distance="350" swimtime="00:04:45.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-14" firstname="Teresa" gender="F" lastname="Żylińska" nation="POL" athleteid="4163">
              <RESULTS>
                <RESULT eventid="1059" points="82" reactiontime="+90" swimtime="00:00:52.66" resultid="4164" heatid="7235" lane="5" entrytime="00:00:52.00" />
                <RESULT eventid="1207" points="79" reactiontime="+71" swimtime="00:00:59.82" resultid="4165" heatid="7307" lane="3" entrytime="00:01:02.00" />
                <RESULT eventid="1272" points="69" swimtime="00:02:02.08" resultid="4166" heatid="7340" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="70" reactiontime="+73" swimtime="00:02:13.42" resultid="4167" heatid="7453" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="72" reactiontime="+71" swimtime="00:04:45.47" resultid="4168" heatid="7524" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.26" />
                    <SPLIT distance="100" swimtime="00:02:18.25" />
                    <SPLIT distance="150" swimtime="00:03:34.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="135" reactiontime="+85" swimtime="00:02:51.18" resultid="4182" heatid="7287" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:01:27.80" />
                    <SPLIT distance="150" swimtime="00:02:21.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4145" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4169" number="2" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4163" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4175" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" status="DNS" swimtime="00:00:00.00" resultid="4183" heatid="7563" lane="0" entrytime="00:03:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4175" number="1" />
                    <RELAYPOSITION athleteid="4145" number="2" />
                    <RELAYPOSITION athleteid="4169" number="3" />
                    <RELAYPOSITION athleteid="4163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="14" clubid="2949" name="SKP Legia Warszawa" shortname="Legia Warszawa">
          <CONTACT name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1993-03-26" firstname="Adrianna" gender="F" lastname="Borowa" nation="POL" athleteid="3026">
              <RESULTS>
                <RESULT eventid="1465" points="235" reactiontime="+79" swimtime="00:01:29.12" resultid="3027" heatid="7455" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="5775">
              <RESULTS>
                <RESULT eventid="1076" points="215" reactiontime="+85" swimtime="00:00:33.80" resultid="5776" heatid="7254" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1188" points="180" reactiontime="+94" swimtime="00:25:00.56" resultid="5777" heatid="7304" lane="8" entrytime="00:27:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:30.65" />
                    <SPLIT distance="150" swimtime="00:02:20.68" />
                    <SPLIT distance="200" swimtime="00:03:10.49" />
                    <SPLIT distance="250" swimtime="00:04:00.21" />
                    <SPLIT distance="300" swimtime="00:04:50.64" />
                    <SPLIT distance="350" swimtime="00:05:40.42" />
                    <SPLIT distance="400" swimtime="00:06:31.14" />
                    <SPLIT distance="450" swimtime="00:07:22.53" />
                    <SPLIT distance="500" swimtime="00:08:13.69" />
                    <SPLIT distance="550" swimtime="00:09:03.89" />
                    <SPLIT distance="600" swimtime="00:09:53.90" />
                    <SPLIT distance="650" swimtime="00:10:45.08" />
                    <SPLIT distance="700" swimtime="00:11:35.92" />
                    <SPLIT distance="750" swimtime="00:12:26.56" />
                    <SPLIT distance="800" swimtime="00:13:17.33" />
                    <SPLIT distance="850" swimtime="00:14:09.36" />
                    <SPLIT distance="900" swimtime="00:15:00.43" />
                    <SPLIT distance="950" swimtime="00:15:51.95" />
                    <SPLIT distance="1000" swimtime="00:16:43.03" />
                    <SPLIT distance="1050" swimtime="00:17:32.90" />
                    <SPLIT distance="1100" swimtime="00:18:23.54" />
                    <SPLIT distance="1150" swimtime="00:19:13.87" />
                    <SPLIT distance="1200" swimtime="00:20:05.81" />
                    <SPLIT distance="1250" swimtime="00:20:56.06" />
                    <SPLIT distance="1300" swimtime="00:21:46.56" />
                    <SPLIT distance="1350" swimtime="00:22:37.44" />
                    <SPLIT distance="1400" swimtime="00:23:27.45" />
                    <SPLIT distance="1450" swimtime="00:24:17.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="172" reactiontime="+81" swimtime="00:00:39.91" resultid="5778" heatid="7319" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1352" points="83" reactiontime="+86" swimtime="00:04:08.01" resultid="5779" heatid="7395" lane="1" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                    <SPLIT distance="100" swimtime="00:01:54.50" />
                    <SPLIT distance="150" swimtime="00:03:01.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="147" reactiontime="+83" swimtime="00:01:32.53" resultid="5780" heatid="7462" lane="2" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="132" swimtime="00:07:41.99" resultid="5781" heatid="8155" lane="0" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                    <SPLIT distance="100" swimtime="00:01:56.25" />
                    <SPLIT distance="150" swimtime="00:02:54.78" />
                    <SPLIT distance="200" swimtime="00:03:50.25" />
                    <SPLIT distance="250" swimtime="00:05:02.81" />
                    <SPLIT distance="300" swimtime="00:06:09.29" />
                    <SPLIT distance="350" swimtime="00:06:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="104" reactiontime="+97" swimtime="00:03:44.53" resultid="5782" heatid="7531" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                    <SPLIT distance="100" swimtime="00:01:49.12" />
                    <SPLIT distance="150" swimtime="00:02:48.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="190" reactiontime="+92" swimtime="00:06:08.58" resultid="5783" heatid="7581" lane="0" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:26.20" />
                    <SPLIT distance="150" swimtime="00:02:13.17" />
                    <SPLIT distance="200" swimtime="00:03:01.45" />
                    <SPLIT distance="250" swimtime="00:03:49.00" />
                    <SPLIT distance="300" swimtime="00:04:36.79" />
                    <SPLIT distance="350" swimtime="00:05:24.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-01" firstname="Stanisław" gender="M" lastname="Fluder" nation="POL" athleteid="2973">
              <RESULTS>
                <RESULT eventid="1076" points="503" swimtime="00:00:25.46" resultid="2974" heatid="7264" lane="0" entrytime="00:00:27.09" />
                <RESULT comment="Rekord Polski Masters kategoria B" eventid="1188" points="527" reactiontime="+85" swimtime="00:17:29.67" resultid="2975" heatid="7302" lane="3" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                    <SPLIT distance="200" swimtime="00:02:16.34" />
                    <SPLIT distance="250" swimtime="00:02:51.84" />
                    <SPLIT distance="300" swimtime="00:03:27.47" />
                    <SPLIT distance="350" swimtime="00:04:03.11" />
                    <SPLIT distance="400" swimtime="00:04:38.27" />
                    <SPLIT distance="450" swimtime="00:05:13.42" />
                    <SPLIT distance="500" swimtime="00:05:48.66" />
                    <SPLIT distance="550" swimtime="00:06:23.57" />
                    <SPLIT distance="600" swimtime="00:06:58.54" />
                    <SPLIT distance="650" swimtime="00:07:33.34" />
                    <SPLIT distance="700" swimtime="00:08:08.20" />
                    <SPLIT distance="750" swimtime="00:08:43.28" />
                    <SPLIT distance="800" swimtime="00:09:18.65" />
                    <SPLIT distance="850" swimtime="00:09:54.07" />
                    <SPLIT distance="900" swimtime="00:10:29.55" />
                    <SPLIT distance="950" swimtime="00:11:05.27" />
                    <SPLIT distance="1000" swimtime="00:11:40.98" />
                    <SPLIT distance="1050" swimtime="00:12:16.49" />
                    <SPLIT distance="1100" swimtime="00:12:51.39" />
                    <SPLIT distance="1150" swimtime="00:13:26.76" />
                    <SPLIT distance="1200" swimtime="00:14:02.06" />
                    <SPLIT distance="1250" swimtime="00:14:37.38" />
                    <SPLIT distance="1300" swimtime="00:15:12.42" />
                    <SPLIT distance="1350" swimtime="00:15:47.54" />
                    <SPLIT distance="1400" swimtime="00:16:22.64" />
                    <SPLIT distance="1450" swimtime="00:16:57.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="549" reactiontime="+72" swimtime="00:00:54.88" resultid="2976" heatid="7364" lane="7" entrytime="00:00:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="488" reactiontime="+72" swimtime="00:00:27.61" resultid="2977" heatid="7446" lane="3" entrytime="00:00:29.20" />
                <RESULT eventid="1513" points="557" reactiontime="+72" swimtime="00:02:00.71" resultid="2978" heatid="7486" lane="5" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:00:59.05" />
                    <SPLIT distance="150" swimtime="00:01:30.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-25" firstname="Adrian" gender="M" lastname="Jagodziński" nation="POL" athleteid="2986">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2987" heatid="7264" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1449" points="282" swimtime="00:00:33.13" resultid="2988" heatid="7441" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="3002">
              <RESULTS>
                <RESULT eventid="1207" points="519" reactiontime="+68" swimtime="00:00:31.94" resultid="3003" heatid="7314" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="3004" heatid="7376" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="1465" points="508" reactiontime="+72" swimtime="00:01:08.95" resultid="3005" heatid="7458" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="452" reactiontime="+84" swimtime="00:05:37.40" resultid="3006" heatid="8151" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:16.95" />
                    <SPLIT distance="150" swimtime="00:01:57.92" />
                    <SPLIT distance="200" swimtime="00:02:40.55" />
                    <SPLIT distance="250" swimtime="00:03:27.58" />
                    <SPLIT distance="300" swimtime="00:04:15.88" />
                    <SPLIT distance="350" swimtime="00:04:57.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="468" reactiontime="+75" swimtime="00:02:33.56" resultid="3007" heatid="7528" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="3008" heatid="7544" lane="4" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="2992">
              <RESULTS>
                <RESULT eventid="1076" points="586" reactiontime="+86" swimtime="00:00:24.20" resultid="2993" heatid="7270" lane="7" entrytime="00:00:23.99" />
                <RESULT eventid="1224" points="633" reactiontime="+63" swimtime="00:00:25.87" resultid="2994" heatid="7326" lane="4" entrytime="00:00:25.99" />
                <RESULT eventid="1449" points="671" reactiontime="+75" swimtime="00:00:24.84" resultid="2995" heatid="7436" lane="0" />
                <RESULT comment="Rekord Europy Masters kategoria D" eventid="1481" points="641" reactiontime="+63" swimtime="00:00:56.69" resultid="2996" heatid="7467" lane="4" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="626" reactiontime="+73" swimtime="00:00:56.20" resultid="2997" heatid="7522" lane="5" entrytime="00:00:55.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-16" firstname="Jacek" gender="M" lastname="Kaczyński" nation="POL" athleteid="2955">
              <RESULTS>
                <RESULT eventid="1076" points="594" reactiontime="+87" swimtime="00:00:24.10" resultid="2956" heatid="7270" lane="8" entrytime="00:00:24.00" />
                <RESULT eventid="1449" points="580" reactiontime="+68" swimtime="00:00:26.07" resultid="2957" heatid="7450" lane="5" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-27" firstname="Agata" gender="F" lastname="Korc" nation="POL" athleteid="2989">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2990" heatid="7245" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="2991" heatid="7434" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-05-18" firstname="Marcin" gender="M" lastname="Kozłowski" nation="POL" athleteid="3014">
              <RESULTS>
                <RESULT eventid="1076" points="522" reactiontime="+84" swimtime="00:00:25.15" resultid="3015" heatid="7247" lane="9" />
                <RESULT eventid="1288" points="477" reactiontime="+75" swimtime="00:00:57.50" resultid="3016" heatid="7349" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="467" reactiontime="+76" swimtime="00:00:28.03" resultid="3017" heatid="7436" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-13" firstname="Romuald" gender="M" lastname="Kozłowski" nation="POL" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1076" points="396" reactiontime="+81" swimtime="00:00:27.58" resultid="3010" heatid="7262" lane="8" entrytime="00:00:28.00" />
                <RESULT comment="Rekord Polski Masters kategoria F" eventid="1256" points="385" reactiontime="+73" swimtime="00:02:45.17" resultid="3011" heatid="7337" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Roekord Polski Masters kategeria F" eventid="1417" points="463" reactiontime="+74" swimtime="00:01:11.88" resultid="3012" heatid="7424" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria F" eventid="1689" points="456" reactiontime="+69" swimtime="00:00:32.79" resultid="3013" heatid="7558" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1320" points="396" reactiontime="+72" swimtime="00:01:08.43" resultid="6479" heatid="7386" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-15" firstname="Aleksandra" gender="F" lastname="Marianek" nation="POL" athleteid="3023">
              <RESULTS>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="3024" heatid="7291" lane="4" entrytime="00:12:00.00" />
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="3025" heatid="7331" lane="1" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-04" firstname="Hubert" gender="M" lastname="Markowski" nation="POL" athleteid="2998">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2999" heatid="7282" lane="6" entrytime="00:02:37.00" />
                <RESULT eventid="1625" points="349" reactiontime="+82" swimtime="00:01:08.27" resultid="3000" heatid="7519" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="303" reactiontime="+72" swimtime="00:02:37.20" resultid="3001" heatid="7534" lane="0" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="150" swimtime="00:01:58.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-27" firstname="Jan" gender="M" lastname="Peńsko" nation="POL" athleteid="2967">
              <RESULTS>
                <RESULT eventid="1449" points="492" reactiontime="+73" swimtime="00:00:27.55" resultid="2968" heatid="7449" lane="7" entrytime="00:00:27.49" />
                <RESULT eventid="1481" points="476" reactiontime="+74" swimtime="00:01:02.59" resultid="2969" heatid="7467" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="510" reactiontime="+81" swimtime="00:01:00.17" resultid="2970" heatid="7522" lane="3" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-12" firstname="Jan" gender="M" lastname="Rekowski" nation="POL" athleteid="3018">
              <RESULTS>
                <RESULT eventid="1076" points="456" reactiontime="+83" swimtime="00:00:26.32" resultid="3019" heatid="7266" lane="6" entrytime="00:00:26.30" />
                <RESULT eventid="1288" points="418" reactiontime="+99" swimtime="00:01:00.06" resultid="3020" heatid="7363" lane="9" entrytime="00:00:59.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="343" reactiontime="+94" swimtime="00:01:11.79" resultid="3021" heatid="7385" lane="8" entrytime="00:01:12.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="381" reactiontime="+92" swimtime="00:00:29.98" resultid="3022" heatid="7446" lane="0" entrytime="00:00:29.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="2958">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2959" heatid="7269" lane="6" entrytime="00:00:24.96" />
                <RESULT eventid="1417" points="589" reactiontime="+70" swimtime="00:01:06.34" resultid="2960" heatid="7425" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="516" reactiontime="+69" swimtime="00:00:27.11" resultid="2961" heatid="7450" lane="1" entrytime="00:00:26.69" />
                <RESULT eventid="1689" points="590" reactiontime="+69" swimtime="00:00:30.09" resultid="2962" heatid="7561" lane="2" entrytime="00:00:28.80" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="5945" heatid="7512" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Maciej" gender="M" lastname="Rybicki" nation="POL" athleteid="2971">
              <RESULTS>
                <RESULT eventid="1076" points="284" reactiontime="+79" swimtime="00:00:30.81" resultid="2972" heatid="7257" lane="7" entrytime="00:00:30.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-04" firstname="Marcin" gender="M" lastname="Walkowicz" nation="POL" athleteid="2984">
              <RESULTS>
                <RESULT eventid="1076" points="223" reactiontime="+84" swimtime="00:00:33.36" resultid="2985" heatid="7255" lane="2" entrytime="00:00:32.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="2963">
              <RESULTS>
                <RESULT eventid="1076" points="465" reactiontime="+76" swimtime="00:00:26.14" resultid="2964" heatid="7266" lane="5" entrytime="00:00:26.25" />
                <RESULT eventid="1288" points="480" reactiontime="+73" swimtime="00:00:57.38" resultid="2965" heatid="7363" lane="1" entrytime="00:00:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2966" heatid="7446" lane="8" entrytime="00:00:29.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="2950">
              <RESULTS>
                <RESULT eventid="1076" points="515" reactiontime="+83" swimtime="00:00:25.27" resultid="2951" heatid="7269" lane="9" entrytime="00:00:25.06" />
                <RESULT eventid="1288" points="509" reactiontime="+68" swimtime="00:00:56.27" resultid="2952" heatid="7366" lane="9" entrytime="00:00:56.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="392" reactiontime="+69" swimtime="00:01:08.67" resultid="2953" heatid="7389" lane="9" entrytime="00:01:04.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="486" reactiontime="+67" swimtime="00:00:27.65" resultid="2954" heatid="7449" lane="1" entrytime="00:00:27.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-23" firstname="Katarzyna" gender="F" lastname="Żołnowska" nation="POL" athleteid="2979">
              <RESULTS>
                <RESULT eventid="1059" points="540" swimtime="00:00:28.15" resultid="2980" heatid="7245" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1272" points="579" reactiontime="+77" swimtime="00:01:00.26" resultid="2981" heatid="7348" lane="3" entrytime="00:00:59.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="641" reactiontime="+75" swimtime="00:02:08.07" resultid="2982" heatid="7474" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="637" reactiontime="+80" swimtime="00:04:31.78" resultid="2983" heatid="7566" lane="4" entrytime="00:04:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:04.71" />
                    <SPLIT distance="150" swimtime="00:01:39.13" />
                    <SPLIT distance="200" swimtime="00:02:13.94" />
                    <SPLIT distance="250" swimtime="00:02:48.66" />
                    <SPLIT distance="300" swimtime="00:03:23.61" />
                    <SPLIT distance="350" swimtime="00:03:58.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="590" reactiontime="+65" swimtime="00:01:37.50" resultid="3031" heatid="7496" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                    <SPLIT distance="100" swimtime="00:00:50.31" />
                    <SPLIT distance="150" swimtime="00:01:14.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2950" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3014" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2955" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2992" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kategoria C" eventid="1391" points="493" reactiontime="+91" swimtime="00:01:54.41" resultid="3037" heatid="7406" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:28.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2973" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="3009" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2955" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="3018" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="461" reactiontime="+88" swimtime="00:01:45.83" resultid="3032" heatid="7496" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:00:54.59" />
                    <SPLIT distance="150" swimtime="00:01:20.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2986" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2967" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="3018" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2963" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="464" reactiontime="+83" swimtime="00:01:56.78" resultid="3033" heatid="7406" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                    <SPLIT distance="150" swimtime="00:01:31.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2958" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2963" number="2" reactiontime="+4" />
                    <RELAYPOSITION athleteid="2950" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3014" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1391" status="WDR" swimtime="00:00:00.00" resultid="3038" heatid="7402" lane="3" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2986" number="1" />
                    <RELAYPOSITION athleteid="3014" number="2" />
                    <RELAYPOSITION athleteid="2973" number="3" />
                    <RELAYPOSITION athleteid="2971" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1545" status="WDR" swimtime="00:00:00.00" resultid="3039" heatid="7495" lane="1" entrytime="00:01:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3014" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" />
                    <RELAYPOSITION athleteid="3018" number="3" />
                    <RELAYPOSITION athleteid="2971" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="3030" heatid="7401" lane="5" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3002" number="1" />
                    <RELAYPOSITION athleteid="3023" number="2" />
                    <RELAYPOSITION athleteid="2989" number="3" />
                    <RELAYPOSITION athleteid="2979" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="3035" heatid="7491" lane="5" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3026" number="1" />
                    <RELAYPOSITION athleteid="3023" number="2" />
                    <RELAYPOSITION athleteid="2979" number="3" />
                    <RELAYPOSITION athleteid="2989" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="3034" heatid="7289" lane="6" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2989" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" />
                    <RELAYPOSITION athleteid="3002" number="3" />
                    <RELAYPOSITION athleteid="2992" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="476" reactiontime="+60" swimtime="00:02:03.41" resultid="3036" heatid="7565" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                    <SPLIT distance="100" swimtime="00:01:02.59" />
                    <SPLIT distance="150" swimtime="00:01:29.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2992" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3002" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2967" number="3" reactiontime="+5" />
                    <RELAYPOSITION athleteid="3026" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="622" reactiontime="+66" swimtime="00:01:42.94" resultid="3028" heatid="7289" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                    <SPLIT distance="100" swimtime="00:00:52.39" />
                    <SPLIT distance="150" swimtime="00:01:19.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2955" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3002" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2979" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2992" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" status="WDR" swimtime="00:00:00.00" resultid="3029" heatid="7565" lane="1" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2998" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" />
                    <RELAYPOSITION athleteid="2979" number="3" />
                    <RELAYPOSITION athleteid="3023" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="3040" name="SP Masters Lublin" shortname="Masters Lublin">
          <CONTACT city="LUBLIN" email="masters_lublin@wp.pl" name="WÓJCICKI" phone="+48501794954" state="LUBEL" street="STANISŁAWA LEMA 18" zip="20-445" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-28" firstname="Anna" gender="F" lastname="Michalska" nation="POL" license="103503700002" athleteid="3062">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3071" heatid="7273" lane="6" entrytime="00:03:10.10" />
                <RESULT eventid="1140" points="264" reactiontime="+75" swimtime="00:12:26.41" resultid="3072" heatid="7291" lane="2" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:04.33" />
                    <SPLIT distance="200" swimtime="00:02:50.45" />
                    <SPLIT distance="250" swimtime="00:03:37.21" />
                    <SPLIT distance="300" swimtime="00:04:24.98" />
                    <SPLIT distance="350" swimtime="00:05:13.36" />
                    <SPLIT distance="400" swimtime="00:06:01.77" />
                    <SPLIT distance="450" swimtime="00:06:49.56" />
                    <SPLIT distance="500" swimtime="00:07:37.64" />
                    <SPLIT distance="550" swimtime="00:08:26.46" />
                    <SPLIT distance="600" swimtime="00:09:14.97" />
                    <SPLIT distance="650" swimtime="00:10:02.62" />
                    <SPLIT distance="700" swimtime="00:10:51.44" />
                    <SPLIT distance="750" swimtime="00:11:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="337" reactiontime="+90" swimtime="00:00:36.87" resultid="3073" heatid="7312" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1304" points="310" reactiontime="+93" swimtime="00:01:23.45" resultid="3074" heatid="7372" lane="6" entrytime="00:01:25.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="308" reactiontime="+94" swimtime="00:01:21.45" resultid="3075" heatid="7456" lane="5" entrytime="00:01:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="296" reactiontime="+73" swimtime="00:02:58.77" resultid="3076" heatid="7527" lane="0" entrytime="00:03:02.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:12.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-11" firstname="Mirosław" gender="M" lastname="Molenda" nation="POL" license="103503700012" athleteid="3057">
              <RESULTS>
                <RESULT eventid="1076" points="186" swimtime="00:00:35.45" resultid="3058" heatid="7250" lane="7" entrytime="00:00:39.40" entrycourse="SCM" />
                <RESULT eventid="1288" points="183" swimtime="00:01:19.03" resultid="3059" heatid="7353" lane="1" entrytime="00:01:20.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="179" swimtime="00:02:56.23" resultid="3060" heatid="7478" lane="3" entrytime="00:02:55.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="183" swimtime="00:06:13.70" resultid="3061" heatid="7581" lane="9" entrytime="00:06:35.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="150" swimtime="00:02:13.79" />
                    <SPLIT distance="200" swimtime="00:03:02.82" />
                    <SPLIT distance="250" swimtime="00:03:51.32" />
                    <SPLIT distance="300" swimtime="00:04:40.34" />
                    <SPLIT distance="350" swimtime="00:05:29.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-06" firstname="Marek" gender="M" lastname="Walencik" nation="POL" license="103503700010" athleteid="3052">
              <RESULTS>
                <RESULT eventid="1224" points="318" reactiontime="+79" swimtime="00:00:32.54" resultid="3053" heatid="7323" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1320" points="352" reactiontime="+86" swimtime="00:01:11.18" resultid="3054" heatid="7385" lane="7" entrytime="00:01:12.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="377" reactiontime="+86" swimtime="00:01:16.92" resultid="3055" heatid="7424" lane="1" entrytime="00:01:15.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="3056" heatid="7465" lane="9" entrytime="00:01:14.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-28" firstname="Rafał" gender="M" lastname="Wójcicki" nation="POL" license="103503700001" athleteid="3041">
              <RESULTS>
                <RESULT eventid="1156" points="282" reactiontime="+78" swimtime="00:11:16.09" resultid="3042" heatid="7296" lane="9" entrytime="00:11:30.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                    <SPLIT distance="200" swimtime="00:02:39.20" />
                    <SPLIT distance="250" swimtime="00:03:21.32" />
                    <SPLIT distance="300" swimtime="00:04:03.40" />
                    <SPLIT distance="350" swimtime="00:04:45.79" />
                    <SPLIT distance="400" swimtime="00:05:28.69" />
                    <SPLIT distance="450" swimtime="00:06:11.81" />
                    <SPLIT distance="500" swimtime="00:06:54.61" />
                    <SPLIT distance="550" swimtime="00:07:38.37" />
                    <SPLIT distance="600" swimtime="00:08:22.26" />
                    <SPLIT distance="650" swimtime="00:09:06.31" />
                    <SPLIT distance="700" swimtime="00:09:49.91" />
                    <SPLIT distance="750" swimtime="00:10:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="260" reactiontime="+74" swimtime="00:00:34.80" resultid="3043" heatid="7323" lane="6" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1481" points="265" reactiontime="+74" swimtime="00:01:16.08" resultid="3044" heatid="7464" lane="7" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="294" reactiontime="+80" swimtime="00:00:37.95" resultid="3045" heatid="7554" lane="0" entrytime="00:00:38.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-28" firstname="Łukasz" gender="M" lastname="Wójcicki" nation="POL" license="103503700004" athleteid="3049">
              <RESULTS>
                <RESULT eventid="1417" points="187" reactiontime="+82" swimtime="00:01:37.11" resultid="3050" heatid="7417" lane="5" entrytime="00:01:41.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="200" reactiontime="+73" swimtime="00:00:43.12" resultid="3051" heatid="7548" lane="4" entrytime="00:00:48.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-07" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" license="103503700005" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1288" points="305" reactiontime="+97" swimtime="00:01:06.74" resultid="3047" heatid="7357" lane="0" entrytime="00:01:08.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3048" heatid="7480" lane="4" entrytime="00:02:35.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="277" reactiontime="+78" swimtime="00:02:18.65" resultid="3069" heatid="7404" lane="4" entrytime="00:02:12.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3052" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3049" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3041" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3046" number="4" reactiontime="+84" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="299" reactiontime="+89" swimtime="00:02:02.26" resultid="3070" heatid="7494" lane="2" entrytime="00:01:55.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:33.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3052" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3057" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3041" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3046" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SPKAR" nation="POL" region="14" clubid="4412" name="SP Sebastiana Karasia W-wa">
          <CONTACT city="Łomianki" email="karas.sebastian@o2.pl" name="Karaś" phone="509425753" street="Irysa 23" zip="05-092" />
          <ATHLETES>
            <ATHLETE birthdate="1989-06-30" firstname="Alan" gender="M" lastname="Bistron" nation="POL" athleteid="4436">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4437" heatid="7333" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1352" points="101" reactiontime="+95" swimtime="00:03:51.68" resultid="4438" heatid="7395" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="4439" heatid="7461" lane="3" entrytime="00:01:45.00" />
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="4440" heatid="8155" lane="3" entrytime="00:07:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-09-20" firstname="Ewa" gender="F" lastname="Borys" nation="POL" athleteid="4431">
              <RESULTS>
                <RESULT eventid="1092" points="207" reactiontime="+85" swimtime="00:03:25.95" resultid="4432" heatid="7271" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                    <SPLIT distance="150" swimtime="00:02:39.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="210" reactiontime="+77" swimtime="00:00:43.17" resultid="4433" heatid="7309" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1304" points="208" reactiontime="+86" swimtime="00:01:35.35" resultid="4434" heatid="7370" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="190" reactiontime="+79" swimtime="00:01:35.58" resultid="4435" heatid="7454" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="4420">
              <RESULTS>
                <RESULT eventid="1076" points="464" reactiontime="+87" swimtime="00:00:26.16" resultid="4421" heatid="7267" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1288" points="475" reactiontime="+85" swimtime="00:00:57.57" resultid="4422" heatid="7363" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="447" reactiontime="+77" swimtime="00:02:09.88" resultid="4423" heatid="7485" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="150" swimtime="00:01:37.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-12" firstname="Tobiasz" gender="M" lastname="Jankowski" nation="POL" athleteid="4451">
              <RESULTS>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="4452" heatid="7379" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1417" points="249" reactiontime="+91" swimtime="00:01:28.38" resultid="4453" heatid="7416" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-03-06" firstname="Aleksandra" gender="F" lastname="Jurczak" nation="POL" athleteid="4444">
              <RESULTS>
                <RESULT eventid="1272" points="199" reactiontime="+99" swimtime="00:01:26.00" resultid="4445" heatid="7343" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="171" swimtime="00:01:41.79" resultid="4446" heatid="7369" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="178" reactiontime="+57" swimtime="00:01:50.82" resultid="4447" heatid="7409" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="167" swimtime="00:03:20.27" resultid="4448" heatid="7470" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:34.63" />
                    <SPLIT distance="150" swimtime="00:02:28.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-07-07" firstname="Piotr" gender="M" lastname="Karczewski" nation="POL" athleteid="4424">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4425" heatid="7253" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1288" points="168" swimtime="00:01:21.44" resultid="4426" heatid="7353" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="4427" heatid="7378" lane="4" entrytime="00:01:45.00" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="4428" heatid="7417" lane="0" entrytime="00:01:50.00" />
                <RESULT eventid="1513" points="178" swimtime="00:02:56.35" resultid="4429" heatid="7478" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:25.20" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4430" heatid="7549" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-08" firstname="Natalia" gender="F" lastname="Konwerska" nation="POL" athleteid="4413">
              <RESULTS>
                <RESULT eventid="1433" points="505" reactiontime="+69" swimtime="00:00:30.60" resultid="4414" heatid="7433" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-29" firstname="Aleksandra" gender="F" lastname="Rudzka" nation="POL" athleteid="4449">
              <RESULTS>
                <RESULT eventid="1465" status="WDR" swimtime="00:00:00.00" resultid="4450" heatid="7457" lane="0" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-10-29" firstname="Dorota" gender="F" lastname="Zembrzuska" nation="POL" athleteid="4441">
              <RESULTS>
                <RESULT eventid="1272" points="395" reactiontime="+99" swimtime="00:01:08.45" resultid="4442" heatid="7346" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4443" heatid="7473" lane="7" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-26" firstname="Radosław" gender="M" lastname="Łopiński" nation="POL" athleteid="8163" />
            <ATHLETE birthdate="1980-01-02" firstname="Ewa" gender="F" lastname="Łukasiuk" nation="POL" athleteid="4415">
              <RESULTS>
                <RESULT eventid="1059" points="391" reactiontime="+75" swimtime="00:00:31.35" resultid="4416" heatid="7242" lane="2" entrytime="00:00:31.90" />
                <RESULT eventid="1272" points="327" reactiontime="+76" swimtime="00:01:12.92" resultid="4417" heatid="7345" lane="0" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="309" reactiontime="+72" swimtime="00:01:32.23" resultid="4418" heatid="7412" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="348" reactiontime="+66" swimtime="00:00:40.58" resultid="4419" heatid="7542" lane="4" entrytime="00:00:41.91" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="290" reactiontime="+78" swimtime="00:02:03.58" resultid="4458" heatid="7492" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:00:56.76" />
                    <SPLIT distance="150" swimtime="00:01:28.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4451" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4420" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="8163" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="4424" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Karaś Team" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="200" reactiontime="+47" swimtime="00:02:34.53" resultid="4456" heatid="7405" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                    <SPLIT distance="150" swimtime="00:02:08.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4424" number="1" reactiontime="+47" status="DSQ" />
                    <RELAYPOSITION athleteid="4451" number="2" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="4436" number="3" reactiontime="-8" status="DSQ" />
                    <RELAYPOSITION athleteid="4420" number="4" reactiontime="+35" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="Karaś Team" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="428" reactiontime="+64" swimtime="00:02:15.84" resultid="4455" heatid="7400" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:45.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4449" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4415" number="2" reactiontime="+10" />
                    <RELAYPOSITION athleteid="4413" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="4441" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Karaś Team" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="317" reactiontime="+70" swimtime="00:02:17.70" resultid="4457" heatid="7489" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="150" swimtime="00:01:45.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4415" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4431" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4444" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4441" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Karaś Team" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="290" reactiontime="+76" swimtime="00:02:12.64" resultid="4454" heatid="7286" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:00:57.74" />
                    <SPLIT distance="150" swimtime="00:01:34.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4415" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4420" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4431" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4424" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02415" nation="POL" region="15" clubid="5573" name="Start Poznań">
          <CONTACT city="Dopiewiec" email="kaczy4@autograf.pl" name="Kaczmarek" phone="603434586" street="Promenada 21" zip="62-070" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-16" firstname="Aneta" gender="F" lastname="Andrzejewska" nation="POL" athleteid="5608">
              <RESULTS>
                <RESULT eventid="1059" points="217" reactiontime="+94" swimtime="00:00:38.12" resultid="5609" heatid="7238" lane="2" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1240" points="234" swimtime="00:03:38.23" resultid="5610" heatid="7329" lane="8" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:44.86" />
                    <SPLIT distance="150" swimtime="00:02:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="162" reactiontime="+98" swimtime="00:01:32.06" resultid="5611" heatid="7341" lane="4" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="224" swimtime="00:01:42.53" resultid="5612" heatid="7410" lane="9" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="189" swimtime="00:03:12.28" resultid="5613" heatid="7469" lane="2" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:31.84" />
                    <SPLIT distance="150" swimtime="00:02:21.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="228" reactiontime="+97" swimtime="00:00:46.69" resultid="5614" heatid="7540" lane="2" entrytime="00:00:47.00" entrycourse="SCM" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5615" heatid="7570" lane="7" entrytime="00:07:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-16" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="5616">
              <RESULTS>
                <RESULT eventid="1076" points="451" reactiontime="+90" swimtime="00:00:26.40" resultid="5617" heatid="7264" lane="8" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5618" heatid="7283" lane="9" entrytime="00:02:35.00" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5619" heatid="7364" lane="9" entrytime="00:00:59.00" entrycourse="SCM" />
                <RESULT eventid="1320" points="470" reactiontime="+73" swimtime="00:01:04.61" resultid="5620" heatid="7387" lane="6" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="450" reactiontime="+72" swimtime="00:00:28.38" resultid="5621" heatid="7446" lane="2" entrytime="00:00:29.50" entrycourse="SCM" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="5622" heatid="7466" lane="9" entrytime="00:01:08.00" entrycourse="SCM" />
                <RESULT eventid="1625" points="431" reactiontime="+79" swimtime="00:01:03.63" resultid="5623" heatid="7519" lane="2" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5624" heatid="7535" lane="0" entrytime="00:02:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-09-10" firstname="Sylwia" gender="F" lastname="Czapla" nation="POL" athleteid="5640">
              <RESULTS>
                <RESULT eventid="1059" points="158" reactiontime="+88" swimtime="00:00:42.38" resultid="5641" heatid="7236" lane="3" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1272" points="131" swimtime="00:01:38.81" resultid="5642" heatid="7340" lane="4" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="103" reactiontime="+86" swimtime="00:00:51.88" resultid="5643" heatid="7427" lane="2" entrytime="00:00:52.00" entrycourse="SCM" />
                <RESULT eventid="1673" points="152" reactiontime="+94" swimtime="00:00:53.47" resultid="5644" heatid="7539" lane="9" entrytime="00:00:54.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-01" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="5650">
              <RESULTS>
                <RESULT eventid="1256" points="291" reactiontime="+90" swimtime="00:03:01.18" resultid="5651" heatid="7336" lane="4" entrytime="00:03:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="344" reactiontime="+86" swimtime="00:01:19.33" resultid="5652" heatid="7420" lane="5" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="352" reactiontime="+76" swimtime="00:00:35.74" resultid="5653" heatid="7553" lane="3" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-03" firstname="Michał" gender="M" lastname="Kaczmarek" nation="POL" athleteid="5583">
              <RESULTS>
                <RESULT eventid="1076" points="341" reactiontime="+98" swimtime="00:00:28.98" resultid="5584" heatid="7259" lane="1" entrytime="00:00:29.14" entrycourse="SCM" />
                <RESULT eventid="1108" points="255" swimtime="00:02:52.72" resultid="5585" heatid="7280" lane="5" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="284" swimtime="00:03:02.76" resultid="5586" heatid="7337" lane="8" entrytime="00:03:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                    <SPLIT distance="150" swimtime="00:02:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="295" swimtime="00:01:15.46" resultid="5587" heatid="7382" lane="8" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="300" reactiontime="+72" swimtime="00:01:23.01" resultid="5588" heatid="7421" lane="8" entrytime="00:01:22.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="233" swimtime="00:06:22.59" resultid="5589" heatid="8156" lane="2" entrytime="00:06:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:31.72" />
                    <SPLIT distance="150" swimtime="00:02:23.99" />
                    <SPLIT distance="200" swimtime="00:03:13.51" />
                    <SPLIT distance="250" swimtime="00:04:05.16" />
                    <SPLIT distance="300" swimtime="00:04:55.84" />
                    <SPLIT distance="350" swimtime="00:05:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="5590" heatid="7515" lane="5" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5591" heatid="7554" lane="5" entrytime="00:00:37.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-16" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="5592">
              <RESULTS>
                <RESULT eventid="1108" points="278" reactiontime="+82" swimtime="00:02:47.88" resultid="5593" heatid="7281" lane="7" entrytime="00:02:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                    <SPLIT distance="150" swimtime="00:02:09.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="288" reactiontime="+82" swimtime="00:03:01.75" resultid="5594" heatid="7337" lane="6" entrytime="00:02:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:26.57" />
                    <SPLIT distance="150" swimtime="00:02:13.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="191" reactiontime="+86" swimtime="00:03:07.64" resultid="5595" heatid="7397" lane="9" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:14.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="280" reactiontime="+81" swimtime="00:01:25.00" resultid="5596" heatid="7421" lane="2" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="266" reactiontime="+88" swimtime="00:06:05.86" resultid="5597" heatid="8157" lane="8" entrytime="00:05:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:12.21" />
                    <SPLIT distance="200" swimtime="00:02:58.01" />
                    <SPLIT distance="250" swimtime="00:03:50.48" />
                    <SPLIT distance="300" swimtime="00:04:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="191" reactiontime="+87" swimtime="00:01:23.41" resultid="5598" heatid="7520" lane="5" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-03" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="5574">
              <RESULTS>
                <RESULT eventid="1059" points="392" swimtime="00:00:31.31" resultid="5575" heatid="7242" lane="3" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1140" points="371" reactiontime="+89" swimtime="00:11:06.68" resultid="5576" heatid="7290" lane="9" entrytime="00:12:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:58.05" />
                    <SPLIT distance="200" swimtime="00:02:39.63" />
                    <SPLIT distance="250" swimtime="00:03:21.73" />
                    <SPLIT distance="300" swimtime="00:04:04.00" />
                    <SPLIT distance="350" swimtime="00:04:46.60" />
                    <SPLIT distance="400" swimtime="00:05:29.52" />
                    <SPLIT distance="450" swimtime="00:06:12.66" />
                    <SPLIT distance="500" swimtime="00:06:55.44" />
                    <SPLIT distance="550" swimtime="00:07:38.67" />
                    <SPLIT distance="600" swimtime="00:08:21.61" />
                    <SPLIT distance="650" swimtime="00:09:04.17" />
                    <SPLIT distance="700" swimtime="00:09:46.03" />
                    <SPLIT distance="750" swimtime="00:10:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="392" reactiontime="+76" swimtime="00:00:35.07" resultid="5577" heatid="7313" lane="8" entrytime="00:00:34.50" entrycourse="SCM" />
                <RESULT eventid="1272" points="412" reactiontime="+86" swimtime="00:01:07.48" resultid="5578" heatid="7346" lane="5" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="382" reactiontime="+79" swimtime="00:01:15.82" resultid="5579" heatid="7455" lane="9" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="401" reactiontime="+87" swimtime="00:02:29.63" resultid="5580" heatid="7473" lane="8" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="411" reactiontime="+79" swimtime="00:02:40.26" resultid="5581" heatid="7528" lane="0" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:01:59.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="386" reactiontime="+83" swimtime="00:05:21.17" resultid="5582" heatid="7569" lane="4" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:55.42" />
                    <SPLIT distance="200" swimtime="00:02:36.72" />
                    <SPLIT distance="250" swimtime="00:03:18.12" />
                    <SPLIT distance="300" swimtime="00:03:59.41" />
                    <SPLIT distance="350" swimtime="00:04:40.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-09" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="5599">
              <RESULTS>
                <RESULT eventid="1059" points="337" reactiontime="+93" swimtime="00:00:32.94" resultid="5600" heatid="7240" lane="1" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1140" points="278" reactiontime="+98" swimtime="00:12:13.80" resultid="5601" heatid="7291" lane="8" entrytime="00:12:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:09.77" />
                    <SPLIT distance="200" swimtime="00:02:55.40" />
                    <SPLIT distance="250" swimtime="00:03:41.41" />
                    <SPLIT distance="300" swimtime="00:04:27.29" />
                    <SPLIT distance="350" swimtime="00:05:13.72" />
                    <SPLIT distance="400" swimtime="00:06:00.08" />
                    <SPLIT distance="450" swimtime="00:06:46.72" />
                    <SPLIT distance="500" swimtime="00:07:34.10" />
                    <SPLIT distance="550" swimtime="00:08:21.30" />
                    <SPLIT distance="600" swimtime="00:09:08.97" />
                    <SPLIT distance="650" swimtime="00:09:56.38" />
                    <SPLIT distance="700" swimtime="00:10:43.51" />
                    <SPLIT distance="750" swimtime="00:11:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="314" reactiontime="+94" swimtime="00:01:13.88" resultid="5602" heatid="7345" lane="9" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="246" reactiontime="+94" swimtime="00:03:10.67" resultid="5603" heatid="7392" lane="4" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                    <SPLIT distance="100" swimtime="00:01:31.55" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="315" reactiontime="+91" swimtime="00:00:35.80" resultid="5604" heatid="7431" lane="6" entrytime="00:00:35.30" entrycourse="SCM" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="5605" heatid="7471" lane="7" entrytime="00:02:55.00" entrycourse="SCM" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="5606" heatid="7509" lane="4" entrytime="00:01:26.00" entrycourse="SCM" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5607" heatid="7568" lane="9" entrytime="00:06:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-02" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="5634">
              <RESULTS>
                <RESULT eventid="1076" points="407" reactiontime="+84" swimtime="00:00:27.32" resultid="5635" heatid="7265" lane="3" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="391" reactiontime="+84" swimtime="00:02:29.84" resultid="5636" heatid="7283" lane="7" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:10.67" />
                    <SPLIT distance="150" swimtime="00:01:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="441" reactiontime="+87" swimtime="00:00:59.00" resultid="5637" heatid="7365" lane="0" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="453" reactiontime="+75" swimtime="00:02:09.36" resultid="5638" heatid="7486" lane="7" entrytime="00:02:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="150" swimtime="00:01:35.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="415" reactiontime="+82" swimtime="00:04:44.33" resultid="5639" heatid="7574" lane="5" entrytime="00:04:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:43.18" />
                    <SPLIT distance="200" swimtime="00:02:20.40" />
                    <SPLIT distance="250" swimtime="00:02:56.07" />
                    <SPLIT distance="300" swimtime="00:03:32.51" />
                    <SPLIT distance="350" swimtime="00:04:08.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-08" firstname="Sławomir" gender="M" lastname="Parysek" nation="POL" athleteid="5625">
              <RESULTS>
                <RESULT eventid="1076" points="320" reactiontime="+79" swimtime="00:00:29.60" resultid="5626" heatid="7257" lane="3" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="278" reactiontime="+78" swimtime="00:02:47.82" resultid="5627" heatid="7281" lane="6" entrytime="00:02:46.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                    <SPLIT distance="150" swimtime="00:02:10.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="320" reactiontime="+72" swimtime="00:01:13.41" resultid="5628" heatid="7384" lane="2" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="176" reactiontime="+89" swimtime="00:03:12.93" resultid="5629" heatid="7396" lane="3" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="150" swimtime="00:02:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="309" reactiontime="+77" swimtime="00:00:32.14" resultid="5630" heatid="7442" lane="0" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1577" points="245" reactiontime="+76" swimtime="00:06:16.02" resultid="5631" heatid="8157" lane="9" entrytime="00:06:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                    <SPLIT distance="200" swimtime="00:03:01.99" />
                    <SPLIT distance="250" swimtime="00:03:57.37" />
                    <SPLIT distance="300" swimtime="00:04:53.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="242" reactiontime="+70" swimtime="00:01:17.09" resultid="5632" heatid="7516" lane="6" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="281" reactiontime="+71" swimtime="00:00:38.52" resultid="5633" heatid="7553" lane="5" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-06-03" firstname="Anna" gender="F" lastname="Rostkowska-Kaczmarek" nation="POL" athleteid="5645">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="5646" heatid="7241" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="5647" heatid="7344" lane="1" entrytime="00:01:17.00" />
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="5648" heatid="7410" lane="8" entrytime="00:01:45.00" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5649" heatid="7539" lane="4" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="341" reactiontime="+53" swimtime="00:02:09.38" resultid="5656" heatid="7403" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                    <SPLIT distance="150" swimtime="00:01:41.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5616" number="1" reactiontime="+53" />
                    <RELAYPOSITION athleteid="5650" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5592" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="5634" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" status="DNS" swimtime="00:00:00.00" resultid="5658" heatid="7492" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5625" number="1" />
                    <RELAYPOSITION athleteid="5583" number="2" />
                    <RELAYPOSITION athleteid="5592" number="3" />
                    <RELAYPOSITION athleteid="5634" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="5655" heatid="7400" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5574" number="1" />
                    <RELAYPOSITION athleteid="5608" number="2" />
                    <RELAYPOSITION athleteid="5599" number="3" />
                    <RELAYPOSITION athleteid="5645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="5657" heatid="7489" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5608" number="1" />
                    <RELAYPOSITION athleteid="5574" number="2" />
                    <RELAYPOSITION athleteid="5599" number="3" />
                    <RELAYPOSITION athleteid="5645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="5654" heatid="7287" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5625" number="1" />
                    <RELAYPOSITION athleteid="5583" number="2" />
                    <RELAYPOSITION athleteid="5599" number="3" />
                    <RELAYPOSITION athleteid="5645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="305" reactiontime="+78" swimtime="00:02:23.11" resultid="5659" heatid="7562" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:10.96" />
                    <SPLIT distance="150" swimtime="00:01:44.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5574" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5650" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5625" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="5608" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STBYD" nation="POL" region="02" clubid="2384" name="Stashky Team Bydgoszcz">
          <ATHLETES>
            <ATHLETE birthdate="1968-04-21" firstname="Radosław" gender="M" lastname="Staszkiewicz" nation="POL" athleteid="2383">
              <RESULTS>
                <RESULT eventid="1108" points="272" swimtime="00:02:49.06" resultid="2385" heatid="7282" lane="9" entrytime="00:02:43.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:02:09.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="281" swimtime="00:21:33.78" resultid="2386" heatid="7303" lane="3" entrytime="00:21:27.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:02.53" />
                    <SPLIT distance="200" swimtime="00:02:46.01" />
                    <SPLIT distance="250" swimtime="00:03:30.01" />
                    <SPLIT distance="300" swimtime="00:04:13.88" />
                    <SPLIT distance="350" swimtime="00:04:57.75" />
                    <SPLIT distance="400" swimtime="00:05:41.60" />
                    <SPLIT distance="450" swimtime="00:06:24.83" />
                    <SPLIT distance="500" swimtime="00:07:08.20" />
                    <SPLIT distance="550" swimtime="00:07:52.31" />
                    <SPLIT distance="600" swimtime="00:08:35.63" />
                    <SPLIT distance="650" swimtime="00:09:19.25" />
                    <SPLIT distance="700" swimtime="00:10:02.86" />
                    <SPLIT distance="750" swimtime="00:10:46.44" />
                    <SPLIT distance="800" swimtime="00:11:30.00" />
                    <SPLIT distance="850" swimtime="00:12:13.31" />
                    <SPLIT distance="900" swimtime="00:12:57.02" />
                    <SPLIT distance="950" swimtime="00:13:40.86" />
                    <SPLIT distance="1000" swimtime="00:14:23.95" />
                    <SPLIT distance="1050" swimtime="00:15:06.99" />
                    <SPLIT distance="1100" swimtime="00:15:50.23" />
                    <SPLIT distance="1150" swimtime="00:16:33.05" />
                    <SPLIT distance="1200" swimtime="00:17:16.31" />
                    <SPLIT distance="1250" swimtime="00:18:00.05" />
                    <SPLIT distance="1300" swimtime="00:18:43.50" />
                    <SPLIT distance="1350" swimtime="00:19:26.43" />
                    <SPLIT distance="1400" swimtime="00:20:10.27" />
                    <SPLIT distance="1450" swimtime="00:20:53.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="276" reactiontime="+86" swimtime="00:01:17.14" resultid="2388" heatid="7384" lane="6" entrytime="00:01:13.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="277" swimtime="00:02:45.99" resultid="2389" heatid="7397" lane="7" entrytime="00:02:46.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:02:00.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="317" swimtime="00:00:31.89" resultid="2390" heatid="7443" lane="6" entrytime="00:00:31.41" />
                <RESULT eventid="1577" points="276" swimtime="00:06:01.43" resultid="2391" heatid="8157" lane="1" entrytime="00:05:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:02:04.38" />
                    <SPLIT distance="200" swimtime="00:02:51.96" />
                    <SPLIT distance="250" swimtime="00:03:45.38" />
                    <SPLIT distance="300" swimtime="00:04:38.99" />
                    <SPLIT distance="350" swimtime="00:05:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="316" swimtime="00:01:10.56" resultid="2392" heatid="7518" lane="2" entrytime="00:01:10.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="283" swimtime="00:05:23.20" resultid="2393" heatid="7577" lane="0" entrytime="00:05:19.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                    <SPLIT distance="200" swimtime="00:02:36.13" />
                    <SPLIT distance="250" swimtime="00:03:18.52" />
                    <SPLIT distance="300" swimtime="00:04:01.14" />
                    <SPLIT distance="350" swimtime="00:04:43.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" nation="POL" region="01" clubid="3442" name="Steef Wrocław">
          <CONTACT city="Wrocław" email="stee1@wp.pl" name="Stefan Skrzypek" street="Edyty Stein 6m1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="3443">
              <RESULTS>
                <RESULT eventid="1092" points="282" swimtime="00:03:05.70" resultid="3444" heatid="7273" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="269" reactiontime="+99" swimtime="00:23:43.73" resultid="3445" heatid="7300" lane="1" entrytime="00:23:52.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="150" swimtime="00:02:14.45" />
                    <SPLIT distance="200" swimtime="00:03:01.33" />
                    <SPLIT distance="250" swimtime="00:03:48.08" />
                    <SPLIT distance="300" swimtime="00:04:35.29" />
                    <SPLIT distance="350" swimtime="00:05:21.07" />
                    <SPLIT distance="400" swimtime="00:06:07.21" />
                    <SPLIT distance="450" swimtime="00:06:54.40" />
                    <SPLIT distance="500" swimtime="00:07:41.52" />
                    <SPLIT distance="550" swimtime="00:08:28.82" />
                    <SPLIT distance="600" swimtime="00:09:17.24" />
                    <SPLIT distance="650" swimtime="00:10:04.83" />
                    <SPLIT distance="700" swimtime="00:10:53.17" />
                    <SPLIT distance="750" swimtime="00:11:42.05" />
                    <SPLIT distance="800" swimtime="00:12:30.07" />
                    <SPLIT distance="850" swimtime="00:13:18.87" />
                    <SPLIT distance="900" swimtime="00:14:07.61" />
                    <SPLIT distance="950" swimtime="00:14:56.04" />
                    <SPLIT distance="1000" swimtime="00:15:44.49" />
                    <SPLIT distance="1050" swimtime="00:16:32.92" />
                    <SPLIT distance="1100" swimtime="00:17:20.60" />
                    <SPLIT distance="1150" swimtime="00:18:08.49" />
                    <SPLIT distance="1200" swimtime="00:18:56.47" />
                    <SPLIT distance="1250" swimtime="00:19:44.30" />
                    <SPLIT distance="1300" swimtime="00:20:32.11" />
                    <SPLIT distance="1350" swimtime="00:21:19.91" />
                    <SPLIT distance="1400" swimtime="00:22:08.00" />
                    <SPLIT distance="1450" swimtime="00:22:56.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="265" reactiontime="+95" swimtime="00:01:27.93" resultid="3446" heatid="7372" lane="7" entrytime="00:01:28.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="241" reactiontime="+88" swimtime="00:01:28.41" resultid="3447" heatid="7455" lane="3" entrytime="00:01:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="276" reactiontime="+99" swimtime="00:06:37.47" resultid="3448" heatid="8150" lane="5" entrytime="00:06:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:37.13" />
                    <SPLIT distance="150" swimtime="00:02:26.94" />
                    <SPLIT distance="200" swimtime="00:03:15.58" />
                    <SPLIT distance="250" swimtime="00:04:12.06" />
                    <SPLIT distance="300" swimtime="00:05:08.42" />
                    <SPLIT distance="350" swimtime="00:05:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="260" reactiontime="+83" swimtime="00:03:06.66" resultid="3449" heatid="7526" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="263" reactiontime="+84" swimtime="00:06:04.86" resultid="3450" heatid="7569" lane="6" entrytime="00:06:02.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:13.52" />
                    <SPLIT distance="200" swimtime="00:03:00.45" />
                    <SPLIT distance="250" swimtime="00:03:47.48" />
                    <SPLIT distance="300" swimtime="00:04:33.80" />
                    <SPLIT distance="350" swimtime="00:05:20.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCMWR" nation="POL" region="01" clubid="6327" name="Swim Club Masters Wrocław">
          <CONTACT city="wrocław" email="stasiaczekmichal@gmail.com" name="Stasiaczek Michał" phone="792883772" street="Dożynkowa 15/7" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="6328">
              <RESULTS>
                <RESULT eventid="1240" points="233" reactiontime="+82" swimtime="00:03:38.62" resultid="6329" heatid="7329" lane="1" entrytime="00:03:48.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                    <SPLIT distance="100" swimtime="00:01:45.31" />
                    <SPLIT distance="150" swimtime="00:02:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="189" reactiontime="+66" swimtime="00:01:38.31" resultid="6330" heatid="7370" lane="2" entrytime="00:01:40.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="234" reactiontime="+69" swimtime="00:01:41.16" resultid="6331" heatid="7410" lane="2" entrytime="00:01:44.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="120" reactiontime="+83" swimtime="00:00:49.32" resultid="6332" heatid="7427" lane="4" entrytime="00:00:49.72" />
                <RESULT eventid="1673" points="262" reactiontime="+70" swimtime="00:00:44.63" resultid="6333" heatid="7540" lane="7" entrytime="00:00:47.02" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWIIR" nation="IRL" clubid="2007" name="Swim Ireland">
          <CONTACT city="Dublin" email="jkk@fusbro.com" name="Kruszyna - Kotulski Jerzy" phone="353879305286" />
          <ATHLETES>
            <ATHLETE birthdate="1979-05-25" firstname="Jerzy" gender="M" lastname="Kruszyna - Kotulski" nation="IRL" license="30019411" athleteid="2008">
              <RESULTS>
                <RESULT eventid="1288" points="385" reactiontime="+80" swimtime="00:01:01.76" resultid="2009" heatid="7360" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="383" reactiontime="+78" swimtime="00:00:29.93" resultid="2011" heatid="7446" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1625" points="358" reactiontime="+79" swimtime="00:01:07.71" resultid="2012" heatid="7519" lane="9" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="322" reactiontime="+63" swimtime="00:00:36.83" resultid="2013" heatid="7555" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1320" points="326" reactiontime="+74" swimtime="00:01:12.97" resultid="2014" heatid="7385" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STRZE" nation="POL" region="08" clubid="5711" name="Swim Tri Rzeszów">
          <CONTACT city="RZESZÓW" email="KLUB@SWIMTRI.PL" name="SWIM TRI RZESZÓW" street="POPIEŁUSZKI  26 C" zip="35-328" />
          <ATHLETES>
            <ATHLETE birthdate="1974-12-10" firstname="Nikodem" gender="M" lastname="Bernacki" nation="POL" athleteid="5720">
              <RESULTS>
                <RESULT eventid="1076" points="247" swimtime="00:00:32.26" resultid="5721" heatid="7253" lane="0" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1156" points="227" reactiontime="+98" swimtime="00:12:06.06" resultid="5722" heatid="7295" lane="6" entrytime="00:10:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:02.36" />
                    <SPLIT distance="200" swimtime="00:02:47.45" />
                    <SPLIT distance="250" swimtime="00:03:33.51" />
                    <SPLIT distance="300" swimtime="00:04:20.46" />
                    <SPLIT distance="350" swimtime="00:05:06.59" />
                    <SPLIT distance="400" swimtime="00:05:53.17" />
                    <SPLIT distance="450" swimtime="00:06:40.56" />
                    <SPLIT distance="500" swimtime="00:07:27.05" />
                    <SPLIT distance="550" swimtime="00:08:14.14" />
                    <SPLIT distance="600" swimtime="00:09:00.94" />
                    <SPLIT distance="650" swimtime="00:09:48.26" />
                    <SPLIT distance="700" swimtime="00:10:35.76" />
                    <SPLIT distance="750" swimtime="00:11:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="235" swimtime="00:01:12.75" resultid="5723" heatid="7354" lane="7" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="218" swimtime="00:02:45.04" resultid="5724" heatid="7480" lane="6" entrytime="00:02:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:02:02.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5725" heatid="7577" lane="3" entrytime="00:05:12.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-04" firstname="Agata" gender="F" lastname="Borcz-Jajuga" nation="POL" athleteid="5734">
              <RESULTS>
                <RESULT eventid="1059" points="197" reactiontime="+92" swimtime="00:00:39.36" resultid="5735" heatid="7236" lane="5" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1207" points="197" reactiontime="+90" swimtime="00:00:44.07" resultid="5736" heatid="7309" lane="0" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1304" points="192" reactiontime="+84" swimtime="00:01:37.86" resultid="5737" heatid="7370" lane="4" entrytime="00:01:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="179" reactiontime="+94" swimtime="00:00:43.23" resultid="5738" heatid="7427" lane="8" entrytime="00:00:55.00" entrycourse="SCM" />
                <RESULT eventid="1497" points="153" reactiontime="+95" swimtime="00:03:26.35" resultid="5739" heatid="7470" lane="3" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:33.19" />
                    <SPLIT distance="150" swimtime="00:02:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5740" heatid="7569" lane="3" entrytime="00:06:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="6497">
              <RESULTS>
                <RESULT eventid="1076" points="254" reactiontime="+88" swimtime="00:00:31.98" resultid="6499" heatid="7255" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1188" points="195" reactiontime="+85" swimtime="00:24:20.45" resultid="6500" heatid="7304" lane="6" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="150" swimtime="00:02:10.18" />
                    <SPLIT distance="200" swimtime="00:02:57.48" />
                    <SPLIT distance="250" swimtime="00:03:45.55" />
                    <SPLIT distance="350" swimtime="00:05:22.35" />
                    <SPLIT distance="400" swimtime="00:06:10.57" />
                    <SPLIT distance="450" swimtime="00:06:58.72" />
                    <SPLIT distance="500" swimtime="00:07:46.92" />
                    <SPLIT distance="550" swimtime="00:08:35.78" />
                    <SPLIT distance="600" swimtime="00:09:24.60" />
                    <SPLIT distance="650" swimtime="00:10:13.59" />
                    <SPLIT distance="700" swimtime="00:11:02.26" />
                    <SPLIT distance="750" swimtime="00:11:51.49" />
                    <SPLIT distance="800" swimtime="00:12:40.99" />
                    <SPLIT distance="850" swimtime="00:13:30.42" />
                    <SPLIT distance="900" swimtime="00:14:20.71" />
                    <SPLIT distance="950" swimtime="00:15:09.96" />
                    <SPLIT distance="1000" swimtime="00:16:01.27" />
                    <SPLIT distance="1100" swimtime="00:17:43.07" />
                    <SPLIT distance="1150" swimtime="00:18:32.69" />
                    <SPLIT distance="1200" swimtime="00:19:24.56" />
                    <SPLIT distance="1250" swimtime="00:20:14.38" />
                    <SPLIT distance="1300" swimtime="00:21:05.49" />
                    <SPLIT distance="1350" swimtime="00:21:56.45" />
                    <SPLIT distance="1400" swimtime="00:22:46.20" />
                    <SPLIT distance="1450" swimtime="00:23:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="246" reactiontime="+69" swimtime="00:01:11.71" resultid="6501" heatid="7355" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="6502" heatid="7380" lane="9" entrytime="00:01:33.00" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6503" heatid="7438" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1513" points="213" reactiontime="+85" swimtime="00:02:46.26" resultid="6504" heatid="7478" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="197" reactiontime="+90" swimtime="00:06:04.30" resultid="6505" heatid="7581" lane="4" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                    <SPLIT distance="150" swimtime="00:02:10.57" />
                    <SPLIT distance="200" swimtime="00:02:56.40" />
                    <SPLIT distance="250" swimtime="00:03:42.18" />
                    <SPLIT distance="300" swimtime="00:04:29.38" />
                    <SPLIT distance="350" swimtime="00:05:15.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-11-15" firstname="Mariusz" gender="M" lastname="Faff" nation="POL" athleteid="5726">
              <RESULTS>
                <RESULT eventid="1076" points="347" swimtime="00:00:28.83" resultid="5727" heatid="7261" lane="0" entrytime="00:00:28.24" entrycourse="SCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5728" heatid="7283" lane="6" entrytime="00:02:28.64" entrycourse="SCM" />
                <RESULT eventid="1224" points="247" reactiontime="+96" swimtime="00:00:35.38" resultid="5729" heatid="7321" lane="4" entrytime="00:00:35.89" entrycourse="SCM" />
                <RESULT eventid="1288" points="343" reactiontime="+87" swimtime="00:01:04.19" resultid="5730" heatid="7359" lane="5" entrytime="00:01:04.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="314" reactiontime="+85" swimtime="00:00:31.98" resultid="5731" heatid="7443" lane="1" entrytime="00:00:31.60" entrycourse="SCM" />
                <RESULT eventid="1513" points="314" reactiontime="+84" swimtime="00:02:26.13" resultid="5732" heatid="7482" lane="7" entrytime="00:02:28.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="150" swimtime="00:01:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="314" reactiontime="+85" swimtime="00:05:12.11" resultid="5733" heatid="7576" lane="1" entrytime="00:05:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                    <SPLIT distance="200" swimtime="00:02:30.98" />
                    <SPLIT distance="250" swimtime="00:03:11.46" />
                    <SPLIT distance="300" swimtime="00:03:51.98" />
                    <SPLIT distance="350" swimtime="00:04:32.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-10-31" firstname="Tomasz" gender="M" lastname="Sarna" nation="POL" athleteid="5712">
              <RESULTS>
                <RESULT eventid="1076" points="405" reactiontime="+87" swimtime="00:00:27.37" resultid="5713" heatid="7263" lane="6" entrytime="00:00:27.28" entrycourse="SCM" />
                <RESULT eventid="1188" points="357" swimtime="00:19:54.87" resultid="5714" heatid="7302" lane="7" entrytime="00:19:40.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:44.66" />
                    <SPLIT distance="200" swimtime="00:02:22.93" />
                    <SPLIT distance="250" swimtime="00:03:01.59" />
                    <SPLIT distance="300" swimtime="00:03:40.31" />
                    <SPLIT distance="350" swimtime="00:04:19.96" />
                    <SPLIT distance="400" swimtime="00:04:59.45" />
                    <SPLIT distance="450" swimtime="00:05:39.21" />
                    <SPLIT distance="500" swimtime="00:06:19.44" />
                    <SPLIT distance="550" swimtime="00:06:59.96" />
                    <SPLIT distance="600" swimtime="00:07:39.66" />
                    <SPLIT distance="650" swimtime="00:08:19.81" />
                    <SPLIT distance="700" swimtime="00:09:00.65" />
                    <SPLIT distance="750" swimtime="00:09:41.20" />
                    <SPLIT distance="800" swimtime="00:10:21.97" />
                    <SPLIT distance="850" swimtime="00:11:02.85" />
                    <SPLIT distance="900" swimtime="00:11:43.58" />
                    <SPLIT distance="950" swimtime="00:12:24.04" />
                    <SPLIT distance="1000" swimtime="00:13:05.15" />
                    <SPLIT distance="1050" swimtime="00:13:45.95" />
                    <SPLIT distance="1100" swimtime="00:14:26.59" />
                    <SPLIT distance="1150" swimtime="00:15:07.97" />
                    <SPLIT distance="1200" swimtime="00:15:49.70" />
                    <SPLIT distance="1250" swimtime="00:16:31.46" />
                    <SPLIT distance="1300" swimtime="00:17:12.58" />
                    <SPLIT distance="1350" swimtime="00:17:53.13" />
                    <SPLIT distance="1400" swimtime="00:18:32.35" />
                    <SPLIT distance="1450" swimtime="00:19:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="423" reactiontime="+97" swimtime="00:00:59.83" resultid="5715" heatid="7362" lane="7" entrytime="00:01:00.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="348" reactiontime="+88" swimtime="00:01:11.41" resultid="5716" heatid="7386" lane="3" entrytime="00:01:10.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="352" reactiontime="+88" swimtime="00:00:30.78" resultid="5717" heatid="7445" lane="9" entrytime="00:00:30.21" entrycourse="SCM" />
                <RESULT eventid="1513" points="405" reactiontime="+86" swimtime="00:02:14.22" resultid="5718" heatid="7484" lane="7" entrytime="00:02:15.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="150" swimtime="00:01:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="408" reactiontime="+87" swimtime="00:04:45.94" resultid="5719" heatid="7574" lane="9" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:07.12" />
                    <SPLIT distance="150" swimtime="00:01:43.55" />
                    <SPLIT distance="200" swimtime="00:02:20.26" />
                    <SPLIT distance="250" swimtime="00:02:57.48" />
                    <SPLIT distance="300" swimtime="00:03:34.62" />
                    <SPLIT distance="350" swimtime="00:04:10.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="312" reactiontime="+94" swimtime="00:02:00.49" resultid="6873" heatid="7492" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:01.48" />
                    <SPLIT distance="150" swimtime="00:01:33.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5726" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="5720" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="6497" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="5712" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="264" reactiontime="+69" swimtime="00:02:20.94" resultid="6874" heatid="7403" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5712" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5726" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5720" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="6497" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SMTSZ" nation="POL" region="16" clubid="4461" name="Swimming Masters Team Szczecin">
          <CONTACT city="Mierzyn" email="marekzet74@gmail.com" name="Zienkiewicz Marek" phone="500641651" state="ZACH." street="Teresy 58" zip="72-006" />
          <ATHLETES>
            <ATHLETE birthdate="1987-08-03" firstname="Edyta" gender="F" lastname="Adamiak" nation="POL" athleteid="4472">
              <RESULTS>
                <RESULT eventid="1059" points="177" reactiontime="+97" swimtime="00:00:40.77" resultid="4473" heatid="7237" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1140" points="156" reactiontime="+98" swimtime="00:14:48.95" resultid="4474" heatid="7292" lane="8" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                    <SPLIT distance="150" swimtime="00:02:33.92" />
                    <SPLIT distance="200" swimtime="00:03:31.44" />
                    <SPLIT distance="250" swimtime="00:04:28.67" />
                    <SPLIT distance="300" swimtime="00:05:25.86" />
                    <SPLIT distance="350" swimtime="00:06:22.32" />
                    <SPLIT distance="400" swimtime="00:07:19.29" />
                    <SPLIT distance="450" swimtime="00:08:16.91" />
                    <SPLIT distance="500" swimtime="00:09:13.87" />
                    <SPLIT distance="550" swimtime="00:10:10.87" />
                    <SPLIT distance="600" swimtime="00:11:07.43" />
                    <SPLIT distance="650" swimtime="00:12:04.34" />
                    <SPLIT distance="700" swimtime="00:13:00.93" />
                    <SPLIT distance="750" swimtime="00:13:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="155" reactiontime="+95" swimtime="00:01:33.46" resultid="4475" heatid="7341" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="157" swimtime="00:01:44.72" resultid="4476" heatid="7370" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="200" reactiontime="+95" swimtime="00:00:48.82" resultid="4477" heatid="7540" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1721" points="163" reactiontime="+90" swimtime="00:07:07.89" resultid="4478" heatid="7570" lane="6" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                    <SPLIT distance="100" swimtime="00:01:40.11" />
                    <SPLIT distance="150" swimtime="00:02:35.03" />
                    <SPLIT distance="200" swimtime="00:03:30.22" />
                    <SPLIT distance="250" swimtime="00:04:25.41" />
                    <SPLIT distance="300" swimtime="00:05:20.94" />
                    <SPLIT distance="350" swimtime="00:06:16.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-26" firstname="Magdalena" gender="F" lastname="Bruzgo" nation="POL" athleteid="4537">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="4538" heatid="7237" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4539" heatid="7340" lane="6" entrytime="00:01:55.00" />
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="4540" heatid="7408" lane="3" entrytime="00:02:10.00" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4541" heatid="7468" lane="7" entrytime="00:04:20.00" />
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="4542" heatid="7539" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="4543" heatid="7572" lane="4" entrytime="00:09:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-31" firstname="Joanna" gender="F" lastname="Głuszyk" nation="POL" athleteid="4491">
              <RESULTS>
                <RESULT eventid="1272" points="81" swimtime="00:01:55.81" resultid="4492" heatid="7341" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="86" swimtime="00:08:49.64" resultid="4493" heatid="7571" lane="7" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.54" />
                    <SPLIT distance="100" swimtime="00:01:56.27" />
                    <SPLIT distance="150" swimtime="00:03:02.70" />
                    <SPLIT distance="200" swimtime="00:04:11.91" />
                    <SPLIT distance="250" swimtime="00:05:21.17" />
                    <SPLIT distance="300" swimtime="00:06:32.01" />
                    <SPLIT distance="350" swimtime="00:07:42.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-31" firstname="Izabela" gender="F" lastname="Kowalczyk" nation="POL" athleteid="4494">
              <RESULTS>
                <RESULT eventid="1092" points="313" reactiontime="+95" swimtime="00:02:59.32" resultid="4495" heatid="7274" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:22.67" />
                    <SPLIT distance="150" swimtime="00:02:15.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="284" reactiontime="+90" swimtime="00:00:39.01" resultid="4496" heatid="7310" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1304" points="340" reactiontime="+87" swimtime="00:01:20.93" resultid="4497" heatid="7372" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="311" reactiontime="+92" swimtime="00:00:35.96" resultid="4498" heatid="7431" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="4499" heatid="7472" lane="0" entrytime="00:02:45.00" />
                <RESULT eventid="1608" points="263" reactiontime="+91" swimtime="00:01:25.22" resultid="4500" heatid="7510" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="306" reactiontime="+90" swimtime="00:00:42.37" resultid="4501" heatid="7541" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="4522">
              <RESULTS>
                <RESULT eventid="1059" points="502" reactiontime="+82" swimtime="00:00:28.84" resultid="4523" heatid="7244" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1207" points="532" reactiontime="+82" swimtime="00:00:31.68" resultid="4524" heatid="7314" lane="9" entrytime="00:00:32.50" />
                <RESULT eventid="1304" points="440" reactiontime="+84" swimtime="00:01:14.25" resultid="4525" heatid="7375" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-26" firstname="Grzegorz" gender="M" lastname="Król" nation="POL" athleteid="4534">
              <RESULTS>
                <RESULT eventid="1513" points="140" reactiontime="+82" swimtime="00:03:11.31" resultid="4535" heatid="7477" lane="6" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                    <SPLIT distance="100" swimtime="00:01:28.36" />
                    <SPLIT distance="150" swimtime="00:02:21.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="127" reactiontime="+91" swimtime="00:07:02.00" resultid="4536" heatid="7582" lane="7" entrytime="00:06:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:40.26" />
                    <SPLIT distance="150" swimtime="00:02:34.97" />
                    <SPLIT distance="200" swimtime="00:03:27.92" />
                    <SPLIT distance="250" swimtime="00:04:23.17" />
                    <SPLIT distance="300" swimtime="00:05:18.50" />
                    <SPLIT distance="350" swimtime="00:06:12.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="4462">
              <RESULTS>
                <RESULT eventid="1092" points="349" reactiontime="+74" swimtime="00:02:53.00" resultid="4463" heatid="7275" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:02:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="406" reactiontime="+69" swimtime="00:00:34.65" resultid="4464" heatid="7313" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="4465" heatid="7375" lane="0" entrytime="00:01:15.00" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="4466" heatid="7432" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="4467" heatid="7511" lane="0" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-27" firstname="Marek" gender="M" lastname="Piotrowski" nation="POL" athleteid="4479">
              <RESULTS>
                <RESULT eventid="1689" points="228" reactiontime="+69" swimtime="00:00:41.29" resultid="4480" heatid="7552" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1737" points="224" reactiontime="+72" swimtime="00:05:49.04" resultid="4481" heatid="7580" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:00.18" />
                    <SPLIT distance="200" swimtime="00:02:44.73" />
                    <SPLIT distance="250" swimtime="00:03:30.29" />
                    <SPLIT distance="300" swimtime="00:04:15.30" />
                    <SPLIT distance="350" swimtime="00:05:02.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-02-15" firstname="Filip" gender="M" lastname="Przybyłowski" nation="POL" athleteid="4510">
              <RESULTS>
                <RESULT eventid="1076" points="440" reactiontime="+63" swimtime="00:00:26.62" resultid="4511" heatid="7262" lane="2" entrytime="00:00:27.92" />
                <RESULT eventid="1156" points="352" reactiontime="+73" swimtime="00:10:27.45" resultid="4512" heatid="7295" lane="7" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:48.17" />
                    <SPLIT distance="200" swimtime="00:02:26.34" />
                    <SPLIT distance="250" swimtime="00:03:05.94" />
                    <SPLIT distance="300" swimtime="00:03:45.95" />
                    <SPLIT distance="350" swimtime="00:04:26.10" />
                    <SPLIT distance="400" swimtime="00:05:06.29" />
                    <SPLIT distance="450" swimtime="00:05:46.83" />
                    <SPLIT distance="500" swimtime="00:06:27.44" />
                    <SPLIT distance="550" swimtime="00:07:08.21" />
                    <SPLIT distance="600" swimtime="00:07:48.98" />
                    <SPLIT distance="650" swimtime="00:08:29.75" />
                    <SPLIT distance="700" swimtime="00:09:10.04" />
                    <SPLIT distance="750" swimtime="00:09:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="409" reactiontime="+60" swimtime="00:00:29.30" resultid="4513" heatid="7444" lane="4" entrytime="00:00:30.26" />
                <RESULT eventid="1513" points="404" reactiontime="+62" swimtime="00:02:14.32" resultid="4514" heatid="7483" lane="3" entrytime="00:02:18.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="100" swimtime="00:01:04.92" />
                    <SPLIT distance="150" swimtime="00:01:40.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="396" reactiontime="+63" swimtime="00:01:05.45" resultid="4515" heatid="7518" lane="8" entrytime="00:01:11.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="188" reactiontime="+88" swimtime="00:06:10.38" resultid="4516" heatid="7576" lane="9" entrytime="00:05:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:23.09" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                    <SPLIT distance="200" swimtime="00:03:00.08" />
                    <SPLIT distance="250" swimtime="00:03:48.46" />
                    <SPLIT distance="300" swimtime="00:04:38.18" />
                    <SPLIT distance="350" swimtime="00:05:26.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="4468">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4469" heatid="7258" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4470" heatid="7357" lane="4" entrytime="00:01:07.07" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4471" heatid="7556" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-09" firstname="Łukasz" gender="M" lastname="Rożek" nation="POL" athleteid="4502">
              <RESULTS>
                <RESULT eventid="1156" points="174" swimtime="00:13:13.06" resultid="4503" heatid="7298" lane="0" entrytime="00:13:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:02:11.36" />
                    <SPLIT distance="200" swimtime="00:02:59.42" />
                    <SPLIT distance="250" swimtime="00:03:48.64" />
                    <SPLIT distance="300" swimtime="00:04:38.66" />
                    <SPLIT distance="350" swimtime="00:05:30.06" />
                    <SPLIT distance="400" swimtime="00:06:21.34" />
                    <SPLIT distance="450" swimtime="00:07:12.13" />
                    <SPLIT distance="500" swimtime="00:08:03.76" />
                    <SPLIT distance="550" swimtime="00:08:55.97" />
                    <SPLIT distance="600" swimtime="00:09:48.24" />
                    <SPLIT distance="650" swimtime="00:10:40.84" />
                    <SPLIT distance="700" swimtime="00:11:32.84" />
                    <SPLIT distance="750" swimtime="00:12:24.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="236" reactiontime="+82" swimtime="00:01:12.65" resultid="4504" heatid="7353" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="162" reactiontime="+80" swimtime="00:01:32.08" resultid="4505" heatid="7379" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="200" reactiontime="+75" swimtime="00:00:37.17" resultid="4506" heatid="7438" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1513" points="198" reactiontime="+79" swimtime="00:02:50.48" resultid="4507" heatid="7479" lane="0" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4508" heatid="7549" lane="2" entrytime="00:00:47.00" />
                <RESULT eventid="1737" points="184" reactiontime="+75" swimtime="00:06:12.71" resultid="4509" heatid="7581" lane="3" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:12.14" />
                    <SPLIT distance="200" swimtime="00:02:59.32" />
                    <SPLIT distance="250" swimtime="00:03:47.38" />
                    <SPLIT distance="300" swimtime="00:04:36.73" />
                    <SPLIT distance="350" swimtime="00:05:26.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-30" firstname="Robert" gender="M" lastname="Zając" nation="POL" athleteid="4517">
              <RESULTS>
                <RESULT eventid="1076" points="245" reactiontime="+98" swimtime="00:00:32.35" resultid="4518" heatid="7256" lane="7" entrytime="00:00:31.47" />
                <RESULT eventid="1288" points="196" reactiontime="+97" swimtime="00:01:17.28" resultid="4519" heatid="7356" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="246" reactiontime="+86" swimtime="00:00:34.70" resultid="4520" heatid="7440" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1689" points="219" reactiontime="+97" swimtime="00:00:41.89" resultid="4521" heatid="7553" lane="2" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="4482">
              <RESULTS>
                <RESULT eventid="1092" points="392" reactiontime="+68" swimtime="00:02:46.48" resultid="4483" heatid="7274" lane="6" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                    <SPLIT distance="150" swimtime="00:02:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="371" reactiontime="+80" swimtime="00:11:06.70" resultid="4484" heatid="7290" lane="8" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                    <SPLIT distance="200" swimtime="00:02:39.19" />
                    <SPLIT distance="250" swimtime="00:03:21.40" />
                    <SPLIT distance="300" swimtime="00:04:03.64" />
                    <SPLIT distance="350" swimtime="00:04:46.11" />
                    <SPLIT distance="400" swimtime="00:05:29.24" />
                    <SPLIT distance="450" swimtime="00:06:12.48" />
                    <SPLIT distance="500" swimtime="00:06:55.54" />
                    <SPLIT distance="550" swimtime="00:07:38.34" />
                    <SPLIT distance="600" swimtime="00:08:21.28" />
                    <SPLIT distance="650" swimtime="00:09:04.30" />
                    <SPLIT distance="700" swimtime="00:09:46.53" />
                    <SPLIT distance="750" swimtime="00:10:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="364" reactiontime="+82" swimtime="00:00:35.92" resultid="4485" heatid="7312" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="1304" points="396" reactiontime="+71" swimtime="00:01:16.95" resultid="4486" heatid="7374" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="375" reactiontime="+81" swimtime="00:01:16.29" resultid="4487" heatid="7457" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="403" reactiontime="+70" swimtime="00:02:29.42" resultid="4488" heatid="7472" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="383" reactiontime="+82" swimtime="00:02:44.09" resultid="4489" heatid="7527" lane="5" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:02.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="377" reactiontime="+71" swimtime="00:05:23.55" resultid="4490" heatid="7567" lane="0" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                    <SPLIT distance="150" swimtime="00:01:57.17" />
                    <SPLIT distance="200" swimtime="00:02:38.95" />
                    <SPLIT distance="250" swimtime="00:03:20.95" />
                    <SPLIT distance="300" swimtime="00:04:03.13" />
                    <SPLIT distance="350" swimtime="00:04:44.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="4526">
              <RESULTS>
                <RESULT eventid="1076" points="336" reactiontime="+78" swimtime="00:00:29.14" resultid="4527" heatid="7260" lane="9" entrytime="00:00:28.80" />
                <RESULT eventid="1288" points="267" reactiontime="+72" swimtime="00:01:09.71" resultid="4528" heatid="7357" lane="6" entrytime="00:01:07.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="244" reactiontime="+75" swimtime="00:01:20.41" resultid="4529" heatid="7382" lane="6" entrytime="00:01:19.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="284" reactiontime="+71" swimtime="00:00:33.07" resultid="4530" heatid="7442" lane="2" entrytime="00:00:32.61" />
                <RESULT eventid="1513" points="224" reactiontime="+72" swimtime="00:02:43.59" resultid="4531" heatid="7480" lane="2" entrytime="00:02:39.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                    <SPLIT distance="150" swimtime="00:02:00.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="222" reactiontime="+73" swimtime="00:01:19.40" resultid="4532" heatid="7517" lane="8" entrytime="00:01:16.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="291" reactiontime="+74" swimtime="00:00:38.08" resultid="4533" heatid="7555" lane="1" entrytime="00:00:37.09" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="252" reactiontime="+75" swimtime="00:02:23.11" resultid="4548" heatid="7404" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:51.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4526" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4468" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4517" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4502" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="290" reactiontime="+71" swimtime="00:02:03.47" resultid="4549" heatid="7494" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:36.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4526" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4534" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4517" number="3" reactiontime="+1" />
                    <RELAYPOSITION athleteid="4468" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="409" reactiontime="+83" swimtime="00:02:17.91" resultid="4546" heatid="7401" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:47.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4522" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="4494" number="2" />
                    <RELAYPOSITION athleteid="4462" number="3" />
                    <RELAYPOSITION athleteid="4482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" points="375" reactiontime="+72" swimtime="00:02:10.18" resultid="4547" heatid="7491" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4482" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4472" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4522" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4462" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="277" reactiontime="+79" swimtime="00:02:14.77" resultid="4544" heatid="7288" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:02.24" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4526" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4494" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4472" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4517" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="341" reactiontime="+80" swimtime="00:02:17.86" resultid="4545" heatid="7564" lane="1" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:45.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4522" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4526" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4517" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4494" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ALVSE" nation="CZE" clubid="6466" name="TJ Alcedo Vsetín z.s." shortname="TJ Alcedo Vsetín">
          <CONTACT city="Vsetín" email="tjvs@czechswimming.cz" name="Pavel Obr" state="CZE" street="Dolní Jasenka 770" zip="75501" />
          <ATHLETES>
            <ATHLETE birthdate="1967-05-03" firstname="Pavel" gender="M" lastname="Obr" nation="CZE" athleteid="6467">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="6468" heatid="7261" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="6469" heatid="7278" lane="1" entrytime="00:02:38.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="6470" heatid="7362" lane="0" entrytime="00:01:01.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="6471" heatid="7385" lane="0" entrytime="00:01:13.00" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6472" heatid="7445" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="6473" heatid="7482" lane="5" entrytime="00:02:27.00" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="6474" heatid="7517" lane="3" entrytime="00:01:11.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="6475" heatid="7557" lane="9" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="5072" name="TKKF Masters Koszalin">
          <CONTACT email="rpieslak@wp.pl" name="Pieślak Roman" phone="600227112" />
          <ATHLETES>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="5124">
              <RESULTS>
                <RESULT eventid="1092" points="187" reactiontime="+90" swimtime="00:03:32.85" resultid="5125" heatid="7272" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                    <SPLIT distance="150" swimtime="00:02:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="242" swimtime="00:24:34.16" resultid="5126" heatid="7300" lane="8" entrytime="00:24:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:18.37" />
                    <SPLIT distance="200" swimtime="00:03:07.56" />
                    <SPLIT distance="250" swimtime="00:03:57.23" />
                    <SPLIT distance="300" swimtime="00:04:46.78" />
                    <SPLIT distance="350" swimtime="00:05:36.54" />
                    <SPLIT distance="400" swimtime="00:06:25.99" />
                    <SPLIT distance="450" swimtime="00:07:15.68" />
                    <SPLIT distance="500" swimtime="00:08:05.69" />
                    <SPLIT distance="550" swimtime="00:08:55.11" />
                    <SPLIT distance="600" swimtime="00:09:44.60" />
                    <SPLIT distance="650" swimtime="00:10:34.15" />
                    <SPLIT distance="700" swimtime="00:11:23.61" />
                    <SPLIT distance="750" swimtime="00:12:13.29" />
                    <SPLIT distance="800" swimtime="00:13:02.61" />
                    <SPLIT distance="850" swimtime="00:13:52.50" />
                    <SPLIT distance="900" swimtime="00:14:41.76" />
                    <SPLIT distance="950" swimtime="00:15:31.57" />
                    <SPLIT distance="1000" swimtime="00:16:21.07" />
                    <SPLIT distance="1050" swimtime="00:17:09.80" />
                    <SPLIT distance="1100" swimtime="00:17:59.79" />
                    <SPLIT distance="1150" swimtime="00:18:49.85" />
                    <SPLIT distance="1200" swimtime="00:19:39.44" />
                    <SPLIT distance="1250" swimtime="00:20:28.67" />
                    <SPLIT distance="1300" swimtime="00:21:18.37" />
                    <SPLIT distance="1350" swimtime="00:22:08.08" />
                    <SPLIT distance="1400" swimtime="00:22:57.80" />
                    <SPLIT distance="1450" swimtime="00:23:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="152" reactiontime="+73" swimtime="00:00:48.05" resultid="5127" heatid="7310" lane="0" entrytime="00:00:43.00" />
                <RESULT eventid="1304" points="198" swimtime="00:01:36.88" resultid="5128" heatid="7371" lane="0" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="183" reactiontime="+71" swimtime="00:01:36.81" resultid="5129" heatid="7454" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="204" reactiontime="+96" swimtime="00:07:19.40" resultid="5130" heatid="8150" lane="7" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                    <SPLIT distance="100" swimtime="00:01:46.71" />
                    <SPLIT distance="150" swimtime="00:02:43.41" />
                    <SPLIT distance="200" swimtime="00:03:39.66" />
                    <SPLIT distance="250" swimtime="00:04:39.99" />
                    <SPLIT distance="300" swimtime="00:05:41.80" />
                    <SPLIT distance="350" swimtime="00:06:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="182" reactiontime="+78" swimtime="00:03:30.31" resultid="5131" heatid="7526" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.24" />
                    <SPLIT distance="100" swimtime="00:01:42.82" />
                    <SPLIT distance="150" swimtime="00:02:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="190" reactiontime="+94" swimtime="00:00:49.65" resultid="5132" heatid="7541" lane="9" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-16" firstname="Katarzyna" gender="F" lastname="Gudaniec" nation="POL" athleteid="5133">
              <RESULTS>
                <RESULT eventid="1172" points="372" reactiontime="+81" swimtime="00:21:18.40" resultid="5134" heatid="7300" lane="5" entrytime="00:21:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:53.41" />
                    <SPLIT distance="200" swimtime="00:02:34.35" />
                    <SPLIT distance="250" swimtime="00:03:15.07" />
                    <SPLIT distance="300" swimtime="00:03:56.46" />
                    <SPLIT distance="350" swimtime="00:04:38.17" />
                    <SPLIT distance="400" swimtime="00:05:20.59" />
                    <SPLIT distance="450" swimtime="00:06:02.56" />
                    <SPLIT distance="500" swimtime="00:06:46.01" />
                    <SPLIT distance="550" swimtime="00:07:29.51" />
                    <SPLIT distance="600" swimtime="00:08:12.84" />
                    <SPLIT distance="650" swimtime="00:08:56.41" />
                    <SPLIT distance="700" swimtime="00:09:39.81" />
                    <SPLIT distance="750" swimtime="00:10:23.36" />
                    <SPLIT distance="800" swimtime="00:11:06.76" />
                    <SPLIT distance="850" swimtime="00:11:50.07" />
                    <SPLIT distance="900" swimtime="00:12:33.66" />
                    <SPLIT distance="950" swimtime="00:13:16.95" />
                    <SPLIT distance="1000" swimtime="00:14:00.69" />
                    <SPLIT distance="1050" swimtime="00:14:44.30" />
                    <SPLIT distance="1100" swimtime="00:15:27.89" />
                    <SPLIT distance="1150" swimtime="00:16:11.58" />
                    <SPLIT distance="1200" swimtime="00:16:55.65" />
                    <SPLIT distance="1250" swimtime="00:17:39.09" />
                    <SPLIT distance="1300" swimtime="00:18:22.90" />
                    <SPLIT distance="1350" swimtime="00:19:07.25" />
                    <SPLIT distance="1400" swimtime="00:19:51.52" />
                    <SPLIT distance="1450" swimtime="00:20:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="361" reactiontime="+77" swimtime="00:01:19.36" resultid="5135" heatid="7374" lane="6" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="420" reactiontime="+78" swimtime="00:02:27.41" resultid="5136" heatid="7472" lane="3" entrytime="00:02:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="399" reactiontime="+88" swimtime="00:05:17.55" resultid="5137" heatid="7568" lane="3" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="150" swimtime="00:01:52.97" />
                    <SPLIT distance="200" swimtime="00:02:33.42" />
                    <SPLIT distance="250" swimtime="00:03:14.52" />
                    <SPLIT distance="300" swimtime="00:03:55.63" />
                    <SPLIT distance="350" swimtime="00:04:36.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-08-24" firstname="Karolina" gender="F" lastname="Janas" nation="POL" athleteid="5118">
              <RESULTS>
                <RESULT eventid="1059" points="224" swimtime="00:00:37.74" resultid="5119" heatid="7238" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1207" points="226" reactiontime="+81" swimtime="00:00:42.13" resultid="5120" heatid="7310" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1304" points="225" reactiontime="+99" swimtime="00:01:32.84" resultid="5121" heatid="7370" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="195" reactiontime="+84" swimtime="00:01:34.83" resultid="5122" heatid="7455" lane="7" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="243" swimtime="00:00:45.75" resultid="5123" heatid="7540" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-23" firstname="Witold" gender="M" lastname="Patan" nation="POL" athleteid="5138">
              <RESULTS>
                <RESULT eventid="1076" points="188" reactiontime="+88" swimtime="00:00:35.36" resultid="5139" heatid="7251" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1224" points="71" reactiontime="+82" swimtime="00:00:53.66" resultid="5140" heatid="7318" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1320" points="116" reactiontime="+82" swimtime="00:01:43.02" resultid="5141" heatid="7378" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="149" reactiontime="+80" swimtime="00:01:44.68" resultid="5142" heatid="7417" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="149" reactiontime="+82" swimtime="00:00:47.61" resultid="5143" heatid="7549" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="5107">
              <RESULTS>
                <RESULT eventid="1059" points="302" reactiontime="+83" swimtime="00:00:34.14" resultid="5108" heatid="7239" lane="4" entrytime="00:00:34.30" />
                <RESULT eventid="1207" points="280" reactiontime="+80" swimtime="00:00:39.22" resultid="5109" heatid="7311" lane="8" entrytime="00:00:39.50" />
                <RESULT eventid="1272" points="298" reactiontime="+86" swimtime="00:01:15.21" resultid="5110" heatid="7344" lane="7" entrytime="00:01:16.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="260" reactiontime="+79" swimtime="00:01:26.14" resultid="5111" heatid="7456" lane="9" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="254" reactiontime="+86" swimtime="00:03:08.16" resultid="5112" heatid="7526" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:30.91" />
                    <SPLIT distance="150" swimtime="00:02:20.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="5087">
              <RESULTS>
                <RESULT eventid="1059" points="320" swimtime="00:00:33.49" resultid="5088" heatid="7242" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1272" points="317" reactiontime="+98" swimtime="00:01:13.64" resultid="5089" heatid="7345" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="5090" heatid="7410" lane="7" entrytime="00:01:45.00" />
                <RESULT eventid="1497" points="297" reactiontime="+87" swimtime="00:02:45.41" resultid="5091" heatid="7471" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:02.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="5092" heatid="7542" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="1721" points="287" reactiontime="+96" swimtime="00:05:54.53" resultid="5093" heatid="7568" lane="7" entrytime="00:05:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:06.42" />
                    <SPLIT distance="200" swimtime="00:02:52.93" />
                    <SPLIT distance="250" swimtime="00:03:39.11" />
                    <SPLIT distance="300" swimtime="00:04:25.81" />
                    <SPLIT distance="350" swimtime="00:05:12.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-28" firstname="Roman" gender="M" lastname="Pieślak" nation="POL" athleteid="5094">
              <RESULTS>
                <RESULT eventid="1076" points="341" reactiontime="+75" swimtime="00:00:28.98" resultid="5095" heatid="7259" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1256" points="335" reactiontime="+74" swimtime="00:02:52.86" resultid="5096" heatid="7338" lane="9" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:22.65" />
                    <SPLIT distance="150" swimtime="00:02:07.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="340" reactiontime="+73" swimtime="00:01:04.34" resultid="5097" heatid="7360" lane="0" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="368" reactiontime="+70" swimtime="00:01:17.58" resultid="5098" heatid="7422" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="325" reactiontime="+72" swimtime="00:02:24.44" resultid="5099" heatid="7482" lane="4" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="365" reactiontime="+77" swimtime="00:00:35.31" resultid="5100" heatid="7557" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5101" heatid="7578" lane="8" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-06" firstname="Joanna" gender="F" lastname="Stankiewicz-Majkowska" nation="POL" athleteid="5113">
              <RESULTS>
                <RESULT eventid="1092" points="214" reactiontime="+91" swimtime="00:03:23.69" resultid="5114" heatid="7273" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:02:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="171" swimtime="00:03:35.35" resultid="5115" heatid="7392" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                    <SPLIT distance="100" swimtime="00:01:40.51" />
                    <SPLIT distance="150" swimtime="00:02:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="210" reactiontime="+98" swimtime="00:07:15.21" resultid="5116" heatid="8150" lane="1" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:41.06" />
                    <SPLIT distance="150" swimtime="00:02:37.01" />
                    <SPLIT distance="200" swimtime="00:03:32.18" />
                    <SPLIT distance="250" swimtime="00:04:30.08" />
                    <SPLIT distance="300" swimtime="00:05:28.62" />
                    <SPLIT distance="350" swimtime="00:06:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="219" reactiontime="+86" swimtime="00:00:47.37" resultid="5117" heatid="7540" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1240" points="242" swimtime="00:03:35.87" resultid="6301" heatid="7330" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:43.58" />
                    <SPLIT distance="150" swimtime="00:02:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-14" firstname="Leszek" gender="M" lastname="Szwed" nation="POL" athleteid="5081">
              <RESULTS>
                <RESULT eventid="1076" points="83" reactiontime="+50" swimtime="00:00:46.38" resultid="5082" heatid="7248" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1224" points="84" swimtime="00:00:50.63" resultid="5083" heatid="7318" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5084" heatid="7351" lane="0" entrytime="00:01:41.00" />
                <RESULT eventid="1481" points="85" swimtime="00:01:51.07" resultid="5085" heatid="7461" lane="7" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="78" reactiontime="+78" swimtime="00:04:06.94" resultid="5086" heatid="7530" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.20" />
                    <SPLIT distance="100" swimtime="00:02:01.40" />
                    <SPLIT distance="150" swimtime="00:04:06.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-16" firstname="Dawid" gender="M" lastname="Wróblewski" nation="POL" athleteid="5144">
              <RESULTS>
                <RESULT eventid="1076" points="580" reactiontime="+73" swimtime="00:00:24.29" resultid="5145" heatid="7268" lane="8" entrytime="00:00:25.50" />
                <RESULT eventid="1108" points="495" reactiontime="+77" swimtime="00:02:18.52" resultid="5146" heatid="7285" lane="9" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:46.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="526" reactiontime="+76" swimtime="00:02:28.79" resultid="5147" heatid="7339" lane="1" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:50.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5148" heatid="7365" lane="5" entrytime="00:00:56.50" />
                <RESULT eventid="1449" points="564" reactiontime="+69" swimtime="00:00:26.32" resultid="5149" heatid="7449" lane="5" entrytime="00:00:27.15" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5150" heatid="7486" lane="1" entrytime="00:02:10.00" />
                <RESULT eventid="1625" points="546" reactiontime="+74" swimtime="00:00:58.80" resultid="5151" heatid="7521" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="477" reactiontime="+72" swimtime="00:04:31.56" resultid="5152" heatid="7573" lane="9" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                    <SPLIT distance="150" swimtime="00:01:39.96" />
                    <SPLIT distance="200" swimtime="00:02:14.22" />
                    <SPLIT distance="250" swimtime="00:02:48.19" />
                    <SPLIT distance="300" swimtime="00:03:22.76" />
                    <SPLIT distance="350" swimtime="00:03:57.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-04-14" firstname="Wiesław" gender="M" lastname="Załuski" nation="POL" athleteid="5102">
              <RESULTS>
                <RESULT eventid="1108" points="232" swimtime="00:02:58.37" resultid="5103" heatid="7280" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="150" swimtime="00:02:15.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="264" reactiontime="+85" swimtime="00:01:18.34" resultid="5104" heatid="7382" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="237" reactiontime="+70" swimtime="00:00:35.12" resultid="5105" heatid="7440" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1625" points="164" reactiontime="+90" swimtime="00:01:27.81" resultid="5106" heatid="7516" lane="0" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="5073">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="5074" heatid="7281" lane="3" entrytime="00:02:45.00" />
                <RESULT eventid="1188" points="261" reactiontime="+89" swimtime="00:22:06.51" resultid="5075" heatid="7303" lane="5" entrytime="00:21:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:02:03.14" />
                    <SPLIT distance="200" swimtime="00:02:46.91" />
                    <SPLIT distance="250" swimtime="00:03:30.84" />
                    <SPLIT distance="300" swimtime="00:04:14.60" />
                    <SPLIT distance="350" swimtime="00:04:58.31" />
                    <SPLIT distance="400" swimtime="00:05:41.60" />
                    <SPLIT distance="450" swimtime="00:06:24.60" />
                    <SPLIT distance="500" swimtime="00:07:07.50" />
                    <SPLIT distance="550" swimtime="00:07:50.59" />
                    <SPLIT distance="600" swimtime="00:08:33.58" />
                    <SPLIT distance="650" swimtime="00:09:17.54" />
                    <SPLIT distance="700" swimtime="00:10:01.59" />
                    <SPLIT distance="750" swimtime="00:10:45.62" />
                    <SPLIT distance="800" swimtime="00:11:30.49" />
                    <SPLIT distance="850" swimtime="00:12:15.32" />
                    <SPLIT distance="900" swimtime="00:13:00.49" />
                    <SPLIT distance="950" swimtime="00:13:46.35" />
                    <SPLIT distance="1000" swimtime="00:14:32.31" />
                    <SPLIT distance="1050" swimtime="00:15:18.46" />
                    <SPLIT distance="1100" swimtime="00:16:04.47" />
                    <SPLIT distance="1150" swimtime="00:16:50.62" />
                    <SPLIT distance="1200" swimtime="00:17:36.97" />
                    <SPLIT distance="1250" swimtime="00:18:22.96" />
                    <SPLIT distance="1300" swimtime="00:19:09.46" />
                    <SPLIT distance="1350" swimtime="00:19:55.91" />
                    <SPLIT distance="1400" swimtime="00:20:41.99" />
                    <SPLIT distance="1450" swimtime="00:21:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="243" reactiontime="+66" swimtime="00:00:35.57" resultid="5076" heatid="7323" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1320" points="319" reactiontime="+76" swimtime="00:01:13.55" resultid="5077" heatid="7384" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="315" reactiontime="+67" swimtime="00:01:11.77" resultid="5078" heatid="7464" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="277" reactiontime="+66" swimtime="00:02:41.98" resultid="5079" heatid="7533" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:19.36" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5080" heatid="7577" lane="7" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="TKKF Koszalin 4" number="4">
              <RESULTS>
                <RESULT eventid="1391" points="383" reactiontime="+74" swimtime="00:02:04.43" resultid="5156" heatid="7405" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:07.79" />
                    <SPLIT distance="150" swimtime="00:01:33.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5073" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5094" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="5144" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="5102" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="TKKF Koszalin 6" number="6">
              <RESULTS>
                <RESULT eventid="1545" status="WDR" swimtime="00:00:00.00" resultid="5158" heatid="7495" lane="0" entrytime="00:01:54.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5094" number="1" />
                    <RELAYPOSITION athleteid="5073" number="2" />
                    <RELAYPOSITION athleteid="5102" number="3" />
                    <RELAYPOSITION athleteid="5144" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="TKKF Koszalin 3" number="3">
              <RESULTS>
                <RESULT eventid="1368" points="292" reactiontime="+78" swimtime="00:02:34.29" resultid="5155" heatid="7400" lane="5" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5107" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5113" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="5133" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5087" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="TKKF Koszalin 5" number="5">
              <RESULTS>
                <RESULT eventid="1529" points="337" reactiontime="+85" swimtime="00:02:14.91" resultid="5157" heatid="7490" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:43.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5107" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5133" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="5124" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="5087" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="TKKF Koszalin 1" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="425" reactiontime="+80" swimtime="00:01:56.86" resultid="5153" heatid="7288" lane="4" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:00.20" />
                    <SPLIT distance="150" swimtime="00:01:32.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5133" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5094" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="5087" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="5144" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TKKF Koszalin 2" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="195" reactiontime="+95" swimtime="00:02:31.39" resultid="5154" heatid="7287" lane="6" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                    <SPLIT distance="150" swimtime="00:01:55.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5081" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="5107" number="2" reactiontime="+2" />
                    <RELAYPOSITION athleteid="5118" number="3" reactiontime="-3" />
                    <RELAYPOSITION athleteid="5138" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="TKKF Koszalin 7" number="7">
              <RESULTS>
                <RESULT eventid="1705" status="DNS" swimtime="00:00:00.00" resultid="5159" heatid="7564" lane="4" entrytime="00:02:11.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5133" number="1" />
                    <RELAYPOSITION athleteid="5094" number="2" />
                    <RELAYPOSITION athleteid="5144" number="3" />
                    <RELAYPOSITION athleteid="5087" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="TKKF Koszalin 8" number="8">
              <RESULTS>
                <RESULT eventid="1705" points="280" reactiontime="+61" swimtime="00:02:27.22" resultid="5161" heatid="7563" lane="4" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:19.20" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5073" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5113" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="5102" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="5107" number="4" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TKKF Koszalin 9" number="9">
              <RESULTS>
                <RESULT eventid="1705" points="157" reactiontime="+85" swimtime="00:02:58.33" resultid="5160" heatid="7563" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:22.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5081" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5118" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5124" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="5138" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05815" nation="POL" region="15" clubid="3954" name="TM Barracuda Kalisz" shortname="Barracuda Kalisz">
          <CONTACT city="KALISZ" email="GALCZYNSKIWOJ@OP.PL" name="GAŁCZYŃSKI WOJCIECH" phone="790690666" state="WLKP" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1996-02-28" firstname="Adam" gender="M" lastname="Białożył" nation="POL" athleteid="3974">
              <RESULTS>
                <RESULT eventid="1076" points="328" reactiontime="+89" swimtime="00:00:29.35" resultid="3975" heatid="7260" lane="2" entrytime="00:00:28.52" />
                <RESULT eventid="1256" points="306" reactiontime="+83" swimtime="00:02:58.17" resultid="3976" heatid="7339" lane="9" entrytime="00:02:42.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:09.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="282" reactiontime="+83" swimtime="00:01:16.62" resultid="3977" heatid="7386" lane="5" entrytime="00:01:10.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="343" reactiontime="+83" swimtime="00:01:19.43" resultid="3978" heatid="7424" lane="6" entrytime="00:01:13.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="269" reactiontime="+87" swimtime="00:02:33.91" resultid="3979" heatid="7481" lane="3" entrytime="00:02:30.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="359" reactiontime="+78" swimtime="00:00:35.51" resultid="3980" heatid="7558" lane="3" entrytime="00:00:34.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-23" firstname="Justyna" gender="F" lastname="Dominiak" nation="POL" athleteid="4022">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="4023" heatid="7241" lane="8" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:02:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="241" reactiontime="+91" swimtime="00:12:49.56" resultid="4024" heatid="7291" lane="6" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:11.70" />
                    <SPLIT distance="200" swimtime="00:02:59.77" />
                    <SPLIT distance="250" swimtime="00:03:49.01" />
                    <SPLIT distance="300" swimtime="00:04:37.95" />
                    <SPLIT distance="350" swimtime="00:05:27.11" />
                    <SPLIT distance="400" swimtime="00:06:17.06" />
                    <SPLIT distance="450" swimtime="00:07:06.27" />
                    <SPLIT distance="500" swimtime="00:07:55.24" />
                    <SPLIT distance="550" swimtime="00:08:44.94" />
                    <SPLIT distance="600" swimtime="00:09:34.19" />
                    <SPLIT distance="650" swimtime="00:10:23.24" />
                    <SPLIT distance="700" swimtime="00:11:12.33" />
                    <SPLIT distance="750" swimtime="00:12:01.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="239" reactiontime="+83" swimtime="00:03:36.67" resultid="4025" heatid="7331" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:41.21" />
                    <SPLIT distance="150" swimtime="00:02:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="4026" heatid="7371" lane="7" entrytime="00:01:35.00" />
                <RESULT eventid="1400" points="245" reactiontime="+77" swimtime="00:01:39.57" resultid="4027" heatid="7411" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="247" reactiontime="+80" swimtime="00:02:55.96" resultid="4028" heatid="7470" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" status="DNS" swimtime="00:00:00.00" resultid="4029" heatid="7543" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1721" status="WDR" swimtime="00:00:00.00" resultid="4030" heatid="7568" lane="0" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-07" firstname="Arkadiusz" gender="M" lastname="Figiel" nation="POL" athleteid="3962">
              <RESULTS>
                <RESULT eventid="1076" points="127" reactiontime="+99" swimtime="00:00:40.21" resultid="3963" heatid="7250" lane="1" entrytime="00:00:39.55" />
                <RESULT eventid="1224" points="83" swimtime="00:00:50.79" resultid="3964" heatid="7317" lane="2" entrytime="00:00:55.93" />
                <RESULT eventid="1320" points="93" swimtime="00:01:50.67" resultid="3965" heatid="7378" lane="1" entrytime="00:01:54.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="135" reactiontime="+94" swimtime="00:01:48.19" resultid="3966" heatid="7416" lane="6" entrytime="00:01:56.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="70" swimtime="00:01:58.17" resultid="3967" heatid="7461" lane="9" entrytime="00:02:01.00" />
                <RESULT eventid="1657" points="66" swimtime="00:04:20.26" resultid="3968" heatid="7529" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.15" />
                    <SPLIT distance="100" swimtime="00:02:07.18" />
                    <SPLIT distance="150" swimtime="00:03:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="155" reactiontime="+94" swimtime="00:00:46.91" resultid="3969" heatid="7548" lane="5" entrytime="00:00:49.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-10-29" firstname="Marzena" gender="F" lastname="Figiel" nation="POL" athleteid="3970">
              <RESULTS>
                <RESULT eventid="1240" points="106" swimtime="00:04:44.11" resultid="3971" heatid="7328" lane="9" entrytime="00:04:46.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.87" />
                    <SPLIT distance="100" swimtime="00:02:18.01" />
                    <SPLIT distance="150" swimtime="00:03:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="50" swimtime="00:02:15.80" resultid="3972" heatid="7340" lane="3" entrytime="00:02:25.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="99" swimtime="00:02:14.72" resultid="3973" heatid="7408" lane="1" entrytime="00:02:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-02" firstname="Anna" gender="F" lastname="Gałczyńska" nation="POL" athleteid="3981">
              <RESULTS>
                <RESULT eventid="1207" points="45" swimtime="00:01:11.88" resultid="3982" heatid="7307" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="1400" points="93" swimtime="00:02:17.42" resultid="3983" heatid="7407" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="53" swimtime="00:02:26.17" resultid="3984" heatid="7453" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="84" swimtime="00:01:05.10" resultid="3985" heatid="7537" lane="4" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-30" firstname="Magdalena" gender="F" lastname="Kolera" nation="POL" athleteid="4006">
              <RESULTS>
                <RESULT eventid="1207" points="218" reactiontime="+88" swimtime="00:00:42.63" resultid="4007" heatid="7310" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1433" status="WDR" swimtime="00:00:00.00" resultid="4008" heatid="7428" lane="9" entrytime="00:00:46.00" />
                <RESULT eventid="1465" points="195" reactiontime="+93" swimtime="00:01:34.86" resultid="4009" heatid="7454" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="182" reactiontime="+98" swimtime="00:03:30.38" resultid="4010" heatid="7525" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                    <SPLIT distance="100" swimtime="00:01:42.52" />
                    <SPLIT distance="150" swimtime="00:02:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-24" firstname="Zofia" gender="F" lastname="Koźlik" nation="POL" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3956" heatid="7235" lane="1" entrytime="00:01:00.36" />
                <RESULT eventid="1207" points="95" reactiontime="+74" swimtime="00:00:56.13" resultid="3957" heatid="7307" lane="0" />
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach. (Time: 11:57)" eventid="1304" status="DSQ" swimtime="00:02:06.26" resultid="3958" heatid="7369" lane="0" entrytime="00:02:08.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="136" reactiontime="+93" swimtime="00:02:01.00" resultid="3959" heatid="7408" lane="4" entrytime="00:02:03.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="58" reactiontime="+98" swimtime="00:01:02.67" resultid="3960" heatid="7426" lane="4" entrytime="00:01:02.20" />
                <RESULT eventid="1673" points="144" swimtime="00:00:54.40" resultid="3961" heatid="7538" lane="5" entrytime="00:00:55.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-09" firstname="Wiktor" gender="M" lastname="Morozowski" nation="POL" athleteid="4000">
              <RESULTS>
                <RESULT eventid="1188" points="211" swimtime="00:23:44.36" resultid="4001" heatid="7303" lane="0" entrytime="00:23:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                    <SPLIT distance="150" swimtime="00:02:03.94" />
                    <SPLIT distance="200" swimtime="00:02:50.19" />
                    <SPLIT distance="250" swimtime="00:03:37.32" />
                    <SPLIT distance="300" swimtime="00:04:25.16" />
                    <SPLIT distance="350" swimtime="00:05:13.11" />
                    <SPLIT distance="400" swimtime="00:06:00.92" />
                    <SPLIT distance="450" swimtime="00:06:48.93" />
                    <SPLIT distance="500" swimtime="00:07:37.40" />
                    <SPLIT distance="550" swimtime="00:08:25.79" />
                    <SPLIT distance="600" swimtime="00:09:14.11" />
                    <SPLIT distance="650" swimtime="00:10:02.72" />
                    <SPLIT distance="700" swimtime="00:10:51.90" />
                    <SPLIT distance="750" swimtime="00:11:41.13" />
                    <SPLIT distance="800" swimtime="00:12:29.62" />
                    <SPLIT distance="850" swimtime="00:13:17.56" />
                    <SPLIT distance="900" swimtime="00:14:05.61" />
                    <SPLIT distance="950" swimtime="00:14:54.36" />
                    <SPLIT distance="1000" swimtime="00:15:43.19" />
                    <SPLIT distance="1050" swimtime="00:16:30.90" />
                    <SPLIT distance="1100" swimtime="00:17:19.36" />
                    <SPLIT distance="1150" swimtime="00:18:07.83" />
                    <SPLIT distance="1200" swimtime="00:18:56.99" />
                    <SPLIT distance="1250" swimtime="00:19:46.05" />
                    <SPLIT distance="1300" swimtime="00:20:34.47" />
                    <SPLIT distance="1350" swimtime="00:21:23.39" />
                    <SPLIT distance="1400" swimtime="00:22:10.81" />
                    <SPLIT distance="1450" swimtime="00:22:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="234" swimtime="00:03:14.92" resultid="4002" heatid="7336" lane="2" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:01:32.07" />
                    <SPLIT distance="150" swimtime="00:02:23.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="222" swimtime="00:01:23.00" resultid="4003" heatid="7381" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="252" swimtime="00:01:28.02" resultid="4004" heatid="7420" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="284" reactiontime="+96" swimtime="00:00:38.37" resultid="4005" heatid="7554" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-20" firstname="Artur" gender="M" lastname="Nowacki" nation="POL" athleteid="3992">
              <RESULTS>
                <RESULT eventid="1076" points="145" swimtime="00:00:38.50" resultid="3993" heatid="7250" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1256" points="171" swimtime="00:03:36.47" resultid="3994" heatid="7336" lane="1" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.04" />
                    <SPLIT distance="100" swimtime="00:01:42.20" />
                    <SPLIT distance="150" swimtime="00:02:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="105" swimtime="00:01:35.18" resultid="3995" heatid="7353" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="182" swimtime="00:01:38.09" resultid="3996" heatid="7418" lane="1" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="81" reactiontime="+87" swimtime="00:03:49.19" resultid="3997" heatid="7479" lane="7" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="100" swimtime="00:01:47.12" />
                    <SPLIT distance="150" swimtime="00:02:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="190" reactiontime="+96" swimtime="00:00:43.91" resultid="3998" heatid="7550" lane="0" entrytime="00:00:45.05" />
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="3999" heatid="7575" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-12" firstname="Karolina" gender="F" lastname="Radomska" nation="POL" athleteid="4011">
              <RESULTS>
                <RESULT eventid="1059" points="260" reactiontime="+91" swimtime="00:00:35.89" resultid="4012" heatid="7239" lane="2" entrytime="00:00:35.15" />
                <RESULT eventid="1140" points="185" reactiontime="+96" swimtime="00:14:01.07" resultid="4013" heatid="7292" lane="7" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.35" />
                    <SPLIT distance="100" swimtime="00:01:38.24" />
                    <SPLIT distance="150" swimtime="00:02:29.23" />
                    <SPLIT distance="200" swimtime="00:03:22.37" />
                    <SPLIT distance="250" swimtime="00:04:14.78" />
                    <SPLIT distance="300" swimtime="00:05:09.26" />
                    <SPLIT distance="350" swimtime="00:06:02.89" />
                    <SPLIT distance="400" swimtime="00:06:56.50" />
                    <SPLIT distance="450" swimtime="00:07:51.75" />
                    <SPLIT distance="500" swimtime="00:08:48.06" />
                    <SPLIT distance="550" swimtime="00:09:45.16" />
                    <SPLIT distance="600" swimtime="00:10:37.43" />
                    <SPLIT distance="650" swimtime="00:11:29.15" />
                    <SPLIT distance="700" swimtime="00:12:20.99" />
                    <SPLIT distance="750" swimtime="00:13:12.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-27" firstname="Małgorzata" gender="F" lastname="Rembowska-Świeboda" nation="POL" athleteid="3986">
              <RESULTS>
                <RESULT eventid="1059" points="347" reactiontime="+76" swimtime="00:00:32.63" resultid="3987" heatid="7241" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1207" points="333" reactiontime="+81" swimtime="00:00:37.00" resultid="3988" heatid="7311" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1304" points="314" reactiontime="+78" swimtime="00:01:23.06" resultid="3989" heatid="7373" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="249" reactiontime="+81" swimtime="00:00:38.74" resultid="3990" heatid="7430" lane="9" entrytime="00:00:37.50" />
                <RESULT eventid="1465" points="308" reactiontime="+80" swimtime="00:01:21.48" resultid="3991" heatid="7456" lane="3" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-11" firstname="Patrycja" gender="F" lastname="Rupa" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1059" points="459" reactiontime="+69" swimtime="00:00:29.71" resultid="4015" heatid="7244" lane="7" entrytime="00:00:29.73" />
                <RESULT eventid="1140" status="DNF" swimtime="00:00:00.00" resultid="4016" heatid="7291" lane="5" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="150" swimtime="00:02:02.98" />
                    <SPLIT distance="200" swimtime="00:02:45.95" />
                    <SPLIT distance="250" swimtime="00:03:38.81" />
                    <SPLIT distance="300" swimtime="00:04:21.61" />
                    <SPLIT distance="350" swimtime="00:05:05.30" />
                    <SPLIT distance="400" swimtime="00:07:43.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="459" reactiontime="+59" swimtime="00:00:33.26" resultid="4017" heatid="7314" lane="8" entrytime="00:00:32.15" />
                <RESULT eventid="1304" points="425" reactiontime="+67" swimtime="00:01:15.14" resultid="4018" heatid="7374" lane="4" entrytime="00:01:15.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="450" reactiontime="+64" swimtime="00:01:11.78" resultid="4019" heatid="7457" lane="4" entrytime="00:01:12.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="413" reactiontime="+63" swimtime="00:02:40.07" resultid="4020" heatid="7528" lane="9" entrytime="00:02:40.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:18.47" />
                    <SPLIT distance="150" swimtime="00:01:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="361" reactiontime="+65" swimtime="00:00:40.10" resultid="4021" heatid="7542" lane="2" entrytime="00:00:42.13" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1368" points="184" reactiontime="+89" swimtime="00:02:59.77" resultid="4033" heatid="7400" lane="6" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:19.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4006" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3981" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="3986" number="3" />
                    <RELAYPOSITION athleteid="4022" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" status="WDR" swimtime="00:00:00.00" resultid="4034" heatid="7490" lane="7" entrytime="00:02:32.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4022" number="1" />
                    <RELAYPOSITION athleteid="3981" number="2" />
                    <RELAYPOSITION athleteid="4006" number="3" />
                    <RELAYPOSITION athleteid="3986" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="258" reactiontime="+99" swimtime="00:02:18.02" resultid="4031" heatid="7287" lane="2" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:45.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3962" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="4011" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="4000" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3986" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1705" points="249" reactiontime="+92" swimtime="00:02:33.21" resultid="4032" heatid="7563" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:25.73" />
                    <SPLIT distance="150" swimtime="00:02:00.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4006" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3992" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4000" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3986" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TORMA" nation="LTU" clubid="5162" name="Torpedos Marijampole">
          <CONTACT city="Marijampole" email="vilmantasenator@gmail.com" name="Vilmantas Krasauskas" phone="+37068746068" street="Jukneviciaus 78-10" />
          <ATHLETES>
            <ATHLETE birthdate="1941-03-14" firstname="Stasys" gender="M" lastname="Grigas" nation="LTU" athleteid="5172">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5173" heatid="7247" lane="5" entrytime="00:00:54.50" entrycourse="SCM" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="5174" heatid="7316" lane="3" entrytime="00:01:10.73" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5175" heatid="7350" lane="7" entrytime="00:02:17.71" entrycourse="SCM" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="5176" heatid="7460" lane="0" entrytime="00:02:34.31" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5177" heatid="7475" lane="3" entrytime="00:05:48.31" entrycourse="SCM" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5178" heatid="7529" lane="3" entrytime="00:05:30.55" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5179" heatid="7547" lane="0" entrytime="00:01:01.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-07-09" firstname="Antanas" gender="M" lastname="Guoga" nation="LTU" athleteid="5163">
              <RESULTS>
                <RESULT eventid="1108" points="95" swimtime="00:03:59.69" resultid="5164" heatid="7278" lane="2" entrytime="00:04:00.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.15" />
                    <SPLIT distance="100" swimtime="00:02:03.29" />
                    <SPLIT distance="150" swimtime="00:03:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="121" swimtime="00:14:54.93" resultid="5165" heatid="7299" lane="1" entrytime="00:15:41.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.76" />
                    <SPLIT distance="100" swimtime="00:01:44.14" />
                    <SPLIT distance="150" swimtime="00:02:39.54" />
                    <SPLIT distance="200" swimtime="00:03:35.52" />
                    <SPLIT distance="250" swimtime="00:04:31.50" />
                    <SPLIT distance="300" swimtime="00:05:27.68" />
                    <SPLIT distance="350" swimtime="00:06:23.94" />
                    <SPLIT distance="400" swimtime="00:07:20.13" />
                    <SPLIT distance="450" swimtime="00:08:16.83" />
                    <SPLIT distance="500" swimtime="00:09:13.49" />
                    <SPLIT distance="550" swimtime="00:10:10.45" />
                    <SPLIT distance="600" swimtime="00:11:07.94" />
                    <SPLIT distance="650" swimtime="00:12:05.19" />
                    <SPLIT distance="700" swimtime="00:13:02.29" />
                    <SPLIT distance="750" swimtime="00:13:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="99" swimtime="00:04:19.62" resultid="5166" heatid="7333" lane="8" entrytime="00:04:35.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.03" />
                    <SPLIT distance="100" swimtime="00:02:03.84" />
                    <SPLIT distance="150" swimtime="00:03:12.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" status="DNS" swimtime="00:00:00.00" resultid="5167" heatid="7394" lane="5" entrytime="00:04:49.16" entrycourse="SCM" />
                <RESULT eventid="1417" points="99" reactiontime="+67" swimtime="00:01:59.84" resultid="5168" heatid="7415" lane="6" entrytime="00:02:14.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="102" reactiontime="+95" swimtime="00:08:23.95" resultid="5169" heatid="8154" lane="6" entrytime="00:08:40.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.10" />
                    <SPLIT distance="100" swimtime="00:02:11.12" />
                    <SPLIT distance="150" swimtime="00:03:16.85" />
                    <SPLIT distance="200" swimtime="00:04:22.95" />
                    <SPLIT distance="250" swimtime="00:05:29.88" />
                    <SPLIT distance="300" swimtime="00:06:37.34" />
                    <SPLIT distance="350" swimtime="00:07:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="63" reactiontime="+94" swimtime="00:02:00.43" resultid="5170" heatid="7513" lane="1" entrytime="00:02:15.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="5171" heatid="7582" lane="9" entrytime="00:07:04.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-07-31" firstname="Vilmantas" gender="M" lastname="Krasauskas" nation="LTU" athleteid="5180">
              <RESULTS>
                <RESULT eventid="1076" points="357" reactiontime="+85" swimtime="00:00:28.54" resultid="5181" heatid="7259" lane="7" entrytime="00:00:29.01" entrycourse="SCM" />
                <RESULT eventid="1188" points="326" reactiontime="+85" swimtime="00:20:31.81" resultid="5182" heatid="7302" lane="9" entrytime="00:20:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:02:32.94" />
                    <SPLIT distance="250" swimtime="00:03:12.59" />
                    <SPLIT distance="300" swimtime="00:03:52.74" />
                    <SPLIT distance="350" swimtime="00:04:32.88" />
                    <SPLIT distance="400" swimtime="00:05:13.16" />
                    <SPLIT distance="450" swimtime="00:05:54.05" />
                    <SPLIT distance="500" swimtime="00:06:35.11" />
                    <SPLIT distance="550" swimtime="00:07:16.23" />
                    <SPLIT distance="600" swimtime="00:07:57.37" />
                    <SPLIT distance="650" swimtime="00:08:38.42" />
                    <SPLIT distance="700" swimtime="00:09:19.72" />
                    <SPLIT distance="750" swimtime="00:10:01.63" />
                    <SPLIT distance="800" swimtime="00:10:43.29" />
                    <SPLIT distance="850" swimtime="00:11:25.15" />
                    <SPLIT distance="900" swimtime="00:12:07.75" />
                    <SPLIT distance="950" swimtime="00:12:49.85" />
                    <SPLIT distance="1000" swimtime="00:13:31.76" />
                    <SPLIT distance="1050" swimtime="00:14:14.73" />
                    <SPLIT distance="1100" swimtime="00:14:56.81" />
                    <SPLIT distance="1150" swimtime="00:15:39.26" />
                    <SPLIT distance="1200" swimtime="00:16:21.45" />
                    <SPLIT distance="1250" swimtime="00:17:03.47" />
                    <SPLIT distance="1300" swimtime="00:17:45.66" />
                    <SPLIT distance="1350" swimtime="00:18:27.49" />
                    <SPLIT distance="1400" swimtime="00:19:09.90" />
                    <SPLIT distance="1450" swimtime="00:19:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="386" reactiontime="+79" swimtime="00:01:01.72" resultid="5183" heatid="7361" lane="9" entrytime="00:01:02.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="362" reactiontime="+81" swimtime="00:02:19.31" resultid="5184" heatid="7483" lane="4" entrytime="00:02:18.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="261" reactiontime="+87" swimtime="00:01:15.23" resultid="5185" heatid="7516" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5186" heatid="7553" lane="8" entrytime="00:00:39.53" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="3850" name="TP Masters Opole" shortname="Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="3867">
              <RESULTS>
                <RESULT eventid="1059" points="473" reactiontime="+79" swimtime="00:00:29.42" resultid="3868" heatid="7239" lane="1" entrytime="00:00:35.40" />
                <RESULT eventid="1092" points="454" reactiontime="+80" swimtime="00:02:38.47" resultid="3869" heatid="7275" lane="7" entrytime="00:02:38.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:02:01.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="561" reactiontime="+63" swimtime="00:00:31.11" resultid="3870" heatid="7313" lane="4" entrytime="00:00:32.85" />
                <RESULT eventid="1304" points="508" reactiontime="+77" swimtime="00:01:10.82" resultid="3871" heatid="7375" lane="2" entrytime="00:01:13.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="432" reactiontime="+70" swimtime="00:00:32.24" resultid="3872" heatid="7430" lane="5" entrytime="00:00:36.80" />
                <RESULT eventid="1465" points="523" reactiontime="+70" swimtime="00:01:08.27" resultid="3873" heatid="7458" lane="6" entrytime="00:01:08.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="514" reactiontime="+57" swimtime="00:02:28.78" resultid="3874" heatid="7528" lane="5" entrytime="00:02:28.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="3851">
              <RESULTS>
                <RESULT eventid="1076" points="394" reactiontime="+81" swimtime="00:00:27.63" resultid="3852" heatid="7255" lane="8" entrytime="00:00:32.55" />
                <RESULT eventid="1108" points="384" reactiontime="+86" swimtime="00:02:30.80" resultid="3853" heatid="7282" lane="2" entrytime="00:02:37.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="390" reactiontime="+76" swimtime="00:00:30.41" resultid="3854" heatid="7324" lane="0" entrytime="00:00:32.78" />
                <RESULT eventid="1320" points="386" reactiontime="+78" swimtime="00:01:08.99" resultid="3855" heatid="7384" lane="4" entrytime="00:01:13.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="400" reactiontime="+81" swimtime="00:00:29.50" resultid="3856" heatid="7440" lane="5" entrytime="00:00:34.66" />
                <RESULT eventid="1481" points="421" reactiontime="+63" swimtime="00:01:05.20" resultid="3857" heatid="7466" lane="6" entrytime="00:01:06.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="410" reactiontime="+68" swimtime="00:02:22.15" resultid="3858" heatid="7535" lane="2" entrytime="00:02:26.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:45.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Samsel" nation="POL" athleteid="3859">
              <RESULTS>
                <RESULT eventid="1076" points="502" reactiontime="+71" swimtime="00:00:25.49" resultid="3860" heatid="7267" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1108" points="400" swimtime="00:02:28.74" resultid="3861" heatid="7283" lane="0" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="329" reactiontime="+71" swimtime="00:00:32.17" resultid="3862" heatid="7323" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1288" points="505" reactiontime="+70" swimtime="00:00:56.41" resultid="3863" heatid="7364" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="330" reactiontime="+74" swimtime="00:01:20.47" resultid="3864" heatid="7422" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="344" reactiontime="+68" swimtime="00:01:09.72" resultid="3865" heatid="7465" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="351" reactiontime="+70" swimtime="00:02:29.71" resultid="3866" heatid="7534" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:51.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMOLA" nation="POL" region="01" clubid="2644" name="Tri Mission Oława">
          <ATHLETES>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba-Gołaszewska" nation="POL" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1059" points="427" reactiontime="+97" swimtime="00:00:30.44" resultid="2645" heatid="7243" lane="3" entrytime="00:00:30.96" />
                <RESULT eventid="1272" points="384" reactiontime="+79" swimtime="00:01:09.10" resultid="2646" heatid="7346" lane="4" entrytime="00:01:07.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="383" reactiontime="+85" swimtime="00:00:33.56" resultid="2647" heatid="7433" lane="9" entrytime="00:00:32.78" />
                <RESULT eventid="1497" points="351" reactiontime="+88" swimtime="00:02:36.44" resultid="2648" heatid="7472" lane="2" entrytime="00:02:38.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="307" reactiontime="+83" swimtime="00:01:20.89" resultid="2649" heatid="7510" lane="3" entrytime="00:01:18.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00215" nation="POL" region="15" clubid="5660" name="TS Olimpia Poznań" shortname="Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-01" firstname="Joanna" gender="F" lastname="Bartosiewicz" nation="POL" athleteid="5670">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters kategoria G" eventid="1240" points="342" swimtime="00:03:12.31" resultid="5671" heatid="7331" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:32.70" />
                    <SPLIT distance="150" swimtime="00:02:22.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria G" eventid="1304" points="349" reactiontime="+96" swimtime="00:01:20.19" resultid="5672" heatid="7374" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="326" reactiontime="+95" swimtime="00:01:30.55" resultid="5673" heatid="7412" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="321" reactiontime="+97" swimtime="00:00:35.60" resultid="5674" heatid="7430" lane="2" entrytime="00:00:37.00" />
                <RESULT comment="Rekord Polski Masters kategoria G" eventid="1721" points="356" reactiontime="+91" swimtime="00:05:29.96" resultid="5675" heatid="7567" lane="9" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:02.79" />
                    <SPLIT distance="200" swimtime="00:02:44.66" />
                    <SPLIT distance="250" swimtime="00:03:26.48" />
                    <SPLIT distance="300" swimtime="00:04:09.15" />
                    <SPLIT distance="350" swimtime="00:04:49.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="5676">
              <RESULTS>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="5677" heatid="7299" lane="6" entrytime="00:14:50.00" />
                <RESULT eventid="1224" status="WDR" swimtime="00:00:00.00" resultid="5678" heatid="7319" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="1481" status="WDR" swimtime="00:00:00.00" resultid="5679" heatid="7461" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="1513" status="WDR" swimtime="00:00:00.00" resultid="5680" heatid="7477" lane="8" entrytime="00:03:20.00" />
                <RESULT eventid="1657" status="WDR" swimtime="00:00:00.00" resultid="5681" heatid="7531" lane="8" entrytime="00:03:44.00" />
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="5682" heatid="7584" lane="4" entrytime="00:07:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="5683">
              <RESULTS>
                <RESULT eventid="1076" points="135" swimtime="00:00:39.41" resultid="5684" heatid="7250" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1108" points="110" swimtime="00:03:48.16" resultid="5685" heatid="7278" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                    <SPLIT distance="100" swimtime="00:01:52.21" />
                    <SPLIT distance="150" swimtime="00:02:56.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria K" eventid="1224" points="112" reactiontime="+75" swimtime="00:00:46.05" resultid="5686" heatid="7318" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1320" points="115" swimtime="00:01:43.20" resultid="5687" heatid="7379" lane="0" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="74" swimtime="00:00:51.61" resultid="5688" heatid="7437" lane="9" entrytime="00:00:53.00" />
                <RESULT comment="Rekord Polski Masters kategoria K" eventid="1481" points="109" reactiontime="+88" swimtime="00:01:42.14" resultid="5689" heatid="7461" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria K" eventid="1657" points="102" reactiontime="+80" swimtime="00:03:45.88" resultid="5690" heatid="7531" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                    <SPLIT distance="100" swimtime="00:01:49.97" />
                    <SPLIT distance="150" swimtime="00:02:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="139" reactiontime="+92" swimtime="00:00:48.72" resultid="5691" heatid="7548" lane="2" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Jacek" gender="M" lastname="Matyszczak" nation="POL" athleteid="5701">
              <RESULTS>
                <RESULT eventid="1076" points="346" swimtime="00:00:28.84" resultid="5702" heatid="7260" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1156" points="242" swimtime="00:11:51.46" resultid="5703" heatid="7297" lane="9" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:02:01.61" />
                    <SPLIT distance="200" swimtime="00:02:46.89" />
                    <SPLIT distance="250" swimtime="00:03:32.20" />
                    <SPLIT distance="300" swimtime="00:04:17.62" />
                    <SPLIT distance="350" swimtime="00:05:03.88" />
                    <SPLIT distance="400" swimtime="00:05:50.27" />
                    <SPLIT distance="450" swimtime="00:06:36.95" />
                    <SPLIT distance="500" swimtime="00:07:21.82" />
                    <SPLIT distance="550" swimtime="00:08:08.08" />
                    <SPLIT distance="600" swimtime="00:08:53.47" />
                    <SPLIT distance="650" swimtime="00:09:39.51" />
                    <SPLIT distance="700" swimtime="00:10:24.34" />
                    <SPLIT distance="750" swimtime="00:11:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="199" reactiontime="+75" swimtime="00:00:38.00" resultid="5704" heatid="7320" lane="5" entrytime="00:00:38.50" />
                <RESULT eventid="1288" points="325" reactiontime="+85" swimtime="00:01:05.36" resultid="5705" heatid="7358" lane="5" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="255" reactiontime="+83" swimtime="00:00:34.29" resultid="5706" heatid="7441" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1513" points="273" reactiontime="+95" swimtime="00:02:33.02" resultid="5707" heatid="7480" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:52.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5708" heatid="7554" lane="8" entrytime="00:00:38.50" />
                <RESULT eventid="1737" points="242" reactiontime="+97" swimtime="00:05:40.22" resultid="5709" heatid="7579" lane="3" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="150" swimtime="00:01:54.68" />
                    <SPLIT distance="200" swimtime="00:02:39.13" />
                    <SPLIT distance="250" swimtime="00:03:23.93" />
                    <SPLIT distance="300" swimtime="00:04:09.91" />
                    <SPLIT distance="350" swimtime="00:04:55.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="5692">
              <RESULTS>
                <RESULT eventid="1108" points="182" reactiontime="+98" swimtime="00:03:13.17" resultid="5693" heatid="7279" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:34.47" />
                    <SPLIT distance="150" swimtime="00:02:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="197" swimtime="00:12:41.91" resultid="5694" heatid="7298" lane="5" entrytime="00:12:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:15.86" />
                    <SPLIT distance="200" swimtime="00:03:04.02" />
                    <SPLIT distance="250" swimtime="00:03:53.19" />
                    <SPLIT distance="300" swimtime="00:04:42.14" />
                    <SPLIT distance="350" swimtime="00:05:30.52" />
                    <SPLIT distance="400" swimtime="00:06:18.52" />
                    <SPLIT distance="450" swimtime="00:07:06.32" />
                    <SPLIT distance="500" swimtime="00:07:54.50" />
                    <SPLIT distance="550" swimtime="00:08:42.62" />
                    <SPLIT distance="600" swimtime="00:09:31.25" />
                    <SPLIT distance="650" swimtime="00:10:19.30" />
                    <SPLIT distance="700" swimtime="00:11:07.17" />
                    <SPLIT distance="750" swimtime="00:11:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="145" reactiontime="+92" swimtime="00:00:42.22" resultid="5695" heatid="7319" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1320" points="188" reactiontime="+94" swimtime="00:01:27.60" resultid="5696" heatid="7381" lane="9" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="168" reactiontime="+96" swimtime="00:01:28.42" resultid="5697" heatid="7462" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="200" swimtime="00:06:42.55" resultid="5698" heatid="8156" lane="7" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                    <SPLIT distance="100" swimtime="00:01:44.66" />
                    <SPLIT distance="150" swimtime="00:02:33.00" />
                    <SPLIT distance="200" swimtime="00:03:21.61" />
                    <SPLIT distance="250" swimtime="00:04:16.95" />
                    <SPLIT distance="300" swimtime="00:05:12.77" />
                    <SPLIT distance="350" swimtime="00:05:58.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="182" reactiontime="+90" swimtime="00:03:06.21" resultid="5699" heatid="7532" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="150" swimtime="00:02:19.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5700" heatid="7580" lane="8" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="5661">
              <RESULTS>
                <RESULT eventid="1059" points="168" reactiontime="+98" swimtime="00:00:41.51" resultid="5662" heatid="7237" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="1092" points="113" reactiontime="+93" swimtime="00:04:11.94" resultid="5663" heatid="7271" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.64" />
                    <SPLIT distance="100" swimtime="00:02:07.31" />
                    <SPLIT distance="150" swimtime="00:03:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="120" reactiontime="+72" swimtime="00:00:52.00" resultid="5664" heatid="7308" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1272" points="142" reactiontime="+90" swimtime="00:01:36.15" resultid="5665" heatid="7342" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="100" reactiontime="+96" swimtime="00:00:52.47" resultid="5666" heatid="7427" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="1497" points="146" reactiontime="+94" swimtime="00:03:29.66" resultid="5667" heatid="7469" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:44.57" />
                    <SPLIT distance="150" swimtime="00:02:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="75" reactiontime="+91" swimtime="00:02:09.03" resultid="5668" heatid="7507" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="145" reactiontime="+91" swimtime="00:07:25.15" resultid="5669" heatid="7570" lane="0" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:44.08" />
                    <SPLIT distance="150" swimtime="00:02:42.84" />
                    <SPLIT distance="200" swimtime="00:03:40.41" />
                    <SPLIT distance="250" swimtime="00:04:37.89" />
                    <SPLIT distance="300" swimtime="00:05:35.61" />
                    <SPLIT distance="350" swimtime="00:06:31.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" points="193" reactiontime="+82" swimtime="00:02:46.71" resultid="5710" heatid="7563" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="150" swimtime="00:02:16.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5683" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5701" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5670" number="3" />
                    <RELAYPOSITION athleteid="5661" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00413" nation="POL" region="13" clubid="4911" name="UKP Jedynka Masters Elbląg " shortname="Jedynka Masters Elbląg ">
          <CONTACT city="Elbląg" name="Wysocki" phone="696427414" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="4912">
              <RESULTS>
                <RESULT eventid="1449" points="364" reactiontime="+72" swimtime="00:00:30.44" resultid="4913" heatid="7444" lane="3" entrytime="00:00:30.33" />
                <RESULT eventid="1513" points="422" reactiontime="+72" swimtime="00:02:12.43" resultid="4914" heatid="7485" lane="7" entrytime="00:02:14.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="378" reactiontime="+76" swimtime="00:01:06.49" resultid="4915" heatid="7519" lane="4" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="392" reactiontime="+73" swimtime="00:04:49.89" resultid="4916" heatid="7574" lane="2" entrytime="00:04:44.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                    <SPLIT distance="200" swimtime="00:02:19.63" />
                    <SPLIT distance="250" swimtime="00:02:56.26" />
                    <SPLIT distance="300" swimtime="00:03:33.80" />
                    <SPLIT distance="350" swimtime="00:04:12.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-18" firstname="Maciej" gender="M" lastname="Pasieczny" nation="POL" athleteid="4917">
              <RESULTS>
                <RESULT eventid="1449" points="464" reactiontime="+75" swimtime="00:00:28.09" resultid="4918" heatid="7444" lane="5" entrytime="00:00:30.32" />
                <RESULT eventid="1513" points="443" reactiontime="+85" swimtime="00:02:10.28" resultid="4919" heatid="7485" lane="1" entrytime="00:02:14.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:02.36" />
                    <SPLIT distance="150" swimtime="00:01:36.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="6425" name="UKS Cityzen Poznań" shortname="Cityzen Poznań">
          <CONTACT city="Poznań" email="t_golembiewski@o2.pl" name="Tadeusz Gołembiewski" phone="792825485" zip="60-761" />
          <ATHLETES>
            <ATHLETE birthdate="1985-03-14" firstname="Tadeusz" gender="M" lastname="Gołembiewski" nation="POL" athleteid="6431">
              <RESULTS>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="6432" heatid="7302" lane="2" entrytime="00:19:15.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="452" reactiontime="+81" swimtime="00:00:58.52" resultid="6433" heatid="7364" lane="6" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="420" reactiontime="+82" swimtime="00:00:29.04" resultid="6434" heatid="7448" lane="3" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="442" reactiontime="+83" swimtime="00:02:10.43" resultid="6435" heatid="7487" lane="7" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:01:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="335" reactiontime="+73" swimtime="00:01:09.19" resultid="6436" heatid="7519" lane="6" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="418" reactiontime="+97" swimtime="00:04:43.74" resultid="6437" heatid="7573" lane="0" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:08.39" />
                    <SPLIT distance="150" swimtime="00:01:44.63" />
                    <SPLIT distance="200" swimtime="00:02:21.23" />
                    <SPLIT distance="250" swimtime="00:02:58.28" />
                    <SPLIT distance="300" swimtime="00:03:34.93" />
                    <SPLIT distance="350" swimtime="00:04:10.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="6444">
              <RESULTS>
                <RESULT eventid="1172" points="285" reactiontime="+98" swimtime="00:23:16.90" resultid="6445" heatid="7301" lane="4" entrytime="00:28:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:23.86" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                    <SPLIT distance="200" swimtime="00:02:56.76" />
                    <SPLIT distance="250" swimtime="00:03:44.06" />
                    <SPLIT distance="300" swimtime="00:04:31.46" />
                    <SPLIT distance="350" swimtime="00:05:18.61" />
                    <SPLIT distance="400" swimtime="00:06:05.83" />
                    <SPLIT distance="450" swimtime="00:06:52.88" />
                    <SPLIT distance="500" swimtime="00:07:40.24" />
                    <SPLIT distance="550" swimtime="00:08:27.19" />
                    <SPLIT distance="600" swimtime="00:09:14.53" />
                    <SPLIT distance="650" swimtime="00:10:01.73" />
                    <SPLIT distance="700" swimtime="00:10:48.50" />
                    <SPLIT distance="750" swimtime="00:11:35.38" />
                    <SPLIT distance="800" swimtime="00:12:22.49" />
                    <SPLIT distance="850" swimtime="00:13:10.05" />
                    <SPLIT distance="900" swimtime="00:13:56.81" />
                    <SPLIT distance="950" swimtime="00:14:43.72" />
                    <SPLIT distance="1000" swimtime="00:15:30.55" />
                    <SPLIT distance="1050" swimtime="00:16:17.29" />
                    <SPLIT distance="1100" swimtime="00:17:04.22" />
                    <SPLIT distance="1150" swimtime="00:17:51.54" />
                    <SPLIT distance="1200" swimtime="00:18:38.23" />
                    <SPLIT distance="1250" swimtime="00:19:25.21" />
                    <SPLIT distance="1300" swimtime="00:20:12.41" />
                    <SPLIT distance="1350" swimtime="00:20:59.46" />
                    <SPLIT distance="1400" swimtime="00:21:46.24" />
                    <SPLIT distance="1450" swimtime="00:22:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="253" reactiontime="+91" swimtime="00:03:32.59" resultid="6446" heatid="7329" lane="3" entrytime="00:03:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="182" reactiontime="+97" swimtime="00:03:30.84" resultid="6447" heatid="7392" lane="3" entrytime="00:03:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.51" />
                    <SPLIT distance="100" swimtime="00:01:40.31" />
                    <SPLIT distance="150" swimtime="00:02:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="230" reactiontime="+88" swimtime="00:07:02.56" resultid="6448" heatid="8150" lane="2" entrytime="00:07:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                    <SPLIT distance="150" swimtime="00:02:34.99" />
                    <SPLIT distance="200" swimtime="00:03:28.92" />
                    <SPLIT distance="250" swimtime="00:04:27.34" />
                    <SPLIT distance="300" swimtime="00:05:27.45" />
                    <SPLIT distance="350" swimtime="00:06:15.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="203" reactiontime="+91" swimtime="00:01:32.79" resultid="6449" heatid="7508" lane="4" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="271" reactiontime="+90" swimtime="00:06:01.37" resultid="6450" heatid="7568" lane="1" entrytime="00:05:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                    <SPLIT distance="200" swimtime="00:02:55.87" />
                    <SPLIT distance="250" swimtime="00:03:42.72" />
                    <SPLIT distance="300" swimtime="00:04:29.72" />
                    <SPLIT distance="350" swimtime="00:05:17.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-06" firstname="Joanna" gender="F" lastname="Krawiec" nation="POL" athleteid="6451">
              <RESULTS>
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="6452" heatid="7301" lane="5" entrytime="00:29:00.00" entrycourse="SCM" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="6453" heatid="7371" lane="5" entrytime="00:01:35.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-26" firstname="Mateusz" gender="M" lastname="Powąska" nation="POL" athleteid="6438">
              <RESULTS>
                <RESULT eventid="1076" points="443" reactiontime="+74" swimtime="00:00:26.56" resultid="6439" heatid="7261" lane="6" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="427" reactiontime="+70" swimtime="00:00:59.64" resultid="6440" heatid="7361" lane="4" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="358" reactiontime="+74" swimtime="00:01:10.75" resultid="6441" heatid="7386" lane="7" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="414" reactiontime="+70" swimtime="00:00:29.17" resultid="6442" heatid="7445" lane="3" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1689" points="318" reactiontime="+68" swimtime="00:00:36.98" resultid="6443" heatid="7553" lane="6" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-10-06" firstname="Anita" gender="F" lastname="Spendowska" nation="POL" athleteid="6458">
              <RESULTS>
                <RESULT eventid="1059" points="306" reactiontime="+87" swimtime="00:00:34.00" resultid="6459" heatid="7240" lane="2" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1272" points="263" reactiontime="+85" swimtime="00:01:18.43" resultid="6460" heatid="7343" lane="0" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="275" reactiontime="+92" swimtime="00:01:26.83" resultid="6461" heatid="7371" lane="3" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="279" reactiontime="+80" swimtime="00:00:37.30" resultid="6462" heatid="7430" lane="6" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1497" points="249" reactiontime="+83" swimtime="00:02:55.49" resultid="6463" heatid="7470" lane="8" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                    <SPLIT distance="150" swimtime="00:02:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="239" reactiontime="+86" swimtime="00:01:27.88" resultid="6464" heatid="7509" lane="0" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="263" reactiontime="+84" swimtime="00:00:44.55" resultid="6465" heatid="7540" lane="4" entrytime="00:00:46.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-14" firstname="Ewa" gender="F" lastname="Stankowska" nation="POL" athleteid="6454">
              <RESULTS>
                <RESULT eventid="1207" points="436" reactiontime="+84" swimtime="00:00:33.83" resultid="6455" heatid="7313" lane="1" entrytime="00:00:34.20" entrycourse="SCM" />
                <RESULT eventid="1304" points="377" reactiontime="+92" swimtime="00:01:18.22" resultid="6456" heatid="7374" lane="2" entrytime="00:01:17.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="425" reactiontime="+84" swimtime="00:01:13.18" resultid="6457" heatid="7457" lane="6" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-21" firstname="Tomasz" gender="M" lastname="Stankowski" nation="POL" athleteid="6426">
              <RESULTS>
                <RESULT eventid="1320" points="522" reactiontime="+77" swimtime="00:01:02.39" resultid="6427" heatid="7390" lane="0" entrytime="00:01:01.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="568" reactiontime="+62" swimtime="00:00:26.25" resultid="6428" heatid="7450" lane="2" entrytime="00:00:26.50" entrycourse="SCM" />
                <RESULT eventid="1625" points="551" reactiontime="+60" swimtime="00:00:58.62" resultid="6429" heatid="7522" lane="9" entrytime="00:00:58.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="560" reactiontime="+63" swimtime="00:00:30.62" resultid="6430" heatid="7561" lane="9" entrytime="00:00:30.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" status="DNS" swimtime="00:00:00.00" resultid="6476" heatid="7401" lane="9" entrytime="00:02:26.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6454" number="1" />
                    <RELAYPOSITION athleteid="6458" number="2" />
                    <RELAYPOSITION athleteid="6444" number="3" />
                    <RELAYPOSITION athleteid="6451" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="6477" heatid="7490" lane="4" entrytime="00:02:14.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6454" number="1" />
                    <RELAYPOSITION athleteid="6458" number="2" />
                    <RELAYPOSITION athleteid="6444" number="3" />
                    <RELAYPOSITION athleteid="6451" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1705" status="DNS" swimtime="00:00:00.00" resultid="6478" heatid="7565" lane="0" entrytime="00:02:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6454" number="1" />
                    <RELAYPOSITION athleteid="6444" number="2" />
                    <RELAYPOSITION athleteid="6426" number="3" />
                    <RELAYPOSITION athleteid="6431" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="14" clubid="3829" name="UKS Delfin Legionowo" shortname="Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="0-601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" license="101414700068" athleteid="3830">
              <RESULTS>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="3831" heatid="7561" lane="5" entrytime="00:00:28.46" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-31" firstname="Joanna" gender="F" lastname="Żbikowska" nation="POL" athleteid="3832">
              <RESULTS>
                <RESULT eventid="1059" reactiontime="+78" status="DNF" swimtime="00:00:00.00" resultid="3833" heatid="7244" lane="9" entrytime="00:00:30.69" />
                <RESULT eventid="1092" points="367" swimtime="00:02:50.15" resultid="3834" heatid="7274" lane="1" entrytime="00:02:59.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="399" reactiontime="+73" swimtime="00:03:02.67" resultid="3835" heatid="7331" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="436" reactiontime="+65" swimtime="00:01:06.23" resultid="3836" heatid="7346" lane="6" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="413" reactiontime="+74" swimtime="00:01:15.83" resultid="3837" heatid="7374" lane="5" entrytime="00:01:15.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="428" reactiontime="+76" swimtime="00:01:22.71" resultid="3838" heatid="7412" lane="4" entrytime="00:01:26.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="408" reactiontime="+67" swimtime="00:00:32.85" resultid="3839" heatid="7432" lane="6" entrytime="00:00:33.61" />
                <RESULT eventid="1497" points="398" reactiontime="+70" swimtime="00:02:30.11" resultid="3840" heatid="7473" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="431" reactiontime="+66" swimtime="00:00:37.79" resultid="3841" heatid="7545" lane="8" entrytime="00:00:36.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-23" firstname="Krzysztof" gender="M" lastname="Żbikowski" nation="POL" athleteid="3842">
              <RESULTS>
                <RESULT eventid="1108" points="411" reactiontime="+79" swimtime="00:02:27.36" resultid="3843" heatid="7285" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:01:07.76" />
                    <SPLIT distance="150" swimtime="00:01:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="461" reactiontime="+77" swimtime="00:02:35.48" resultid="3844" heatid="7339" lane="3" entrytime="00:02:30.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="489" reactiontime="+73" swimtime="00:00:57.02" resultid="3845" heatid="7364" lane="1" entrytime="00:00:58.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="510" reactiontime="+74" swimtime="00:01:02.88" resultid="3846" heatid="7390" lane="9" entrytime="00:01:02.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="603" reactiontime="+79" swimtime="00:01:05.82" resultid="3847" heatid="7425" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3848" heatid="7486" lane="0" entrytime="00:02:10.00" />
                <RESULT eventid="1689" points="618" reactiontime="+73" swimtime="00:00:29.64" resultid="3849" heatid="7561" lane="1" entrytime="00:00:29.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="08" clubid="3657" name="UKS Delfin Masters Tarnobrzeg" shortname="Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="3658">
              <RESULTS>
                <RESULT eventid="1108" points="455" swimtime="00:02:22.51" resultid="3659" heatid="7284" lane="0" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="479" reactiontime="+79" swimtime="00:02:33.55" resultid="3660" heatid="7339" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="500" reactiontime="+77" swimtime="00:01:10.06" resultid="3661" heatid="7424" lane="3" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="433" reactiontime="+82" swimtime="00:05:11.15" resultid="3662" heatid="8158" lane="1" entrytime="00:05:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:51.60" />
                    <SPLIT distance="200" swimtime="00:02:33.17" />
                    <SPLIT distance="250" swimtime="00:03:15.17" />
                    <SPLIT distance="300" swimtime="00:03:58.21" />
                    <SPLIT distance="350" swimtime="00:04:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="485" reactiontime="+71" swimtime="00:00:32.13" resultid="3663" heatid="7559" lane="6" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="3690">
              <RESULTS>
                <RESULT eventid="1059" points="363" reactiontime="+73" swimtime="00:00:32.14" resultid="3691" heatid="7243" lane="9" entrytime="00:00:31.20" />
                <RESULT eventid="1207" points="276" reactiontime="+73" swimtime="00:00:39.38" resultid="3692" heatid="7311" lane="7" entrytime="00:00:39.20" />
                <RESULT eventid="1272" points="337" reactiontime="+80" swimtime="00:01:12.14" resultid="3693" heatid="7345" lane="5" entrytime="00:01:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="276" reactiontime="+77" swimtime="00:00:37.44" resultid="3694" heatid="7429" lane="3" entrytime="00:00:38.25" />
                <RESULT eventid="1497" points="305" reactiontime="+75" swimtime="00:02:44.01" resultid="3695" heatid="7472" lane="8" entrytime="00:02:42.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="265" reactiontime="+72" swimtime="00:00:44.44" resultid="3696" heatid="7542" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="3672">
              <RESULTS>
                <RESULT eventid="1076" points="332" reactiontime="+73" swimtime="00:00:29.23" resultid="3673" heatid="7258" lane="6" entrytime="00:00:29.92" />
                <RESULT eventid="1188" points="264" reactiontime="+80" swimtime="00:22:00.99" resultid="3674" heatid="7303" lane="1" entrytime="00:22:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:19.19" />
                    <SPLIT distance="150" swimtime="00:02:02.56" />
                    <SPLIT distance="200" swimtime="00:02:46.39" />
                    <SPLIT distance="250" swimtime="00:03:30.15" />
                    <SPLIT distance="300" swimtime="00:04:14.06" />
                    <SPLIT distance="350" swimtime="00:04:58.25" />
                    <SPLIT distance="400" swimtime="00:05:42.18" />
                    <SPLIT distance="450" swimtime="00:06:26.75" />
                    <SPLIT distance="500" swimtime="00:07:11.64" />
                    <SPLIT distance="550" swimtime="00:07:56.21" />
                    <SPLIT distance="600" swimtime="00:08:41.07" />
                    <SPLIT distance="650" swimtime="00:09:25.64" />
                    <SPLIT distance="700" swimtime="00:10:10.20" />
                    <SPLIT distance="750" swimtime="00:10:54.61" />
                    <SPLIT distance="800" swimtime="00:11:39.71" />
                    <SPLIT distance="850" swimtime="00:12:24.45" />
                    <SPLIT distance="900" swimtime="00:13:08.80" />
                    <SPLIT distance="950" swimtime="00:13:53.79" />
                    <SPLIT distance="1000" swimtime="00:14:38.82" />
                    <SPLIT distance="1050" swimtime="00:15:23.14" />
                    <SPLIT distance="1100" swimtime="00:16:07.32" />
                    <SPLIT distance="1150" swimtime="00:16:52.00" />
                    <SPLIT distance="1200" swimtime="00:17:36.76" />
                    <SPLIT distance="1250" swimtime="00:18:21.25" />
                    <SPLIT distance="1300" swimtime="00:19:06.02" />
                    <SPLIT distance="1350" swimtime="00:19:50.72" />
                    <SPLIT distance="1400" swimtime="00:20:35.84" />
                    <SPLIT distance="1450" swimtime="00:21:20.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="324" reactiontime="+82" swimtime="00:01:05.39" resultid="3675" heatid="7358" lane="2" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="203" reactiontime="+78" swimtime="00:03:03.93" resultid="3676" heatid="7396" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                    <SPLIT distance="150" swimtime="00:02:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="208" reactiontime="+79" swimtime="00:01:22.44" resultid="3677" heatid="7464" lane="8" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="283" reactiontime="+74" swimtime="00:02:31.34" resultid="3678" heatid="7482" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:51.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="201" reactiontime="+84" swimtime="00:03:00.16" resultid="3679" heatid="7532" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:15.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="276" reactiontime="+73" swimtime="00:05:25.76" resultid="3680" heatid="7577" lane="9" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:57.46" />
                    <SPLIT distance="200" swimtime="00:02:39.24" />
                    <SPLIT distance="250" swimtime="00:03:21.53" />
                    <SPLIT distance="300" swimtime="00:04:04.00" />
                    <SPLIT distance="350" swimtime="00:04:46.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="3664">
              <RESULTS>
                <RESULT eventid="1092" points="304" reactiontime="+87" swimtime="00:03:01.05" resultid="3665" heatid="7274" lane="9" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                    <SPLIT distance="150" swimtime="00:02:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="278" reactiontime="+88" swimtime="00:03:25.95" resultid="3666" heatid="7330" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:38.43" />
                    <SPLIT distance="150" swimtime="00:02:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="297" reactiontime="+85" swimtime="00:01:24.63" resultid="3667" heatid="7373" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="305" reactiontime="+82" swimtime="00:01:32.59" resultid="3668" heatid="7411" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="279" reactiontime="+96" swimtime="00:06:35.84" resultid="3669" heatid="8150" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="150" swimtime="00:02:26.56" />
                    <SPLIT distance="200" swimtime="00:03:16.71" />
                    <SPLIT distance="250" swimtime="00:04:12.55" />
                    <SPLIT distance="300" swimtime="00:05:08.42" />
                    <SPLIT distance="350" swimtime="00:05:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="232" reactiontime="+88" swimtime="00:01:28.82" resultid="3670" heatid="7509" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="317" reactiontime="+80" swimtime="00:00:41.85" resultid="3671" heatid="7542" lane="3" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="3681">
              <RESULTS>
                <RESULT eventid="1076" points="447" reactiontime="+91" swimtime="00:00:26.48" resultid="3682" heatid="7257" lane="1" entrytime="00:00:30.34" />
                <RESULT eventid="1108" points="397" reactiontime="+83" swimtime="00:02:29.15" resultid="3683" heatid="7283" lane="8" entrytime="00:02:34.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:10.96" />
                    <SPLIT distance="150" swimtime="00:01:55.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="460" reactiontime="+77" swimtime="00:00:58.18" resultid="3684" heatid="7359" lane="4" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="415" reactiontime="+72" swimtime="00:01:07.35" resultid="3685" heatid="7386" lane="6" entrytime="00:01:10.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="417" reactiontime="+74" swimtime="00:01:14.43" resultid="3686" heatid="7421" lane="5" entrytime="00:01:20.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="459" reactiontime="+80" swimtime="00:02:08.75" resultid="3687" heatid="7483" lane="6" entrytime="00:02:18.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:02.53" />
                    <SPLIT distance="150" swimtime="00:01:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="375" reactiontime="+77" swimtime="00:01:06.63" resultid="3688" heatid="7518" lane="6" entrytime="00:01:10.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="427" reactiontime="+76" swimtime="00:00:33.51" resultid="3689" heatid="7557" lane="1" entrytime="00:00:35.83" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="385" reactiontime="+81" swimtime="00:02:00.81" resultid="3697" heatid="7289" lane="7" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                    <SPLIT distance="150" swimtime="00:01:27.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3681" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3658" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3690" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3664" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="364" reactiontime="+84" swimtime="00:02:14.95" resultid="3698" heatid="7565" lane="9" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:04.82" />
                    <SPLIT distance="150" swimtime="00:01:42.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3681" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3658" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3664" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="3690" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="01" clubid="2417" name="UKS Enegetyk Zgorzelec" shortname="Enegetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska" street2="2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="2418">
              <RESULTS>
                <RESULT eventid="1108" points="77" reactiontime="+87" swimtime="00:04:16.66" resultid="2419" heatid="7278" lane="7" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.69" />
                    <SPLIT distance="100" swimtime="00:02:07.16" />
                    <SPLIT distance="150" swimtime="00:03:20.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="81" reactiontime="+83" swimtime="00:17:01.23" resultid="2420" heatid="7299" lane="8" entrytime="00:17:33.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                    <SPLIT distance="100" swimtime="00:01:58.55" />
                    <SPLIT distance="150" swimtime="00:03:03.87" />
                    <SPLIT distance="200" swimtime="00:04:09.93" />
                    <SPLIT distance="250" swimtime="00:05:15.41" />
                    <SPLIT distance="300" swimtime="00:06:20.60" />
                    <SPLIT distance="350" swimtime="00:07:24.10" />
                    <SPLIT distance="400" swimtime="00:08:29.23" />
                    <SPLIT distance="450" swimtime="00:09:34.24" />
                    <SPLIT distance="500" swimtime="00:10:39.14" />
                    <SPLIT distance="550" swimtime="00:11:43.04" />
                    <SPLIT distance="600" swimtime="00:12:46.52" />
                    <SPLIT distance="650" swimtime="00:13:51.03" />
                    <SPLIT distance="700" swimtime="00:14:57.09" />
                    <SPLIT distance="750" swimtime="00:15:56.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="79" swimtime="00:04:39.79" resultid="2421" heatid="7333" lane="0" entrytime="00:04:49.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.12" />
                    <SPLIT distance="100" swimtime="00:02:16.58" />
                    <SPLIT distance="150" swimtime="00:03:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="43" reactiontime="+90" swimtime="00:05:07.09" resultid="2422" heatid="7395" lane="9" entrytime="00:04:41.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.67" />
                    <SPLIT distance="100" swimtime="00:02:24.09" />
                    <SPLIT distance="150" swimtime="00:03:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="72" swimtime="00:01:56.98" resultid="2423" heatid="7461" lane="1" entrytime="00:01:55.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="74" reactiontime="+94" swimtime="00:09:18.55" resultid="2424" heatid="8154" lane="8" entrytime="00:08:58.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.17" />
                    <SPLIT distance="100" swimtime="00:02:26.26" />
                    <SPLIT distance="150" swimtime="00:03:36.18" />
                    <SPLIT distance="200" swimtime="00:04:41.87" />
                    <SPLIT distance="250" swimtime="00:06:00.55" />
                    <SPLIT distance="300" swimtime="00:07:16.60" />
                    <SPLIT distance="350" swimtime="00:08:15.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="44" reactiontime="+86" swimtime="00:02:15.68" resultid="2425" heatid="7513" lane="5" entrytime="00:02:09.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="82" reactiontime="+93" swimtime="00:04:02.75" resultid="2426" heatid="7530" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.30" />
                    <SPLIT distance="100" swimtime="00:02:03.03" />
                    <SPLIT distance="150" swimtime="00:03:04.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00706" nation="POL" region="06" clubid="2086" name="UKS SP8 Chrzanów Chrzanów">
          <CONTACT city="CHRZANÓW" email="aba;p@poczta.onet.pl" name="ZABRZAŃSKI ALFRED" phone="692076808" state="MAŁ" street="Niepodległości 7 / 46" zip="32-500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2087">
              <RESULTS>
                <RESULT eventid="1076" points="265" reactiontime="+92" swimtime="00:00:31.54" resultid="2088" heatid="7255" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1156" points="144" reactiontime="+65" swimtime="00:14:05.25" resultid="2089" heatid="7299" lane="4" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:35.66" />
                    <SPLIT distance="150" swimtime="00:02:28.09" />
                    <SPLIT distance="200" swimtime="00:03:22.66" />
                    <SPLIT distance="250" swimtime="00:04:16.88" />
                    <SPLIT distance="300" swimtime="00:05:12.06" />
                    <SPLIT distance="350" swimtime="00:06:06.20" />
                    <SPLIT distance="400" swimtime="00:07:00.91" />
                    <SPLIT distance="450" swimtime="00:07:55.18" />
                    <SPLIT distance="500" swimtime="00:08:48.67" />
                    <SPLIT distance="550" swimtime="00:09:42.50" />
                    <SPLIT distance="600" swimtime="00:10:35.71" />
                    <SPLIT distance="650" swimtime="00:11:28.39" />
                    <SPLIT distance="700" swimtime="00:12:21.13" />
                    <SPLIT distance="750" swimtime="00:13:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="235" reactiontime="+92" swimtime="00:01:12.77" resultid="2090" heatid="7354" lane="0" entrytime="00:01:16.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2091" heatid="7380" lane="6" entrytime="00:01:29.80" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="2092" heatid="7478" lane="2" entrytime="00:02:59.03" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="2093" heatid="7582" lane="5" entrytime="00:06:39.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04814" nation="POL" region="14" clubid="3404" name="UKS Sparta Masters Grodzisk Maz." shortname="Sparta Masters Grodzisk Maz.">
          <CONTACT email="sherry@interia.pl" name="Wolnicki" phone="533544534" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-15" firstname="Dariusz" gender="M" lastname="Dziczek" nation="POL" athleteid="3428">
              <RESULTS>
                <RESULT eventid="1076" points="305" reactiontime="+89" swimtime="00:00:30.08" resultid="3429" heatid="7258" lane="1" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="348" reactiontime="+87" swimtime="00:01:03.85" resultid="3430" heatid="7358" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="301" reactiontime="+86" swimtime="00:00:32.45" resultid="3431" heatid="7441" lane="5" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="1625" points="291" reactiontime="+93" swimtime="00:01:12.51" resultid="3432" heatid="7517" lane="5" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-10-08" firstname="Michał" gender="M" lastname="Głowa" nation="POL" athleteid="3420">
              <RESULTS>
                <RESULT eventid="1288" points="318" reactiontime="+92" swimtime="00:01:05.81" resultid="3421" heatid="7359" lane="6" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="317" reactiontime="+84" swimtime="00:00:31.88" resultid="3422" heatid="7443" lane="2" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3423" heatid="7484" lane="1" entrytime="00:02:16.00" entrycourse="SCM" />
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="3424" heatid="7518" lane="5" entrytime="00:01:10.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Maciej" gender="M" lastname="Kracher" nation="POL" athleteid="3433">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3434" heatid="7258" lane="9" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3435" heatid="7358" lane="6" entrytime="00:01:06.00" entrycourse="SCM" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3436" heatid="7383" lane="3" entrytime="00:01:16.00" entrycourse="SCM" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="3437" heatid="7421" lane="7" entrytime="00:01:22.00" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3438" heatid="7482" lane="0" entrytime="00:02:30.00" entrycourse="SCM" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="3439" heatid="7556" lane="5" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-03-21" firstname="Jakub" gender="M" lastname="Stadnik" nation="POL" athleteid="3425">
              <RESULTS>
                <RESULT eventid="1288" points="273" reactiontime="+84" swimtime="00:01:09.22" resultid="3426" heatid="7354" lane="5" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="287" reactiontime="+81" swimtime="00:01:24.25" resultid="3427" heatid="7419" lane="6" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-17" firstname="Robert" gender="M" lastname="Wolnicki" nation="POL" athleteid="3410">
              <RESULTS>
                <RESULT eventid="1076" points="348" reactiontime="+95" swimtime="00:00:28.79" resultid="3411" heatid="7257" lane="6" entrytime="00:00:30.12" entrycourse="SCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="3412" heatid="7337" lane="9" entrytime="00:03:05.00" entrycourse="SCM" />
                <RESULT eventid="1417" points="362" reactiontime="+91" swimtime="00:01:17.96" resultid="3413" heatid="7421" lane="3" entrytime="00:01:20.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="384" reactiontime="+88" swimtime="00:00:34.72" resultid="3414" heatid="7556" lane="1" entrytime="00:00:36.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-18" firstname="Karol" gender="M" lastname="Zieliński" nation="POL" athleteid="3415">
              <RESULTS>
                <RESULT eventid="1256" points="295" reactiontime="+86" swimtime="00:03:00.35" resultid="3416" heatid="7335" lane="8" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:09.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="297" reactiontime="+83" swimtime="00:01:15.29" resultid="3417" heatid="7384" lane="7" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="326" reactiontime="+87" swimtime="00:01:20.75" resultid="3418" heatid="7422" lane="0" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="367" reactiontime="+79" swimtime="00:00:35.25" resultid="3419" heatid="7556" lane="6" entrytime="00:00:36.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-06-10" firstname="Ewa" gender="F" lastname="Łatkowska" nation="POL" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1172" points="145" swimtime="00:29:07.78" resultid="3406" heatid="7301" lane="3" entrytime="00:30:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                    <SPLIT distance="150" swimtime="00:02:33.16" />
                    <SPLIT distance="200" swimtime="00:03:30.66" />
                    <SPLIT distance="250" swimtime="00:04:29.15" />
                    <SPLIT distance="300" swimtime="00:05:27.97" />
                    <SPLIT distance="400" swimtime="00:07:28.54" />
                    <SPLIT distance="450" swimtime="00:08:28.51" />
                    <SPLIT distance="500" swimtime="00:09:29.19" />
                    <SPLIT distance="550" swimtime="00:10:29.79" />
                    <SPLIT distance="600" swimtime="00:11:30.33" />
                    <SPLIT distance="650" swimtime="00:12:30.71" />
                    <SPLIT distance="700" swimtime="00:13:31.55" />
                    <SPLIT distance="750" swimtime="00:14:31.80" />
                    <SPLIT distance="800" swimtime="00:15:32.16" />
                    <SPLIT distance="850" swimtime="00:16:31.79" />
                    <SPLIT distance="900" swimtime="00:17:31.55" />
                    <SPLIT distance="950" swimtime="00:18:31.45" />
                    <SPLIT distance="1000" swimtime="00:19:31.26" />
                    <SPLIT distance="1050" swimtime="00:20:29.99" />
                    <SPLIT distance="1100" swimtime="00:21:28.72" />
                    <SPLIT distance="1150" swimtime="00:22:26.89" />
                    <SPLIT distance="1200" swimtime="00:23:25.29" />
                    <SPLIT distance="1250" swimtime="00:24:23.92" />
                    <SPLIT distance="1300" swimtime="00:25:21.01" />
                    <SPLIT distance="1350" swimtime="00:26:18.92" />
                    <SPLIT distance="1400" swimtime="00:27:17.41" />
                    <SPLIT distance="1450" swimtime="00:28:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="156" swimtime="00:01:44.76" resultid="3407" heatid="7369" lane="7" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="138" swimtime="00:00:47.09" resultid="3408" heatid="7426" lane="5" entrytime="00:01:05.00" entrycourse="SCM" />
                <RESULT eventid="1721" points="147" reactiontime="+93" swimtime="00:07:23.01" resultid="3409" heatid="7571" lane="5" entrytime="00:08:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:37.86" />
                    <SPLIT distance="200" swimtime="00:03:35.69" />
                    <SPLIT distance="250" swimtime="00:04:33.64" />
                    <SPLIT distance="300" swimtime="00:05:31.66" />
                    <SPLIT distance="350" swimtime="00:06:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="357" reactiontime="+85" swimtime="00:01:55.25" resultid="3440" heatid="7494" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:00:58.41" />
                    <SPLIT distance="150" swimtime="00:01:27.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3428" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3415" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="3420" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3410" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" status="DNS" swimtime="00:00:00.00" resultid="3441" heatid="7404" lane="5" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3428" number="1" />
                    <RELAYPOSITION athleteid="3433" number="2" />
                    <RELAYPOSITION athleteid="3420" number="3" />
                    <RELAYPOSITION athleteid="3410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="11" clubid="2607" name="UKS Trójka Częstochowa" shortname="Trójka Częstochowa">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@o2.pl" name="Gawda" phone="511181791" state="ŚL" street="Schillera 5" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1995-06-07" firstname="Mateusz" gender="M" lastname="Chowaniec" nation="POL" license="100111700079" athleteid="2626">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2627" heatid="7268" lane="3" entrytime="00:00:25.34" />
                <RESULT eventid="1108" points="470" reactiontime="+76" swimtime="00:02:20.95" resultid="2628" heatid="7283" lane="5" entrytime="00:02:27.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:47.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="501" reactiontime="+73" swimtime="00:01:03.25" resultid="2629" heatid="7387" lane="2" entrytime="00:01:08.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="530" reactiontime="+77" swimtime="00:01:08.70" resultid="2630" heatid="7425" lane="9" entrytime="00:01:09.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="496" reactiontime="+75" swimtime="00:00:31.88" resultid="2631" heatid="7560" lane="6" entrytime="00:00:31.90" />
                <RESULT eventid="1737" points="422" reactiontime="+77" swimtime="00:04:42.85" resultid="2632" heatid="7576" lane="5" entrytime="00:04:55.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:42.22" />
                    <SPLIT distance="200" swimtime="00:02:18.41" />
                    <SPLIT distance="250" swimtime="00:02:54.83" />
                    <SPLIT distance="300" swimtime="00:03:31.55" />
                    <SPLIT distance="350" swimtime="00:04:08.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-04-23" firstname="Maciej" gender="M" lastname="Gajda" nation="POL" license="100111700062" athleteid="2608">
              <RESULTS>
                <RESULT eventid="1076" points="532" reactiontime="+77" swimtime="00:00:25.00" resultid="2609" heatid="7269" lane="3" entrytime="00:00:24.72" />
                <RESULT eventid="1108" points="423" reactiontime="+80" swimtime="00:02:26.01" resultid="2610" heatid="7284" lane="8" entrytime="00:02:25.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="518" reactiontime="+79" swimtime="00:00:55.95" resultid="2611" heatid="7366" lane="7" entrytime="00:00:55.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="454" reactiontime="+77" swimtime="00:01:05.36" resultid="2612" heatid="7388" lane="1" entrytime="00:01:06.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="503" reactiontime="+73" swimtime="00:00:27.34" resultid="2613" heatid="7450" lane="8" entrytime="00:00:26.92" />
                <RESULT eventid="1513" points="500" reactiontime="+75" swimtime="00:02:05.18" resultid="2614" heatid="7487" lane="6" entrytime="00:02:04.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:01:00.36" />
                    <SPLIT distance="150" swimtime="00:01:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="451" reactiontime="+78" swimtime="00:01:02.69" resultid="2615" heatid="7520" lane="6" entrytime="00:01:02.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="483" reactiontime="+81" swimtime="00:04:30.49" resultid="2616" heatid="7574" lane="3" entrytime="00:04:41.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:03.12" />
                    <SPLIT distance="150" swimtime="00:01:37.60" />
                    <SPLIT distance="200" swimtime="00:02:12.65" />
                    <SPLIT distance="250" swimtime="00:02:47.61" />
                    <SPLIT distance="300" swimtime="00:03:22.30" />
                    <SPLIT distance="350" swimtime="00:03:57.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-08-04" firstname="Wiktoria" gender="F" lastname="Musik" nation="POL" license="100111600053" athleteid="2617">
              <RESULTS>
                <RESULT eventid="1059" points="588" reactiontime="+87" swimtime="00:00:27.36" resultid="2618" heatid="7245" lane="9" entrytime="00:00:28.10" />
                <RESULT eventid="1092" points="506" reactiontime="+80" swimtime="00:02:32.88" resultid="2619" heatid="7275" lane="6" entrytime="00:02:36.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:56.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="575" reactiontime="+78" swimtime="00:01:00.40" resultid="2620" heatid="7347" lane="4" entrytime="00:01:01.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="535" reactiontime="+79" swimtime="00:01:09.61" resultid="2621" heatid="7376" lane="0" entrytime="00:01:10.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="530" reactiontime="+78" swimtime="00:00:30.12" resultid="2622" heatid="7433" lane="4" entrytime="00:00:30.63" />
                <RESULT eventid="1465" points="443" reactiontime="+77" swimtime="00:01:12.16" resultid="2623" heatid="7457" lane="3" entrytime="00:01:13.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="471" reactiontime="+78" swimtime="00:01:10.17" resultid="2624" heatid="7511" lane="1" entrytime="00:01:10.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="471" reactiontime="+76" swimtime="00:00:36.70" resultid="2625" heatid="7544" lane="8" entrytime="00:00:38.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="2876" name="UKS Trójka Puławy" shortname="Trójka Puławy">
          <CONTACT name="Gogacz" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" license="501203700057" athleteid="2877">
              <RESULTS>
                <RESULT eventid="1156" points="367" reactiontime="+90" swimtime="00:10:19.28" resultid="2878" heatid="7296" lane="6" entrytime="00:11:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="150" swimtime="00:01:50.61" />
                    <SPLIT distance="200" swimtime="00:02:29.23" />
                    <SPLIT distance="250" swimtime="00:03:08.12" />
                    <SPLIT distance="300" swimtime="00:03:46.83" />
                    <SPLIT distance="350" swimtime="00:04:25.43" />
                    <SPLIT distance="400" swimtime="00:05:04.21" />
                    <SPLIT distance="450" swimtime="00:05:43.44" />
                    <SPLIT distance="500" swimtime="00:06:22.37" />
                    <SPLIT distance="550" swimtime="00:07:01.72" />
                    <SPLIT distance="600" swimtime="00:07:41.45" />
                    <SPLIT distance="650" swimtime="00:08:21.36" />
                    <SPLIT distance="700" swimtime="00:09:01.04" />
                    <SPLIT distance="750" swimtime="00:09:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="343" reactiontime="+86" swimtime="00:02:51.65" resultid="2879" heatid="7332" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                    <SPLIT distance="150" swimtime="00:02:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="338" reactiontime="+82" swimtime="00:01:12.10" resultid="2880" heatid="7385" lane="5" entrytime="00:01:11.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="348" reactiontime="+90" swimtime="00:02:33.76" resultid="2881" heatid="7394" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:01:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="342" reactiontime="+83" swimtime="00:05:36.71" resultid="2882" heatid="8157" lane="6" entrytime="00:05:38.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:57.96" />
                    <SPLIT distance="200" swimtime="00:02:42.92" />
                    <SPLIT distance="250" swimtime="00:03:28.54" />
                    <SPLIT distance="300" swimtime="00:04:16.33" />
                    <SPLIT distance="350" swimtime="00:04:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="355" reactiontime="+79" swimtime="00:01:07.88" resultid="2883" heatid="7512" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-08" firstname="Andrzej" gender="M" lastname="Maciejczak" nation="POL" athleteid="2884">
              <RESULTS>
                <RESULT eventid="1188" points="161" reactiontime="+99" swimtime="00:25:57.27" resultid="2885" heatid="7304" lane="1" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:28.81" />
                    <SPLIT distance="150" swimtime="00:02:19.24" />
                    <SPLIT distance="200" swimtime="00:03:11.13" />
                    <SPLIT distance="250" swimtime="00:04:03.39" />
                    <SPLIT distance="300" swimtime="00:04:55.75" />
                    <SPLIT distance="350" swimtime="00:05:48.04" />
                    <SPLIT distance="400" swimtime="00:06:40.57" />
                    <SPLIT distance="450" swimtime="00:07:33.00" />
                    <SPLIT distance="500" swimtime="00:08:25.85" />
                    <SPLIT distance="550" swimtime="00:09:18.30" />
                    <SPLIT distance="600" swimtime="00:10:11.17" />
                    <SPLIT distance="650" swimtime="00:11:03.87" />
                    <SPLIT distance="700" swimtime="00:11:57.13" />
                    <SPLIT distance="750" swimtime="00:12:50.16" />
                    <SPLIT distance="800" swimtime="00:13:41.90" />
                    <SPLIT distance="850" swimtime="00:14:34.39" />
                    <SPLIT distance="900" swimtime="00:15:26.68" />
                    <SPLIT distance="950" swimtime="00:16:19.02" />
                    <SPLIT distance="1000" swimtime="00:17:11.40" />
                    <SPLIT distance="1050" swimtime="00:18:04.53" />
                    <SPLIT distance="1100" swimtime="00:18:56.88" />
                    <SPLIT distance="1150" swimtime="00:19:49.09" />
                    <SPLIT distance="1200" swimtime="00:20:42.22" />
                    <SPLIT distance="1250" swimtime="00:21:35.49" />
                    <SPLIT distance="1300" swimtime="00:22:28.90" />
                    <SPLIT distance="1350" swimtime="00:23:21.96" />
                    <SPLIT distance="1400" swimtime="00:24:15.21" />
                    <SPLIT distance="1450" swimtime="00:25:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="110" swimtime="00:08:11.48" resultid="2886" heatid="8155" lane="9" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:56.39" />
                    <SPLIT distance="150" swimtime="00:03:09.11" />
                    <SPLIT distance="200" swimtime="00:04:22.47" />
                    <SPLIT distance="250" swimtime="00:05:29.26" />
                    <SPLIT distance="300" swimtime="00:06:36.04" />
                    <SPLIT distance="350" swimtime="00:07:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="171" swimtime="00:06:21.86" resultid="2887" heatid="7582" lane="2" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:26.15" />
                    <SPLIT distance="150" swimtime="00:02:15.44" />
                    <SPLIT distance="200" swimtime="00:03:04.82" />
                    <SPLIT distance="250" swimtime="00:03:54.43" />
                    <SPLIT distance="300" swimtime="00:04:44.68" />
                    <SPLIT distance="350" swimtime="00:05:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="11" clubid="5518" name="UKS Wodnik 29 Katowice" shortname="Wodnik 29 Katowice">
          <CONTACT name="Skoczylas" />
          <ATHLETES>
            <ATHLETE birthdate="1987-04-21" firstname="Agnieszka" gender="F" lastname="Koenig" nation="POL" athleteid="5534">
              <RESULTS>
                <RESULT eventid="1207" points="56" reactiontime="+83" swimtime="00:01:06.87" resultid="5535" heatid="7307" lane="2" entrytime="00:01:08.50" />
                <RESULT eventid="1240" points="96" swimtime="00:04:53.35" resultid="5536" heatid="7327" lane="6" entrytime="00:05:15.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.69" />
                    <SPLIT distance="100" swimtime="00:02:20.74" />
                    <SPLIT distance="150" swimtime="00:03:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="90" swimtime="00:02:18.92" resultid="5537" heatid="7408" lane="2" entrytime="00:02:15.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" reactiontime="+95" status="DNF" swimtime="00:00:00.00" resultid="5538" heatid="7538" lane="9" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="5528">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5529" heatid="7256" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1256" points="291" reactiontime="+91" swimtime="00:03:01.23" resultid="5530" heatid="7337" lane="3" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                    <SPLIT distance="150" swimtime="00:02:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="283" reactiontime="+81" swimtime="00:01:16.49" resultid="5531" heatid="7383" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="324" reactiontime="+77" swimtime="00:01:20.96" resultid="5532" heatid="7422" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="342" reactiontime="+82" swimtime="00:00:36.08" resultid="5533" heatid="7557" lane="7" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-09" firstname="Edyta" gender="F" lastname="Mróz" nation="POL" athleteid="5556">
              <RESULTS>
                <RESULT eventid="1140" points="316" reactiontime="+94" swimtime="00:11:43.16" resultid="5557" heatid="7290" lane="1" entrytime="00:11:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:02:04.35" />
                    <SPLIT distance="200" swimtime="00:02:48.66" />
                    <SPLIT distance="250" swimtime="00:03:33.34" />
                    <SPLIT distance="300" swimtime="00:04:18.33" />
                    <SPLIT distance="350" swimtime="00:05:03.17" />
                    <SPLIT distance="400" swimtime="00:05:48.03" />
                    <SPLIT distance="450" swimtime="00:06:32.64" />
                    <SPLIT distance="500" swimtime="00:07:17.31" />
                    <SPLIT distance="550" swimtime="00:08:02.15" />
                    <SPLIT distance="600" swimtime="00:08:47.16" />
                    <SPLIT distance="650" swimtime="00:09:32.25" />
                    <SPLIT distance="700" swimtime="00:10:16.89" />
                    <SPLIT distance="750" swimtime="00:11:00.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="323" reactiontime="+85" swimtime="00:00:37.38" resultid="5558" heatid="7313" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1272" points="323" reactiontime="+95" swimtime="00:01:13.20" resultid="5559" heatid="7345" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="276" reactiontime="+90" swimtime="00:00:37.42" resultid="5560" heatid="7431" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1465" points="305" reactiontime="+81" swimtime="00:01:21.71" resultid="5561" heatid="7456" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="318" reactiontime="+88" swimtime="00:02:54.64" resultid="5562" heatid="7527" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:25.62" />
                    <SPLIT distance="150" swimtime="00:02:10.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="310" reactiontime="+95" swimtime="00:05:45.57" resultid="5563" heatid="7567" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:04.72" />
                    <SPLIT distance="200" swimtime="00:02:49.62" />
                    <SPLIT distance="250" swimtime="00:03:34.60" />
                    <SPLIT distance="300" swimtime="00:04:19.41" />
                    <SPLIT distance="350" swimtime="00:05:03.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="5519">
              <RESULTS>
                <RESULT eventid="1076" points="341" reactiontime="+89" swimtime="00:00:28.98" resultid="5520" heatid="7259" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1156" points="314" reactiontime="+99" swimtime="00:10:52.28" resultid="5521" heatid="7295" lane="1" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:52.46" />
                    <SPLIT distance="200" swimtime="00:02:32.82" />
                    <SPLIT distance="250" swimtime="00:03:13.87" />
                    <SPLIT distance="300" swimtime="00:03:55.00" />
                    <SPLIT distance="350" swimtime="00:04:36.37" />
                    <SPLIT distance="400" swimtime="00:05:17.97" />
                    <SPLIT distance="450" swimtime="00:05:59.68" />
                    <SPLIT distance="500" swimtime="00:06:41.58" />
                    <SPLIT distance="550" swimtime="00:07:23.70" />
                    <SPLIT distance="600" swimtime="00:08:05.47" />
                    <SPLIT distance="650" swimtime="00:08:47.68" />
                    <SPLIT distance="700" swimtime="00:09:29.81" />
                    <SPLIT distance="750" swimtime="00:10:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="359" reactiontime="+96" swimtime="00:01:03.22" resultid="5522" heatid="7359" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="224" reactiontime="+97" swimtime="00:02:58.14" resultid="5523" heatid="7396" lane="4" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:08.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="255" reactiontime="+87" swimtime="00:01:17.04" resultid="5524" heatid="7463" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5525" heatid="7482" lane="1" entrytime="00:02:30.00" />
                <RESULT eventid="1657" points="240" reactiontime="+93" swimtime="00:02:49.97" resultid="5526" heatid="7533" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:21.53" />
                    <SPLIT distance="150" swimtime="00:02:05.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="327" reactiontime="+97" swimtime="00:05:08.00" resultid="5527" heatid="7578" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:50.01" />
                    <SPLIT distance="200" swimtime="00:02:29.63" />
                    <SPLIT distance="250" swimtime="00:03:09.30" />
                    <SPLIT distance="300" swimtime="00:03:48.88" />
                    <SPLIT distance="350" swimtime="00:04:29.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-15" firstname="Jolanta" gender="F" lastname="Stefanek" nation="POL" athleteid="5547">
              <RESULTS>
                <RESULT eventid="1240" points="237" reactiontime="+76" swimtime="00:03:37.22" resultid="5548" heatid="7329" lane="2" entrytime="00:03:42.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:43.19" />
                    <SPLIT distance="150" swimtime="00:02:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="233" reactiontime="+82" swimtime="00:01:41.25" resultid="5549" heatid="7410" lane="4" entrytime="00:01:41.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="252" reactiontime="+75" swimtime="00:00:45.16" resultid="5550" heatid="7540" lane="3" entrytime="00:00:46.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="5539">
              <RESULTS>
                <RESULT eventid="1059" points="27" swimtime="00:01:15.62" resultid="5540" heatid="7234" lane="4" />
                <RESULT eventid="1140" status="DNF" swimtime="00:00:00.00" resultid="5541" heatid="7293" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.32" />
                    <SPLIT distance="100" swimtime="00:03:02.15" />
                    <SPLIT distance="150" swimtime="00:04:39.24" />
                    <SPLIT distance="200" swimtime="00:06:16.37" />
                    <SPLIT distance="250" swimtime="00:07:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="47" reactiontime="+86" swimtime="00:01:11.08" resultid="5542" heatid="7306" lane="5" />
                <RESULT eventid="1272" points="26" reactiontime="+98" swimtime="00:02:49.49" resultid="5543" heatid="7341" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="5544" heatid="7452" lane="2" />
                <RESULT eventid="1641" points="35" swimtime="00:06:01.64" resultid="5545" heatid="7524" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.60" />
                    <SPLIT distance="100" swimtime="00:03:03.56" />
                    <SPLIT distance="150" swimtime="00:04:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="5546" heatid="7572" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="5551">
              <RESULTS>
                <RESULT eventid="1076" points="298" swimtime="00:00:30.33" resultid="5552" heatid="7259" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1352" points="177" reactiontime="+95" swimtime="00:03:12.50" resultid="5553" heatid="7396" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:01:33.79" />
                    <SPLIT distance="150" swimtime="00:02:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="290" swimtime="00:00:32.83" resultid="5554" heatid="7442" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1625" points="236" reactiontime="+99" swimtime="00:01:17.73" resultid="5555" heatid="7517" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="2342" name="Unia Masters Oświęcim ">
          <ATHLETES>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" license="101006700340" athleteid="2343">
              <RESULTS>
                <RESULT eventid="1224" points="198" reactiontime="+84" swimtime="00:00:38.07" resultid="2344" heatid="7320" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1481" points="213" reactiontime="+94" swimtime="00:01:21.77" resultid="2345" heatid="7462" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="200" reactiontime="+82" swimtime="00:03:00.49" resultid="2346" heatid="7532" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:25.14" />
                    <SPLIT distance="150" swimtime="00:02:11.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-01" firstname="Barbara" gender="F" lastname="Lipniarska-Skubis" nation="POL" license="501006600377" athleteid="2347">
              <RESULTS>
                <RESULT eventid="1240" points="106" swimtime="00:04:43.47" resultid="2348" heatid="7327" lane="4" entrytime="00:04:46.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.73" />
                    <SPLIT distance="100" swimtime="00:02:18.04" />
                    <SPLIT distance="150" swimtime="00:03:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="89" swimtime="00:01:52.28" resultid="2349" heatid="7341" lane="7" entrytime="00:01:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="95" swimtime="00:02:16.52" resultid="2350" heatid="7408" lane="7" entrytime="00:02:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="84" swimtime="00:04:12.04" resultid="2351" heatid="7468" lane="3" entrytime="00:04:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                    <SPLIT distance="100" swimtime="00:01:58.85" />
                    <SPLIT distance="150" swimtime="00:03:04.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="98" swimtime="00:01:01.88" resultid="2352" heatid="7538" lane="1" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" nation="POL" license="101006600341" athleteid="2353">
              <RESULTS>
                <RESULT eventid="1207" points="312" reactiontime="+85" swimtime="00:00:37.82" resultid="2354" heatid="7310" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1465" points="285" reactiontime="+81" swimtime="00:01:23.62" resultid="2355" heatid="7455" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="279" reactiontime="+87" swimtime="00:03:02.32" resultid="2356" heatid="7526" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:02:15.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03105" nation="POL" region="05" clubid="3094" name="UTW Masters Zgierz" shortname="Masters Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ROMAN" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1997-05-30" firstname="Rzewuska" gender="F" lastname="Adrianna" nation="POL" license="503105600062" athleteid="3270">
              <RESULTS>
                <RESULT eventid="1207" points="493" reactiontime="+76" swimtime="00:00:32.48" resultid="3271" heatid="7314" lane="0" entrytime="00:00:32.30" entrycourse="SCM" />
                <RESULT eventid="1465" points="465" reactiontime="+77" swimtime="00:01:10.99" resultid="3272" heatid="7458" lane="0" entrytime="00:01:11.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="3273" heatid="7528" lane="7" entrytime="00:02:38.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-01" firstname="Justyna" gender="F" lastname="Barańska" nation="POL" license="503105600" athleteid="3274">
              <RESULTS>
                <RESULT eventid="1059" points="160" reactiontime="+98" swimtime="00:00:42.23" resultid="3275" heatid="7242" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1207" points="135" reactiontime="+86" swimtime="00:00:50.02" resultid="3276" heatid="7312" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1304" points="151" reactiontime="+98" swimtime="00:01:46.04" resultid="3277" heatid="7373" lane="7" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="165" reactiontime="+98" swimtime="00:01:53.49" resultid="3278" heatid="7412" lane="8" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-03-24" firstname="Krzysztof" gender="M" lastname="Bednarek" nation="POL" license="503105700" athleteid="3135">
              <RESULTS>
                <RESULT eventid="1076" points="175" swimtime="00:00:36.21" resultid="3136" heatid="7253" lane="4" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="168" reactiontime="+98" swimtime="00:01:21.42" resultid="3137" heatid="7354" lane="9" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="152" reactiontime="+95" swimtime="00:03:06.00" resultid="3138" heatid="7477" lane="1" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                    <SPLIT distance="150" swimtime="00:02:17.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="151" swimtime="00:06:38.23" resultid="3139" heatid="7582" lane="0" entrytime="00:07:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:17.30" />
                    <SPLIT distance="200" swimtime="00:03:08.38" />
                    <SPLIT distance="250" swimtime="00:04:01.15" />
                    <SPLIT distance="300" swimtime="00:04:53.90" />
                    <SPLIT distance="350" swimtime="00:05:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-12-27" firstname="Sławomir" gender="M" lastname="Bielawski" nation="POL" license="503105700" athleteid="3140">
              <RESULTS>
                <RESULT eventid="1076" points="183" reactiontime="+93" swimtime="00:00:35.67" resultid="3141" heatid="7251" lane="7" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1449" points="144" reactiontime="+96" swimtime="00:00:41.48" resultid="3142" heatid="7437" lane="5" entrytime="00:00:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="3238">
              <RESULTS>
                <RESULT eventid="1076" points="116" reactiontime="+99" swimtime="00:00:41.51" resultid="3239" heatid="7249" lane="2" entrytime="00:00:40.91" entrycourse="SCM" />
                <RESULT eventid="1108" points="75" swimtime="00:04:19.27" resultid="3240" heatid="7278" lane="0" entrytime="00:04:18.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.55" />
                    <SPLIT distance="100" swimtime="00:02:05.55" />
                    <SPLIT distance="150" swimtime="00:03:24.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="101" reactiontime="+83" swimtime="00:01:36.31" resultid="3241" heatid="7351" lane="7" entrytime="00:01:36.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="36" reactiontime="+86" swimtime="00:05:26.88" resultid="3242" heatid="7394" lane="6" entrytime="00:05:08.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.68" />
                    <SPLIT distance="100" swimtime="00:02:36.36" />
                    <SPLIT distance="150" swimtime="00:04:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="106" reactiontime="+82" swimtime="00:03:29.37" resultid="3243" heatid="7476" lane="6" entrytime="00:03:42.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="150" swimtime="00:02:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="66" reactiontime="+92" swimtime="00:09:39.93" resultid="3244" heatid="8154" lane="0" entrytime="00:09:16.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.41" />
                    <SPLIT distance="100" swimtime="00:02:43.08" />
                    <SPLIT distance="150" swimtime="00:03:57.19" />
                    <SPLIT distance="200" swimtime="00:05:07.66" />
                    <SPLIT distance="250" swimtime="00:06:28.72" />
                    <SPLIT distance="300" swimtime="00:07:50.99" />
                    <SPLIT distance="350" swimtime="00:08:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="33" reactiontime="+92" swimtime="00:02:28.95" resultid="3245" heatid="7513" lane="0" entrytime="00:02:19.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="59" reactiontime="+97" swimtime="00:04:30.37" resultid="3246" heatid="7530" lane="8" entrytime="00:04:30.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.77" />
                    <SPLIT distance="150" swimtime="00:03:25.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105700035" athleteid="3288">
              <RESULTS>
                <RESULT eventid="1076" points="211" reactiontime="+85" swimtime="00:00:34.00" resultid="3289" heatid="7254" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1417" points="148" reactiontime="+90" swimtime="00:01:45.06" resultid="3290" heatid="7418" lane="8" entrytime="00:01:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="180" swimtime="00:00:44.72" resultid="3291" heatid="7550" lane="6" entrytime="00:00:43.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-09" firstname="Łukasz" gender="M" lastname="Chwiałkowski" nation="POL" license="503105700057" athleteid="3263">
              <RESULTS>
                <RESULT eventid="1076" points="284" reactiontime="+92" swimtime="00:00:30.82" resultid="3264" heatid="7251" lane="5" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1156" points="245" reactiontime="+96" swimtime="00:11:48.56" resultid="3265" heatid="7296" lane="3" entrytime="00:11:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                    <SPLIT distance="200" swimtime="00:02:42.03" />
                    <SPLIT distance="250" swimtime="00:03:25.49" />
                    <SPLIT distance="300" swimtime="00:04:09.14" />
                    <SPLIT distance="350" swimtime="00:04:54.29" />
                    <SPLIT distance="400" swimtime="00:05:40.09" />
                    <SPLIT distance="450" swimtime="00:06:25.50" />
                    <SPLIT distance="500" swimtime="00:07:11.03" />
                    <SPLIT distance="550" swimtime="00:07:57.45" />
                    <SPLIT distance="600" swimtime="00:08:43.83" />
                    <SPLIT distance="650" swimtime="00:09:30.17" />
                    <SPLIT distance="700" swimtime="00:10:17.32" />
                    <SPLIT distance="750" swimtime="00:11:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="3266" heatid="7320" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3267" heatid="7353" lane="0" entrytime="00:01:21.00" entrycourse="SCM" />
                <RESULT eventid="1513" points="262" reactiontime="+94" swimtime="00:02:35.14" resultid="3268" heatid="7479" lane="8" entrytime="00:02:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="220" reactiontime="+97" swimtime="00:05:51.15" resultid="3269" heatid="7580" lane="2" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                    <SPLIT distance="200" swimtime="00:02:43.36" />
                    <SPLIT distance="250" swimtime="00:03:27.48" />
                    <SPLIT distance="300" swimtime="00:04:11.46" />
                    <SPLIT distance="350" swimtime="00:04:54.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-02-19" firstname="Jacek" gender="M" lastname="Dziarek" nation="POL" license="503105700061" athleteid="3257">
              <RESULTS>
                <RESULT eventid="1076" points="261" swimtime="00:00:31.68" resultid="3258" heatid="7255" lane="5" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1188" points="226" swimtime="00:23:10.26" resultid="3259" heatid="7304" lane="5" entrytime="00:24:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:23.79" />
                    <SPLIT distance="150" swimtime="00:02:08.42" />
                    <SPLIT distance="200" swimtime="00:02:53.63" />
                    <SPLIT distance="250" swimtime="00:03:39.22" />
                    <SPLIT distance="300" swimtime="00:04:24.21" />
                    <SPLIT distance="350" swimtime="00:05:10.03" />
                    <SPLIT distance="400" swimtime="00:05:55.88" />
                    <SPLIT distance="450" swimtime="00:06:41.86" />
                    <SPLIT distance="500" swimtime="00:07:27.86" />
                    <SPLIT distance="550" swimtime="00:08:13.41" />
                    <SPLIT distance="600" swimtime="00:08:58.99" />
                    <SPLIT distance="650" swimtime="00:09:45.20" />
                    <SPLIT distance="700" swimtime="00:10:31.43" />
                    <SPLIT distance="750" swimtime="00:11:18.43" />
                    <SPLIT distance="800" swimtime="00:12:05.32" />
                    <SPLIT distance="900" swimtime="00:13:40.53" />
                    <SPLIT distance="950" swimtime="00:14:27.99" />
                    <SPLIT distance="1050" swimtime="00:16:02.88" />
                    <SPLIT distance="1100" swimtime="00:16:51.15" />
                    <SPLIT distance="1150" swimtime="00:17:38.75" />
                    <SPLIT distance="1200" swimtime="00:18:25.95" />
                    <SPLIT distance="1250" swimtime="00:19:13.16" />
                    <SPLIT distance="1300" swimtime="00:20:01.44" />
                    <SPLIT distance="1350" swimtime="00:20:49.33" />
                    <SPLIT distance="1400" swimtime="00:21:36.71" />
                    <SPLIT distance="1450" swimtime="00:22:24.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="261" reactiontime="+98" swimtime="00:01:10.24" resultid="3260" heatid="7355" lane="3" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="231" swimtime="00:02:41.83" resultid="3261" heatid="7479" lane="4" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="228" swimtime="00:05:47.23" resultid="3262" heatid="7579" lane="9" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                    <SPLIT distance="200" swimtime="00:02:52.89" />
                    <SPLIT distance="250" swimtime="00:03:37.07" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:05:05.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="3153">
              <RESULTS>
                <RESULT eventid="1059" points="498" reactiontime="+90" swimtime="00:00:28.92" resultid="3154" heatid="7244" lane="1" entrytime="00:00:29.90" entrycourse="SCM" />
                <RESULT eventid="1207" points="505" reactiontime="+83" swimtime="00:00:32.23" resultid="3155" heatid="7313" lane="6" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1304" points="481" reactiontime="+82" swimtime="00:01:12.11" resultid="3156" heatid="7375" lane="6" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="468" reactiontime="+76" swimtime="00:01:10.86" resultid="3157" heatid="7458" lane="9" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="426" reactiontime="+89" swimtime="00:05:44.04" resultid="3158" heatid="8151" lane="8" entrytime="00:06:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                    <SPLIT distance="200" swimtime="00:02:44.20" />
                    <SPLIT distance="250" swimtime="00:03:33.68" />
                    <SPLIT distance="300" swimtime="00:04:23.15" />
                    <SPLIT distance="350" swimtime="00:05:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="436" reactiontime="+79" swimtime="00:02:37.23" resultid="3159" heatid="7527" lane="4" entrytime="00:02:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-08-03" firstname="Katarzyna" gender="F" lastname="Izert" nation="POL" license="503105600" athleteid="3292">
              <RESULTS>
                <RESULT eventid="1059" points="278" reactiontime="+85" swimtime="00:00:35.10" resultid="3293" heatid="7240" lane="8" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1207" points="187" swimtime="00:00:44.87" resultid="3294" heatid="7306" lane="4" />
                <RESULT eventid="1272" points="247" reactiontime="+77" swimtime="00:01:20.03" resultid="3295" heatid="7344" lane="6" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" status="DNS" swimtime="00:00:00.00" resultid="3296" heatid="7452" lane="0" />
                <RESULT eventid="1497" points="202" reactiontime="+93" swimtime="00:03:08.00" resultid="3297" heatid="7471" lane="9" entrytime="00:02:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:25.22" />
                    <SPLIT distance="150" swimtime="00:02:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="188" reactiontime="+84" swimtime="00:00:49.81" resultid="3298" heatid="7537" lane="8" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="3299" heatid="7569" lane="5" entrytime="00:06:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="3198">
              <RESULTS>
                <RESULT eventid="1076" points="498" reactiontime="+82" swimtime="00:00:25.56" resultid="3199" heatid="7267" lane="9" entrytime="00:00:26.20" entrycourse="SCM" />
                <RESULT eventid="1108" points="426" reactiontime="+88" swimtime="00:02:25.64" resultid="3200" heatid="7283" lane="3" entrytime="00:02:27.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="414" reactiontime="+95" swimtime="00:02:41.16" resultid="3201" heatid="7339" lane="0" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="478" reactiontime="+86" swimtime="00:01:04.24" resultid="3202" heatid="7388" lane="5" entrytime="00:01:05.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="492" reactiontime="+88" swimtime="00:01:10.44" resultid="3203" heatid="7424" lane="4" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="443" reactiontime="+88" swimtime="00:02:10.35" resultid="3204" heatid="7484" lane="4" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:01:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" status="DNS" swimtime="00:00:00.00" resultid="3205" heatid="7517" lane="1" entrytime="00:01:07.00" entrycourse="SCM" />
                <RESULT eventid="1689" points="489" reactiontime="+71" swimtime="00:00:32.03" resultid="3206" heatid="7560" lane="9" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-23" firstname="Zdzisław" gender="M" lastname="Jasiński" nation="POL" license="503105700064" athleteid="3117">
              <RESULTS>
                <RESULT eventid="1076" points="190" swimtime="00:00:35.22" resultid="3118" heatid="7253" lane="6" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="192" reactiontime="+76" swimtime="00:01:17.84" resultid="3119" heatid="7353" lane="2" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="152" swimtime="00:01:34.04" resultid="3120" heatid="7380" lane="0" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="131" reactiontime="+90" swimtime="00:00:42.74" resultid="3121" heatid="7438" lane="8" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3122" heatid="7478" lane="1" entrytime="00:03:00.00" entrycourse="SCM" />
                <RESULT eventid="1689" points="153" reactiontime="+91" swimtime="00:00:47.12" resultid="3123" heatid="7552" lane="9" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-08" firstname="Piotr" gender="M" lastname="Kapczyński" nation="POL" license="503105700043" athleteid="3219">
              <RESULTS>
                <RESULT eventid="1076" points="292" reactiontime="+80" swimtime="00:00:30.53" resultid="3220" heatid="7259" lane="4" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1256" points="238" reactiontime="+82" swimtime="00:03:13.86" resultid="3221" heatid="7336" lane="9" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:33.64" />
                    <SPLIT distance="150" swimtime="00:02:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="284" reactiontime="+73" swimtime="00:01:24.58" resultid="3222" heatid="7420" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="302" reactiontime="+92" swimtime="00:00:37.63" resultid="3223" heatid="7556" lane="8" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-25" firstname="Joanna" gender="F" lastname="Kańska-Papiernik" nation="POL" license="503105600058" athleteid="3172">
              <RESULTS>
                <RESULT eventid="1059" points="411" reactiontime="+85" swimtime="00:00:30.84" resultid="3173" heatid="7243" lane="8" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1207" points="371" reactiontime="+82" swimtime="00:00:35.71" resultid="3174" heatid="7312" lane="3" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1400" points="393" reactiontime="+78" swimtime="00:01:25.07" resultid="3175" heatid="7412" lane="5" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="344" reactiontime="+75" swimtime="00:01:18.52" resultid="3176" heatid="7457" lane="9" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="324" reactiontime="+71" swimtime="00:02:53.42" resultid="3177" heatid="7527" lane="7" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="410" reactiontime="+72" swimtime="00:00:38.42" resultid="3178" heatid="7544" lane="7" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Maja" gender="F" lastname="Klusek" nation="POL" license="503105600059" athleteid="3166">
              <RESULTS>
                <RESULT eventid="1092" points="315" reactiontime="+96" swimtime="00:02:58.91" resultid="3167" heatid="7273" lane="5" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="282" swimtime="00:03:02.37" resultid="3168" heatid="7393" lane="7" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="310" reactiontime="+93" swimtime="00:00:36.02" resultid="3169" heatid="7431" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1561" points="328" swimtime="00:06:15.37" resultid="3170" heatid="8151" lane="1" entrytime="00:06:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                    <SPLIT distance="250" swimtime="00:03:55.68" />
                    <SPLIT distance="300" swimtime="00:04:49.08" />
                    <SPLIT distance="350" swimtime="00:05:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="324" reactiontime="+92" swimtime="00:01:19.47" resultid="3171" heatid="7510" lane="7" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="3124">
              <RESULTS>
                <RESULT eventid="1076" points="199" swimtime="00:00:34.67" resultid="3125" heatid="7252" lane="0" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1108" points="106" reactiontime="+91" swimtime="00:03:51.03" resultid="3126" heatid="7278" lane="6" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.27" />
                    <SPLIT distance="100" swimtime="00:01:56.04" />
                    <SPLIT distance="150" swimtime="00:03:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="127" reactiontime="+84" swimtime="00:01:39.77" resultid="3127" heatid="7379" lane="2" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="147" reactiontime="+80" swimtime="00:00:41.19" resultid="3128" heatid="7438" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1625" points="80" swimtime="00:01:51.39" resultid="3129" heatid="7514" lane="0" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="Maciejewski" nation="POL" license="503105700063" athleteid="3130">
              <RESULTS>
                <RESULT eventid="1076" points="274" reactiontime="+87" swimtime="00:00:31.17" resultid="3131" heatid="7254" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="272" reactiontime="+89" swimtime="00:01:09.30" resultid="3132" heatid="7356" lane="4" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="259" reactiontime="+90" swimtime="00:01:27.18" resultid="3133" heatid="7419" lane="9" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="262" reactiontime="+93" swimtime="00:00:39.45" resultid="3134" heatid="7553" lane="9" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="3102">
              <RESULTS>
                <RESULT eventid="1059" points="338" reactiontime="+87" swimtime="00:00:32.91" resultid="3103" heatid="7242" lane="5" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1207" points="279" reactiontime="+79" swimtime="00:00:39.27" resultid="3104" heatid="7312" lane="1" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1304" points="322" reactiontime="+88" swimtime="00:01:22.41" resultid="3105" heatid="7372" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="348" reactiontime="+91" swimtime="00:00:34.65" resultid="3106" heatid="7431" lane="2" entrytime="00:00:35.30" entrycourse="SCM" />
                <RESULT eventid="1465" points="259" reactiontime="+81" swimtime="00:01:26.23" resultid="3107" heatid="7456" lane="8" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="3108" heatid="7510" lane="0" entrytime="00:01:25.00" entrycourse="SCM" />
                <RESULT eventid="1641" points="239" reactiontime="+80" swimtime="00:03:12.06" resultid="3109" heatid="7526" lane="4" entrytime="00:03:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                    <SPLIT distance="100" swimtime="00:01:32.44" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-07-18" firstname="Tomasz" gender="M" lastname="Niedźwiedź" nation="POL" license="503105700031" athleteid="3279">
              <RESULTS>
                <RESULT eventid="1352" points="88" swimtime="00:04:03.00" resultid="3280" heatid="7395" lane="3" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:55.83" />
                    <SPLIT distance="150" swimtime="00:03:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" status="DNS" swimtime="00:00:00.00" resultid="3281" heatid="8155" lane="1" entrytime="00:07:40.00" entrycourse="SCM" />
                <RESULT eventid="1657" points="102" reactiontime="+97" swimtime="00:03:45.39" resultid="3282" heatid="7530" lane="6" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.14" />
                    <SPLIT distance="100" swimtime="00:01:50.09" />
                    <SPLIT distance="150" swimtime="00:02:47.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="3143">
              <RESULTS>
                <RESULT eventid="1256" status="WDR" swimtime="00:00:00.00" resultid="3144" heatid="7334" lane="7" entrytime="00:03:48.00" entrycourse="SCM" />
                <RESULT eventid="1417" status="WDR" swimtime="00:00:00.00" resultid="3145" heatid="7415" lane="5" entrytime="00:01:37.00" entrycourse="SCM" />
                <RESULT eventid="1689" status="WDR" swimtime="00:00:00.00" resultid="3146" heatid="7550" lane="4" entrytime="00:00:42.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-12-01" firstname="Sergiusz" gender="M" lastname="Olejniczak" nation="POL" license="503105700" athleteid="3232">
              <RESULTS>
                <RESULT eventid="1188" points="373" reactiontime="+80" swimtime="00:19:37.96" resultid="3233" heatid="7303" lane="8" entrytime="00:22:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                    <SPLIT distance="200" swimtime="00:02:28.77" />
                    <SPLIT distance="250" swimtime="00:03:07.19" />
                    <SPLIT distance="300" swimtime="00:03:45.69" />
                    <SPLIT distance="350" swimtime="00:04:24.36" />
                    <SPLIT distance="400" swimtime="00:05:03.29" />
                    <SPLIT distance="450" swimtime="00:05:42.23" />
                    <SPLIT distance="500" swimtime="00:06:21.61" />
                    <SPLIT distance="550" swimtime="00:07:01.23" />
                    <SPLIT distance="600" swimtime="00:07:40.52" />
                    <SPLIT distance="650" swimtime="00:08:19.71" />
                    <SPLIT distance="700" swimtime="00:08:59.25" />
                    <SPLIT distance="750" swimtime="00:09:39.00" />
                    <SPLIT distance="800" swimtime="00:10:18.40" />
                    <SPLIT distance="850" swimtime="00:10:57.64" />
                    <SPLIT distance="900" swimtime="00:11:36.97" />
                    <SPLIT distance="950" swimtime="00:12:16.71" />
                    <SPLIT distance="1000" swimtime="00:12:56.86" />
                    <SPLIT distance="1050" swimtime="00:13:36.19" />
                    <SPLIT distance="1100" swimtime="00:14:16.61" />
                    <SPLIT distance="1150" swimtime="00:14:55.93" />
                    <SPLIT distance="1200" swimtime="00:15:35.75" />
                    <SPLIT distance="1250" swimtime="00:16:15.88" />
                    <SPLIT distance="1300" swimtime="00:16:56.23" />
                    <SPLIT distance="1350" swimtime="00:17:36.65" />
                    <SPLIT distance="1400" swimtime="00:18:17.60" />
                    <SPLIT distance="1450" swimtime="00:18:58.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="369" reactiontime="+73" swimtime="00:02:47.47" resultid="3234" heatid="7339" lane="8" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="296" reactiontime="+75" swimtime="00:02:42.36" resultid="3235" heatid="7397" lane="4" entrytime="00:02:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:02:01.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="373" reactiontime="+73" swimtime="00:05:27.14" resultid="3236" heatid="8157" lane="0" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:01:59.88" />
                    <SPLIT distance="200" swimtime="00:02:39.98" />
                    <SPLIT distance="250" swimtime="00:03:24.86" />
                    <SPLIT distance="300" swimtime="00:04:11.26" />
                    <SPLIT distance="350" swimtime="00:04:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="368" reactiontime="+69" swimtime="00:04:56.01" resultid="3237" heatid="7578" lane="1" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:47.26" />
                    <SPLIT distance="200" swimtime="00:02:25.15" />
                    <SPLIT distance="250" swimtime="00:03:03.46" />
                    <SPLIT distance="300" swimtime="00:03:41.73" />
                    <SPLIT distance="350" swimtime="00:04:19.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-11-22" firstname="Jakub" gender="M" lastname="Papiernik" nation="POL" license="503105700" athleteid="3252">
              <RESULTS>
                <RESULT eventid="1076" points="299" reactiontime="+80" swimtime="00:00:30.29" resultid="3253" heatid="7257" lane="9" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1320" points="290" reactiontime="+80" swimtime="00:01:15.87" resultid="3254" heatid="7382" lane="7" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="222" reactiontime="+82" swimtime="00:02:44.03" resultid="3255" heatid="7479" lane="6" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="274" reactiontime="+79" swimtime="00:00:38.87" resultid="3256" heatid="7554" lane="7" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="3210">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="3211" heatid="7280" lane="2" entrytime="00:03:05.00" entrycourse="SCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="3212" heatid="7297" lane="6" entrytime="00:12:00.00" entrycourse="SCM" />
                <RESULT eventid="1224" points="234" reactiontime="+75" swimtime="00:00:36.05" resultid="3213" heatid="7321" lane="8" entrytime="00:00:37.50" entrycourse="SCM" />
                <RESULT eventid="1288" points="284" reactiontime="+88" swimtime="00:01:08.29" resultid="3214" heatid="7357" lane="9" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="204" reactiontime="+91" swimtime="00:01:22.91" resultid="3215" heatid="7463" lane="1" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="3216" heatid="7480" lane="9" entrytime="00:02:40.00" entrycourse="SCM" />
                <RESULT eventid="1657" points="190" reactiontime="+81" swimtime="00:03:03.68" resultid="3217" heatid="7532" lane="4" entrytime="00:03:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="3218" heatid="7579" lane="1" entrytime="00:05:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-03" firstname="Stanisław" gender="M" lastname="Sikorski" nation="POL" license="503105700054" athleteid="3247">
              <RESULTS>
                <RESULT eventid="1224" points="57" reactiontime="+93" swimtime="00:00:57.60" resultid="3248" heatid="7318" lane="8" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1417" points="98" swimtime="00:02:00.45" resultid="3249" heatid="7415" lane="4" entrytime="00:02:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="45" swimtime="00:02:16.51" resultid="3250" heatid="7460" lane="5" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="118" swimtime="00:00:51.39" resultid="3251" heatid="7548" lane="3" entrytime="00:00:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="3224">
              <RESULTS>
                <RESULT eventid="1108" points="519" reactiontime="+82" swimtime="00:02:16.34" resultid="3225" heatid="7284" lane="6" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:01:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="545" reactiontime="+75" swimtime="00:00:55.00" resultid="3226" heatid="7363" lane="6" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="580" reactiontime="+77" swimtime="00:01:00.26" resultid="3227" heatid="7388" lane="9" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="595" reactiontime="+84" swimtime="00:01:06.10" resultid="3228" heatid="7425" lane="0" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="543" reactiontime="+80" swimtime="00:00:26.65" resultid="3229" heatid="7448" lane="0" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1625" points="565" reactiontime="+80" swimtime="00:00:58.13" resultid="3230" heatid="7519" lane="3" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="593" reactiontime="+71" swimtime="00:00:30.04" resultid="3231" heatid="7560" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" license="503105700060" athleteid="3183">
              <RESULTS>
                <RESULT eventid="1076" points="261" reactiontime="+82" swimtime="00:00:31.70" resultid="3184" heatid="7256" lane="1" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="1108" points="222" reactiontime="+82" swimtime="00:03:00.81" resultid="3185" heatid="7280" lane="6" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="150" swimtime="00:02:15.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="218" reactiontime="+79" swimtime="00:03:19.47" resultid="3186" heatid="7335" lane="9" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="150" swimtime="00:02:26.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="250" reactiontime="+81" swimtime="00:01:19.69" resultid="3187" heatid="7381" lane="1" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="240" reactiontime="+80" swimtime="00:01:29.46" resultid="3188" heatid="7419" lane="7" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="171" reactiontime="+69" swimtime="00:07:03.64" resultid="3189" heatid="8155" lane="4" entrytime="00:07:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:42.85" />
                    <SPLIT distance="150" swimtime="00:02:37.23" />
                    <SPLIT distance="200" swimtime="00:03:31.80" />
                    <SPLIT distance="250" swimtime="00:04:29.38" />
                    <SPLIT distance="300" swimtime="00:05:26.58" />
                    <SPLIT distance="350" swimtime="00:06:15.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="167" reactiontime="+79" swimtime="00:01:27.26" resultid="3190" heatid="7515" lane="4" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="264" reactiontime="+69" swimtime="00:00:39.36" resultid="3191" heatid="7552" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-06" firstname="Robert" gender="M" lastname="Szalbierz" nation="POL" license="503105700056" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1076" points="286" reactiontime="+92" swimtime="00:00:30.74" resultid="3180" heatid="7257" lane="5" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3181" heatid="7381" lane="4" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="1449" points="279" reactiontime="+94" swimtime="00:00:33.27" resultid="3182" heatid="7442" lane="9" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="Szcęsnowicz" nation="POL" license="503105600052" athleteid="3110">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3111" heatid="7244" lane="8" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1207" status="WDR" swimtime="00:00:00.00" resultid="3112" heatid="7310" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1304" status="WDR" swimtime="00:00:00.00" resultid="3113" heatid="7372" lane="1" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1400" status="WDR" swimtime="00:00:00.00" resultid="3114" heatid="7412" lane="2" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1433" status="WDR" swimtime="00:00:00.00" resultid="3115" heatid="7432" lane="0" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1673" status="WDR" swimtime="00:00:00.00" resultid="3116" heatid="7544" lane="1" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-06" firstname="Wojciech" gender="M" lastname="Szymański" nation="POL" license="503105700037" athleteid="3207">
              <RESULTS>
                <RESULT eventid="1224" points="62" reactiontime="+79" swimtime="00:00:55.94" resultid="3208" heatid="7318" lane="0" entrytime="00:00:51.00" entrycourse="SCM" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="3209" heatid="7460" lane="6" entrytime="00:02:06.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700032" athleteid="3095">
              <RESULTS>
                <RESULT eventid="1156" points="124" reactiontime="+70" swimtime="00:14:48.96" resultid="3096" heatid="7299" lane="2" entrytime="00:15:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:42.93" />
                    <SPLIT distance="150" swimtime="00:02:39.42" />
                    <SPLIT distance="200" swimtime="00:03:35.43" />
                    <SPLIT distance="250" swimtime="00:04:30.97" />
                    <SPLIT distance="300" swimtime="00:05:26.48" />
                    <SPLIT distance="350" swimtime="00:06:21.48" />
                    <SPLIT distance="400" swimtime="00:07:17.44" />
                    <SPLIT distance="450" swimtime="00:08:13.50" />
                    <SPLIT distance="500" swimtime="00:09:09.21" />
                    <SPLIT distance="550" swimtime="00:10:07.53" />
                    <SPLIT distance="600" swimtime="00:11:05.84" />
                    <SPLIT distance="650" swimtime="00:12:02.49" />
                    <SPLIT distance="700" swimtime="00:13:01.02" />
                    <SPLIT distance="750" swimtime="00:13:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="172" swimtime="00:03:35.80" resultid="3097" heatid="7334" lane="4" entrytime="00:03:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                    <SPLIT distance="100" swimtime="00:01:44.19" />
                    <SPLIT distance="150" swimtime="00:02:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="181" reactiontime="+94" swimtime="00:01:38.25" resultid="3098" heatid="7419" lane="0" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="120" reactiontime="+83" swimtime="00:01:38.85" resultid="3099" heatid="7462" lane="7" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="120" reactiontime="+81" swimtime="00:03:34.09" resultid="3100" heatid="7531" lane="6" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                    <SPLIT distance="100" swimtime="00:01:44.14" />
                    <SPLIT distance="150" swimtime="00:02:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="200" reactiontime="+99" swimtime="00:00:43.16" resultid="3101" heatid="7551" lane="8" entrytime="00:00:42.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Woźniak" nation="POL" license="503105700039" athleteid="3192">
              <RESULTS>
                <RESULT eventid="1224" points="442" reactiontime="+51" swimtime="00:00:29.16" resultid="3193" heatid="7326" lane="9" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1449" points="452" reactiontime="+80" swimtime="00:00:28.32" resultid="3194" heatid="7436" lane="7" entrytime="00:02:00.00" entrycourse="SCM" />
                <RESULT eventid="1481" points="455" reactiontime="+55" swimtime="00:01:03.51" resultid="3195" heatid="7466" lane="3" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="420" reactiontime="+84" swimtime="00:01:04.16" resultid="3196" heatid="7512" lane="3" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="419" reactiontime="+56" swimtime="00:02:21.07" resultid="3197" heatid="7535" lane="5" entrytime="00:02:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                    <SPLIT distance="150" swimtime="00:01:46.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-26" firstname="Katarzyna" gender="F" lastname="Węgrzycka" nation="POL" license="503105600" athleteid="3300">
              <RESULTS>
                <RESULT eventid="1059" points="88" swimtime="00:00:51.51" resultid="3301" heatid="7240" lane="6" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1400" points="119" swimtime="00:02:06.53" resultid="3302" heatid="7411" lane="7" entrytime="00:01:38.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="407" swimtime="00:00:38.51" resultid="3303" heatid="7543" lane="9" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-08" firstname="Ewa" gender="F" lastname="Zimna-Walendzik" nation="POL" license="503105600019" athleteid="3283">
              <RESULTS>
                <RESULT eventid="1092" points="123" swimtime="00:04:04.39" resultid="3284" heatid="7271" lane="2" entrytime="00:04:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                    <SPLIT distance="100" swimtime="00:01:57.89" />
                    <SPLIT distance="150" swimtime="00:03:08.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="118" swimtime="00:08:47.72" resultid="3285" heatid="8149" lane="1" entrytime="00:08:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                    <SPLIT distance="100" swimtime="00:02:05.81" />
                    <SPLIT distance="150" swimtime="00:03:15.37" />
                    <SPLIT distance="200" swimtime="00:04:23.58" />
                    <SPLIT distance="250" swimtime="00:05:34.11" />
                    <SPLIT distance="300" swimtime="00:06:47.91" />
                    <SPLIT distance="350" swimtime="00:07:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="3286" heatid="7508" lane="9" entrytime="00:02:09.00" entrycourse="SCM" />
                <RESULT eventid="1721" points="128" reactiontime="+99" swimtime="00:07:43.13" resultid="3287" heatid="7571" lane="4" entrytime="00:07:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:44.22" />
                    <SPLIT distance="150" swimtime="00:02:43.20" />
                    <SPLIT distance="200" swimtime="00:03:43.44" />
                    <SPLIT distance="250" swimtime="00:04:43.68" />
                    <SPLIT distance="300" swimtime="00:05:43.75" />
                    <SPLIT distance="350" swimtime="00:06:43.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-05-25" firstname="Włodzimierz" gender="M" lastname="Łatecki" nation="POL" license="503105700032" athleteid="3147">
              <RESULTS>
                <RESULT eventid="1108" points="43" swimtime="00:05:10.94" resultid="3148" heatid="7278" lane="8" entrytime="00:04:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:04:07.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="59" reactiontime="+99" swimtime="00:01:55.19" resultid="3149" heatid="7352" lane="9" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="32" reactiontime="+96" swimtime="00:05:39.37" resultid="3150" heatid="7394" lane="3" entrytime="00:05:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.36" />
                    <SPLIT distance="100" swimtime="00:02:35.16" />
                    <SPLIT distance="150" swimtime="00:04:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="62" reactiontime="+98" swimtime="00:04:10.00" resultid="3151" heatid="7476" lane="7" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.57" />
                    <SPLIT distance="100" swimtime="00:01:57.06" />
                    <SPLIT distance="150" swimtime="00:03:04.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="70" swimtime="00:08:33.08" resultid="3152" heatid="7583" lane="1" entrytime="00:07:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.49" />
                    <SPLIT distance="200" swimtime="00:04:10.68" />
                    <SPLIT distance="300" swimtime="00:06:23.30" />
                    <SPLIT distance="350" swimtime="00:07:28.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="3160">
              <RESULTS>
                <RESULT eventid="1092" points="439" reactiontime="+80" swimtime="00:02:40.25" resultid="3161" heatid="7274" lane="4" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:02:02.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="378" reactiontime="+82" swimtime="00:02:45.29" resultid="3162" heatid="7393" lane="6" entrytime="00:02:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="446" reactiontime="+75" swimtime="00:00:31.90" resultid="3163" heatid="7432" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1608" points="466" reactiontime="+81" swimtime="00:01:10.39" resultid="3164" heatid="7511" lane="9" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="415" reactiontime="+76" swimtime="00:00:38.28" resultid="3165" heatid="7543" lane="5" entrytime="00:00:39.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="130" reactiontime="+83" swimtime="00:02:58.10" resultid="3304" heatid="7403" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:38.28" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3207" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3095" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3124" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3135" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="132" swimtime="00:02:40.51" resultid="3305" heatid="7493" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                    <SPLIT distance="100" swimtime="00:01:28.62" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3207" number="1" />
                    <RELAYPOSITION athleteid="3095" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3124" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3135" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="222" reactiontime="+80" swimtime="00:02:29.14" resultid="3306" heatid="7404" lane="1" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:01:56.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3210" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3288" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3183" number="3" reactiontime="+11" />
                    <RELAYPOSITION athleteid="3257" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="264" reactiontime="+89" swimtime="00:02:07.45" resultid="3307" heatid="7494" lane="0" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="150" swimtime="00:01:36.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3117" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3257" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3183" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="3210" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="413" reactiontime="+64" swimtime="00:02:01.36" resultid="3308" heatid="7405" lane="6" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:33.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3192" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3219" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="3224" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3232" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1545" points="434" reactiontime="+75" swimtime="00:01:48.01" resultid="3309" heatid="7495" lane="2" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.82" />
                    <SPLIT distance="100" swimtime="00:00:54.99" />
                    <SPLIT distance="150" swimtime="00:01:22.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3224" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3219" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3232" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3198" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1545" points="221" reactiontime="+88" swimtime="00:02:15.18" resultid="3320" heatid="7494" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:48.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3130" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3288" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3238" number="3" reactiontime="+11" />
                    <RELAYPOSITION athleteid="3192" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1368" points="430" reactiontime="+76" swimtime="00:02:15.61" resultid="3316" heatid="7401" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:10.96" />
                    <SPLIT distance="150" swimtime="00:01:43.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3153" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3172" number="2" />
                    <RELAYPOSITION athleteid="3160" number="3" />
                    <RELAYPOSITION athleteid="3102" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1529" points="450" reactiontime="+81" swimtime="00:02:02.48" resultid="3317" heatid="7491" lane="2" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:33.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3160" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3110" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3172" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3153" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1529" status="DNS" swimtime="00:00:00.00" resultid="3318" heatid="7491" lane="0" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3274" number="1" />
                    <RELAYPOSITION athleteid="3292" number="2" />
                    <RELAYPOSITION athleteid="3300" number="3" />
                    <RELAYPOSITION athleteid="3166" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1368" points="189" reactiontime="+75" swimtime="00:02:58.11" resultid="3319" heatid="7400" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:46.50" />
                    <SPLIT distance="150" swimtime="00:02:22.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3274" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3300" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3166" number="3" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3292" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="281" reactiontime="+96" swimtime="00:02:14.10" resultid="3310" heatid="7288" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:32.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3124" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="3102" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="3135" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3153" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="288" reactiontime="+81" swimtime="00:02:25.95" resultid="3311" heatid="7564" lane="0" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3153" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3095" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3102" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3124" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="370" reactiontime="+76" swimtime="00:02:02.32" resultid="3312" heatid="7289" lane="1" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.72" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:35.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3198" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3274" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3160" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3224" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="492" reactiontime="+56" swimtime="00:02:02.11" resultid="3313" heatid="7565" lane="6" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:00:58.89" />
                    <SPLIT distance="150" swimtime="00:01:31.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3192" number="1" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3224" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="3160" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3172" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="333" reactiontime="+81" swimtime="00:02:06.80" resultid="3314" heatid="7288" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="150" swimtime="00:01:35.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3183" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3166" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3172" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3210" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="234" reactiontime="+85" swimtime="00:02:36.23" resultid="3315" heatid="7565" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:28.38" />
                    <SPLIT distance="150" swimtime="00:02:04.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3210" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3274" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3166" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3183" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="4550" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="marlena@masters.waw.pl" name="Dobrasiewicz" phone="516120337" street="Zólkiewskiego 40/11" zip="04-305" />
          <ATHLETES>
            <ATHLETE birthdate="1977-08-13" firstname="Dymitr" gender="M" lastname="Bielski" nation="POL" athleteid="4551">
              <RESULTS>
                <RESULT eventid="1256" points="295" reactiontime="+89" swimtime="00:03:00.45" resultid="4552" heatid="7337" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                    <SPLIT distance="150" swimtime="00:02:12.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="248" reactiontime="+88" swimtime="00:01:19.96" resultid="4553" heatid="7381" lane="2" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="295" reactiontime="+90" swimtime="00:01:23.51" resultid="4554" heatid="7422" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="245" reactiontime="+84" swimtime="00:02:38.77" resultid="4555" heatid="7480" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="205" reactiontime="+86" swimtime="00:01:21.51" resultid="4556" heatid="7516" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="4647">
              <RESULTS>
                <RESULT eventid="1076" points="128" reactiontime="+88" swimtime="00:00:40.16" resultid="4648" heatid="7250" lane="8" entrytime="00:00:39.90" />
                <RESULT eventid="1224" points="69" reactiontime="+81" swimtime="00:00:53.97" resultid="4649" heatid="7317" lane="5" entrytime="00:00:53.00" />
                <RESULT eventid="1288" points="114" reactiontime="+90" swimtime="00:01:32.63" resultid="4650" heatid="7352" lane="1" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-13" firstname="Justyna" gender="F" lastname="Dabrowska- Bien" nation="POL" athleteid="4592">
              <RESULTS>
                <RESULT eventid="1240" points="268" reactiontime="+82" swimtime="00:03:28.50" resultid="4593" heatid="7329" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.28" />
                    <SPLIT distance="100" swimtime="00:01:41.11" />
                    <SPLIT distance="150" swimtime="00:02:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="286" reactiontime="+90" swimtime="00:01:34.57" resultid="4594" heatid="7410" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="254" reactiontime="+79" swimtime="00:00:45.06" resultid="4595" heatid="7541" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-24" firstname="Marlena" gender="F" lastname="Dobrasiewicz" nation="POL" athleteid="4741">
              <RESULTS>
                <RESULT eventid="1240" points="482" reactiontime="+88" swimtime="00:02:51.54" resultid="4742" heatid="7331" lane="8" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="479" reactiontime="+90" swimtime="00:01:04.18" resultid="4743" heatid="7347" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="465" reactiontime="+84" swimtime="00:01:20.49" resultid="4744" heatid="7412" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="464" reactiontime="+88" swimtime="00:02:22.63" resultid="4745" heatid="7474" lane="8" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:46.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="4608">
              <RESULTS>
                <RESULT eventid="1240" points="305" reactiontime="+79" swimtime="00:03:19.78" resultid="4609" heatid="7330" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:36.16" />
                    <SPLIT distance="150" swimtime="00:02:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="332" reactiontime="+81" swimtime="00:01:21.54" resultid="4610" heatid="7374" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="323" reactiontime="+74" swimtime="00:00:35.51" resultid="4611" heatid="7432" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1561" points="291" reactiontime="+74" swimtime="00:06:30.58" resultid="4612" heatid="8151" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:30.56" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                    <SPLIT distance="200" swimtime="00:03:09.74" />
                    <SPLIT distance="250" swimtime="00:04:04.34" />
                    <SPLIT distance="300" swimtime="00:04:59.77" />
                    <SPLIT distance="350" swimtime="00:05:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="305" reactiontime="+78" swimtime="00:02:57.06" resultid="4613" heatid="7527" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                    <SPLIT distance="150" swimtime="00:02:11.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-26" firstname="Ewa" gender="F" lastname="Galica" nation="POL" athleteid="4659">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="4660" heatid="7242" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="4661" heatid="7344" lane="3" entrytime="00:01:15.50" />
                <RESULT eventid="1433" points="300" reactiontime="+83" swimtime="00:00:36.41" resultid="4662" heatid="7431" lane="9" entrytime="00:00:36.80" />
                <RESULT eventid="1497" points="345" reactiontime="+78" swimtime="00:02:37.36" resultid="4663" heatid="7472" lane="1" entrytime="00:02:41.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" status="DNS" swimtime="00:00:00.00" resultid="4664" heatid="7508" lane="1" entrytime="00:01:55.00" />
                <RESULT eventid="1721" points="379" reactiontime="+78" swimtime="00:05:23.18" resultid="4665" heatid="7567" lane="7" entrytime="00:05:34.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:57.13" />
                    <SPLIT distance="200" swimtime="00:02:39.09" />
                    <SPLIT distance="250" swimtime="00:03:21.13" />
                    <SPLIT distance="300" swimtime="00:04:02.76" />
                    <SPLIT distance="350" swimtime="00:04:44.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="4623">
              <RESULTS>
                <RESULT eventid="1156" points="394" reactiontime="+79" swimtime="00:10:04.72" resultid="4624" heatid="7294" lane="1" entrytime="00:10:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:44.48" />
                    <SPLIT distance="200" swimtime="00:02:21.91" />
                    <SPLIT distance="250" swimtime="00:02:59.93" />
                    <SPLIT distance="300" swimtime="00:03:38.29" />
                    <SPLIT distance="350" swimtime="00:04:16.61" />
                    <SPLIT distance="400" swimtime="00:04:54.89" />
                    <SPLIT distance="450" swimtime="00:05:33.50" />
                    <SPLIT distance="500" swimtime="00:06:13.03" />
                    <SPLIT distance="550" swimtime="00:06:52.10" />
                    <SPLIT distance="600" swimtime="00:07:32.03" />
                    <SPLIT distance="650" swimtime="00:08:11.76" />
                    <SPLIT distance="700" swimtime="00:08:50.20" />
                    <SPLIT distance="750" swimtime="00:09:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="430" reactiontime="+80" swimtime="00:00:59.53" resultid="4625" heatid="7361" lane="0" entrytime="00:01:02.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="368" reactiontime="+72" swimtime="00:00:30.34" resultid="4626" heatid="7442" lane="3" entrytime="00:00:32.30" />
                <RESULT eventid="1513" points="432" reactiontime="+72" swimtime="00:02:11.39" resultid="4627" heatid="7484" lane="8" entrytime="00:02:16.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="416" reactiontime="+68" swimtime="00:04:44.15" resultid="4628" heatid="7575" lane="1" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:06.34" />
                    <SPLIT distance="150" swimtime="00:01:42.52" />
                    <SPLIT distance="200" swimtime="00:02:18.48" />
                    <SPLIT distance="250" swimtime="00:02:54.52" />
                    <SPLIT distance="300" swimtime="00:03:31.44" />
                    <SPLIT distance="350" swimtime="00:04:08.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="4634">
              <RESULTS>
                <RESULT eventid="1256" points="90" swimtime="00:04:27.37" resultid="4635" heatid="7333" lane="6" entrytime="00:04:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.04" />
                    <SPLIT distance="100" swimtime="00:02:13.14" />
                    <SPLIT distance="150" swimtime="00:03:23.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="39" swimtime="00:05:18.75" resultid="4636" heatid="7394" lane="4" entrytime="00:04:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.65" />
                    <SPLIT distance="100" swimtime="00:02:40.83" />
                    <SPLIT distance="150" swimtime="00:04:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="90" swimtime="00:02:04.07" resultid="4637" heatid="7418" lane="9" entrytime="00:01:48.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="73" swimtime="00:00:51.89" resultid="4638" heatid="7437" lane="6" entrytime="00:00:46.55" />
                <RESULT eventid="1625" points="59" swimtime="00:02:03.09" resultid="4639" heatid="7514" lane="9" entrytime="00:01:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="145" swimtime="00:00:47.96" resultid="4640" heatid="7549" lane="4" entrytime="00:00:45.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-07-18" firstname="Damian" gender="M" lastname="Iwaniuk" nation="POL" athleteid="4746">
              <RESULTS>
                <RESULT eventid="1224" points="405" reactiontime="+85" swimtime="00:00:30.01" resultid="4747" heatid="7325" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1288" points="540" reactiontime="+82" swimtime="00:00:55.16" resultid="4748" heatid="7365" lane="3" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="488" reactiontime="+80" swimtime="00:00:27.61" resultid="4749" heatid="7448" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1513" points="486" reactiontime="+82" swimtime="00:02:06.33" resultid="4750" heatid="7487" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:01.97" />
                    <SPLIT distance="150" swimtime="00:01:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-13" firstname="Michal" gender="M" lastname="Jablonski" nation="POL" athleteid="4681">
              <RESULTS>
                <RESULT eventid="1288" points="315" reactiontime="+88" swimtime="00:01:05.99" resultid="4682" heatid="7358" lane="3" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="4683" heatid="7444" lane="6" entrytime="00:00:30.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="Jakalski" nation="POL" athleteid="4666">
              <RESULTS>
                <RESULT eventid="1224" points="400" reactiontime="+70" swimtime="00:00:30.15" resultid="4667" heatid="7324" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1288" points="412" reactiontime="+85" swimtime="00:01:00.37" resultid="4668" heatid="7363" lane="0" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="470" reactiontime="+84" swimtime="00:00:27.97" resultid="4669" heatid="7436" lane="1" />
                <RESULT eventid="1481" points="370" reactiontime="+70" swimtime="00:01:08.08" resultid="4670" heatid="7466" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="388" reactiontime="+83" swimtime="00:01:05.90" resultid="4671" heatid="7518" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="4672" heatid="7534" lane="3" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="4700">
              <RESULTS>
                <RESULT eventid="1059" points="364" reactiontime="+81" swimtime="00:00:32.09" resultid="4701" heatid="7239" lane="5" entrytime="00:00:34.90" />
                <RESULT eventid="1240" points="286" reactiontime="+84" swimtime="00:03:24.17" resultid="4702" heatid="7329" lane="5" entrytime="00:03:40.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:36.75" />
                    <SPLIT distance="150" swimtime="00:02:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="350" reactiontime="+75" swimtime="00:01:28.47" resultid="4703" heatid="7411" lane="9" entrytime="00:01:40.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="358" reactiontime="+77" swimtime="00:00:40.19" resultid="4704" heatid="7542" lane="8" entrytime="00:00:43.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-07" firstname="Daniel" gender="M" lastname="Julian Aguilar" nation="POL" athleteid="4586">
              <RESULTS>
                <RESULT eventid="1224" points="362" reactiontime="+63" swimtime="00:00:31.17" resultid="4587" heatid="7325" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1288" points="438" reactiontime="+71" swimtime="00:00:59.14" resultid="4588" heatid="7363" lane="8" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="4589" heatid="7387" lane="5" entrytime="00:01:07.50" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="4590" heatid="7466" lane="8" entrytime="00:01:07.50" />
                <RESULT eventid="1513" points="410" reactiontime="+70" swimtime="00:02:13.74" resultid="4591" heatid="7485" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:39.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-28" firstname="Konrad" gender="M" lastname="Karnaszewski" nation="POL" athleteid="4629">
              <RESULTS>
                <RESULT eventid="1076" points="635" reactiontime="+66" swimtime="00:00:23.57" resultid="4630" heatid="7270" lane="6" entrytime="00:00:23.30" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4631" heatid="7332" lane="1" />
                <RESULT eventid="1288" points="614" reactiontime="+63" swimtime="00:00:52.85" resultid="4632" heatid="7367" lane="1" entrytime="00:00:53.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="4633" heatid="7449" lane="8" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-05" firstname="Marta" gender="F" lastname="Kosla" nation="POL" athleteid="4684">
              <RESULTS>
                <RESULT eventid="1059" points="472" reactiontime="+83" swimtime="00:00:29.45" resultid="4685" heatid="7244" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1207" points="503" reactiontime="+79" swimtime="00:00:32.26" resultid="4686" heatid="7314" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1304" points="379" reactiontime="+83" swimtime="00:01:18.02" resultid="4687" heatid="7375" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="434" reactiontime="+78" swimtime="00:00:32.19" resultid="4688" heatid="7433" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1465" points="482" reactiontime="+72" swimtime="00:01:10.14" resultid="4689" heatid="7458" lane="4" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="410" reactiontime="+84" swimtime="00:02:40.49" resultid="4690" heatid="7528" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:01:59.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-27" firstname="Wojciech" gender="M" lastname="Kossowski" nation="POL" athleteid="4602">
              <RESULTS>
                <RESULT eventid="1108" points="156" reactiontime="+95" swimtime="00:03:23.60" resultid="4603" heatid="7279" lane="8" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                    <SPLIT distance="100" swimtime="00:01:43.28" />
                    <SPLIT distance="150" swimtime="00:02:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="4604" heatid="7335" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="1320" points="169" swimtime="00:01:30.82" resultid="4605" heatid="7380" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="217" swimtime="00:01:32.40" resultid="4606" heatid="7418" lane="5" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="226" swimtime="00:00:41.42" resultid="4607" heatid="7551" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="4614">
              <RESULTS>
                <RESULT eventid="1076" points="392" reactiontime="+86" swimtime="00:00:27.68" resultid="4615" heatid="7260" lane="7" entrytime="00:00:28.53" />
                <RESULT eventid="1108" points="353" reactiontime="+89" swimtime="00:02:35.02" resultid="4616" heatid="7282" lane="8" entrytime="00:02:38.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="409" reactiontime="+84" swimtime="00:01:00.50" resultid="4617" heatid="7360" lane="4" entrytime="00:01:02.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="360" reactiontime="+80" swimtime="00:01:10.64" resultid="4618" heatid="7387" lane="7" entrytime="00:01:09.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="4619" heatid="7421" lane="4" entrytime="00:01:20.24" />
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="4620" heatid="7483" lane="1" entrytime="00:02:19.87" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4621" heatid="7555" lane="8" entrytime="00:00:37.18" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="4622" heatid="7577" lane="5" entrytime="00:05:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="4641">
              <RESULTS>
                <RESULT eventid="1272" points="367" reactiontime="+77" swimtime="00:01:10.15" resultid="4642" heatid="7344" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="327" reactiontime="+79" swimtime="00:01:22.00" resultid="4643" heatid="7372" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="365" reactiontime="+78" swimtime="00:00:34.10" resultid="4644" heatid="7432" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1497" points="375" reactiontime="+77" swimtime="00:02:33.10" resultid="4645" heatid="7472" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:52.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="379" reactiontime="+78" swimtime="00:05:23.13" resultid="4646" heatid="7567" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                    <SPLIT distance="200" swimtime="00:02:37.96" />
                    <SPLIT distance="250" swimtime="00:03:20.24" />
                    <SPLIT distance="300" swimtime="00:04:02.24" />
                    <SPLIT distance="350" swimtime="00:04:43.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michal" gender="M" lastname="Nowak" nation="POL" athleteid="4723">
              <RESULTS>
                <RESULT eventid="1108" points="181" reactiontime="+96" swimtime="00:03:13.51" resultid="4724" heatid="7280" lane="7" entrytime="00:03:06.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:39.90" />
                    <SPLIT distance="150" swimtime="00:02:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="222" swimtime="00:03:18.35" resultid="4725" heatid="7336" lane="6" entrytime="00:03:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="100" swimtime="00:01:34.31" />
                    <SPLIT distance="150" swimtime="00:02:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="224" reactiontime="+88" swimtime="00:01:22.68" resultid="4726" heatid="7382" lane="5" entrytime="00:01:18.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="283" reactiontime="+90" swimtime="00:01:24.68" resultid="4727" heatid="7421" lane="0" entrytime="00:01:22.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="170" reactiontime="+88" swimtime="00:07:04.53" resultid="4728" heatid="8155" lane="5" entrytime="00:07:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:47.51" />
                    <SPLIT distance="200" swimtime="00:03:42.95" />
                    <SPLIT distance="250" swimtime="00:04:37.37" />
                    <SPLIT distance="300" swimtime="00:05:31.75" />
                    <SPLIT distance="350" swimtime="00:06:20.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="300" reactiontime="+81" swimtime="00:00:37.68" resultid="4729" heatid="7555" lane="0" entrytime="00:00:37.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="4712">
              <RESULTS>
                <RESULT eventid="1224" points="401" reactiontime="+74" swimtime="00:00:30.12" resultid="4713" heatid="7325" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1481" points="429" reactiontime="+71" swimtime="00:01:04.78" resultid="4714" heatid="7467" lane="0" entrytime="00:01:04.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="354" reactiontime="+67" swimtime="00:02:29.26" resultid="4715" heatid="7536" lane="1" entrytime="00:02:22.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:48.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-14" firstname="Bartosz" gender="M" lastname="Ostrowski" nation="POL" athleteid="4691">
              <RESULTS>
                <RESULT eventid="1076" points="438" reactiontime="+78" swimtime="00:00:26.66" resultid="4692" heatid="7260" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1156" points="345" reactiontime="+91" swimtime="00:10:32.14" resultid="4693" heatid="7297" lane="7" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                    <SPLIT distance="200" swimtime="00:02:30.96" />
                    <SPLIT distance="250" swimtime="00:03:11.00" />
                    <SPLIT distance="300" swimtime="00:03:51.51" />
                    <SPLIT distance="350" swimtime="00:04:32.16" />
                    <SPLIT distance="400" swimtime="00:05:12.56" />
                    <SPLIT distance="450" swimtime="00:05:53.14" />
                    <SPLIT distance="500" swimtime="00:06:33.51" />
                    <SPLIT distance="550" swimtime="00:07:14.25" />
                    <SPLIT distance="600" swimtime="00:07:54.56" />
                    <SPLIT distance="650" swimtime="00:08:34.69" />
                    <SPLIT distance="700" swimtime="00:09:14.67" />
                    <SPLIT distance="750" swimtime="00:09:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="252" reactiontime="+94" swimtime="00:00:35.16" resultid="4694" heatid="7321" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1288" points="447" reactiontime="+74" swimtime="00:00:58.77" resultid="4695" heatid="7359" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="481" reactiontime="+75" swimtime="00:01:10.97" resultid="4696" heatid="7423" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="372" reactiontime="+77" swimtime="00:00:30.24" resultid="4697" heatid="7441" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1625" points="316" reactiontime="+80" swimtime="00:01:10.55" resultid="4698" heatid="7516" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="494" reactiontime="+74" swimtime="00:00:31.93" resultid="4699" heatid="7558" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-02-17" firstname="Zbigniew" gender="M" lastname="Paluszak" nation="POL" athleteid="4570">
              <RESULTS>
                <RESULT eventid="1256" points="145" reactiontime="+80" swimtime="00:03:48.60" resultid="4571" heatid="7334" lane="8" entrytime="00:03:51.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.10" />
                    <SPLIT distance="100" swimtime="00:01:44.62" />
                    <SPLIT distance="150" swimtime="00:02:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="108" reactiontime="+76" swimtime="00:01:45.33" resultid="4572" heatid="7377" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="157" reactiontime="+84" swimtime="00:01:43.04" resultid="4573" heatid="7417" lane="2" entrytime="00:01:47.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="103" reactiontime="+84" swimtime="00:03:31.55" resultid="4574" heatid="7476" lane="3" entrytime="00:03:30.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                    <SPLIT distance="100" swimtime="00:01:41.09" />
                    <SPLIT distance="150" swimtime="00:02:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="160" reactiontime="+76" swimtime="00:00:46.48" resultid="4575" heatid="7549" lane="1" entrytime="00:00:47.36" />
                <RESULT eventid="1737" points="123" reactiontime="+71" swimtime="00:07:06.00" resultid="4576" heatid="7583" lane="7" entrytime="00:07:37.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="100" swimtime="00:01:38.46" />
                    <SPLIT distance="150" swimtime="00:02:33.29" />
                    <SPLIT distance="200" swimtime="00:03:27.20" />
                    <SPLIT distance="250" swimtime="00:04:21.33" />
                    <SPLIT distance="300" swimtime="00:05:15.45" />
                    <SPLIT distance="350" swimtime="00:06:11.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="4673">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4674" heatid="7266" lane="2" entrytime="00:00:26.45" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="4675" heatid="7325" lane="3" entrytime="00:00:30.45" />
                <RESULT eventid="1288" points="437" reactiontime="+76" swimtime="00:00:59.20" resultid="4676" heatid="7365" lane="8" entrytime="00:00:57.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="4677" heatid="7448" lane="2" entrytime="00:00:28.45" />
                <RESULT eventid="1513" points="440" reactiontime="+72" swimtime="00:02:10.57" resultid="4678" heatid="7486" lane="4" entrytime="00:02:06.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:02.46" />
                    <SPLIT distance="150" swimtime="00:01:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="390" reactiontime="+72" swimtime="00:00:34.55" resultid="4679" heatid="7553" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1737" points="429" reactiontime="+78" swimtime="00:04:41.23" resultid="4680" heatid="7573" lane="8" entrytime="00:04:39.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                    <SPLIT distance="150" swimtime="00:01:40.64" />
                    <SPLIT distance="200" swimtime="00:02:17.61" />
                    <SPLIT distance="250" swimtime="00:02:53.84" />
                    <SPLIT distance="300" swimtime="00:03:30.88" />
                    <SPLIT distance="350" swimtime="00:04:06.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-19" firstname="Emilia" gender="F" lastname="Saczynska" nation="POL" athleteid="4716">
              <RESULTS>
                <RESULT eventid="1092" points="351" swimtime="00:02:52.66" resultid="4717" heatid="7274" lane="0" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="150" swimtime="00:02:11.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="363" reactiontime="+94" swimtime="00:00:35.97" resultid="4718" heatid="7312" lane="5" entrytime="00:00:35.80" />
                <RESULT eventid="1304" points="340" reactiontime="+89" swimtime="00:01:20.92" resultid="4719" heatid="7373" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="296" reactiontime="+92" swimtime="00:00:36.56" resultid="4720" heatid="7431" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1465" points="357" reactiontime="+79" swimtime="00:01:17.55" resultid="4721" heatid="7456" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="375" reactiontime="+80" swimtime="00:02:45.22" resultid="4722" heatid="7527" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:02.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="4562">
              <RESULTS>
                <RESULT eventid="1076" points="21" swimtime="00:01:13.13" resultid="4563" heatid="7247" lane="6" entrytime="00:01:05.00" />
                <RESULT eventid="1224" points="16" reactiontime="+88" swimtime="00:01:27.98" resultid="4564" heatid="7316" lane="7" entrytime="00:01:20.00" />
                <RESULT eventid="1320" points="17" swimtime="00:03:12.18" resultid="4565" heatid="7377" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="21" swimtime="00:03:19.12" resultid="4566" heatid="7415" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="16" reactiontime="+90" swimtime="00:03:11.46" resultid="4567" heatid="7459" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="4568" heatid="7529" lane="2" entrytime="00:05:55.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="4569" heatid="7546" lane="3" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafal" gender="M" lastname="Skoskiewicz" nation="POL" athleteid="4577">
              <RESULTS>
                <RESULT eventid="1076" points="377" reactiontime="+89" swimtime="00:00:28.04" resultid="4578" heatid="7261" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1108" points="384" reactiontime="+89" swimtime="00:02:30.71" resultid="4579" heatid="7282" lane="1" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="315" reactiontime="+77" swimtime="00:00:32.64" resultid="4580" heatid="7324" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1320" points="403" reactiontime="+75" swimtime="00:01:08.00" resultid="4581" heatid="7386" lane="8" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="390" reactiontime="+76" swimtime="00:00:29.75" resultid="4582" heatid="7447" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1481" points="395" reactiontime="+71" swimtime="00:01:06.61" resultid="4583" heatid="7465" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="379" reactiontime="+79" swimtime="00:01:06.43" resultid="4584" heatid="7518" lane="0" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="348" reactiontime="+70" swimtime="00:02:30.11" resultid="4585" heatid="7534" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="4651">
              <RESULTS>
                <RESULT eventid="1076" points="134" reactiontime="+99" swimtime="00:00:39.52" resultid="4652" heatid="7250" lane="5" entrytime="00:00:38.57" />
                <RESULT eventid="1156" points="154" swimtime="00:13:46.59" resultid="4653" heatid="7298" lane="2" entrytime="00:13:10.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="150" swimtime="00:02:26.89" />
                    <SPLIT distance="200" swimtime="00:03:19.38" />
                    <SPLIT distance="250" swimtime="00:04:11.63" />
                    <SPLIT distance="300" swimtime="00:05:03.66" />
                    <SPLIT distance="450" swimtime="00:07:40.64" />
                    <SPLIT distance="500" swimtime="00:08:32.47" />
                    <SPLIT distance="550" swimtime="00:09:25.07" />
                    <SPLIT distance="600" swimtime="00:10:18.38" />
                    <SPLIT distance="650" swimtime="00:11:11.57" />
                    <SPLIT distance="700" swimtime="00:12:05.30" />
                    <SPLIT distance="750" swimtime="00:12:57.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="151" swimtime="00:01:24.34" resultid="4654" heatid="7352" lane="7" entrytime="00:01:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="92" reactiontime="+65" swimtime="00:01:51.20" resultid="4655" heatid="7377" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="100" swimtime="00:00:46.75" resultid="4656" heatid="7437" lane="7" entrytime="00:00:48.10" />
                <RESULT eventid="1513" points="158" swimtime="00:03:03.54" resultid="4657" heatid="7477" lane="5" entrytime="00:03:03.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="161" swimtime="00:06:29.88" resultid="4658" heatid="7581" lane="7" entrytime="00:06:27.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:32.90" />
                    <SPLIT distance="150" swimtime="00:02:23.10" />
                    <SPLIT distance="200" swimtime="00:03:14.36" />
                    <SPLIT distance="250" swimtime="00:04:04.52" />
                    <SPLIT distance="300" swimtime="00:04:54.57" />
                    <SPLIT distance="350" swimtime="00:05:43.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="4738">
              <RESULTS>
                <RESULT eventid="1140" points="96" swimtime="00:17:23.69" resultid="4739" heatid="7293" lane="4" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.69" />
                    <SPLIT distance="100" swimtime="00:02:04.77" />
                    <SPLIT distance="150" swimtime="00:03:11.09" />
                    <SPLIT distance="200" swimtime="00:04:17.47" />
                    <SPLIT distance="250" swimtime="00:05:23.55" />
                    <SPLIT distance="300" swimtime="00:06:29.23" />
                    <SPLIT distance="350" swimtime="00:07:34.20" />
                    <SPLIT distance="400" swimtime="00:08:39.55" />
                    <SPLIT distance="450" swimtime="00:09:45.20" />
                    <SPLIT distance="500" swimtime="00:10:50.52" />
                    <SPLIT distance="550" swimtime="00:11:55.72" />
                    <SPLIT distance="600" swimtime="00:13:00.44" />
                    <SPLIT distance="650" swimtime="00:14:06.29" />
                    <SPLIT distance="700" swimtime="00:15:12.21" />
                    <SPLIT distance="750" swimtime="00:16:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="84" reactiontime="+93" swimtime="00:08:53.52" resultid="4740" heatid="7571" lane="8" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="100" swimtime="00:02:07.76" />
                    <SPLIT distance="150" swimtime="00:03:15.87" />
                    <SPLIT distance="200" swimtime="00:04:23.77" />
                    <SPLIT distance="250" swimtime="00:05:30.66" />
                    <SPLIT distance="300" swimtime="00:06:38.27" />
                    <SPLIT distance="350" swimtime="00:07:49.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="4705">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4706" heatid="7262" lane="3" entrytime="00:00:27.80" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="4707" heatid="7322" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1288" points="418" reactiontime="+77" swimtime="00:01:00.10" resultid="4708" heatid="7361" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="365" reactiontime="+78" swimtime="00:00:30.42" resultid="4709" heatid="7443" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1513" points="398" reactiontime="+77" swimtime="00:02:15.07" resultid="4710" heatid="7484" lane="0" entrytime="00:02:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" status="WDR" swimtime="00:00:00.00" resultid="4711" heatid="7576" lane="2" entrytime="00:05:01.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-11" firstname="Bolek" gender="M" lastname="Szuter" nation="POL" athleteid="4557">
              <RESULTS>
                <RESULT eventid="1076" points="491" reactiontime="+74" swimtime="00:00:25.67" resultid="4558" heatid="7269" lane="7" entrytime="00:00:24.99" />
                <RESULT eventid="1288" points="547" reactiontime="+77" swimtime="00:00:54.95" resultid="4559" heatid="7367" lane="0" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters kategoria E" eventid="1513" points="549" reactiontime="+65" swimtime="00:02:01.34" resultid="4560" heatid="7488" lane="0" entrytime="00:02:02.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:00:59.89" />
                    <SPLIT distance="150" swimtime="00:01:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="497" reactiontime="+71" swimtime="00:04:27.91" resultid="4561" heatid="7574" lane="4" entrytime="00:04:40.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:39.19" />
                    <SPLIT distance="200" swimtime="00:02:14.04" />
                    <SPLIT distance="250" swimtime="00:02:48.67" />
                    <SPLIT distance="300" swimtime="00:03:23.47" />
                    <SPLIT distance="350" swimtime="00:03:56.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="4730">
              <RESULTS>
                <RESULT eventid="1076" points="531" reactiontime="+82" swimtime="00:00:25.01" resultid="4731" heatid="7269" lane="5" entrytime="00:00:24.60" />
                <RESULT eventid="1224" points="498" reactiontime="+66" swimtime="00:00:28.02" resultid="4732" heatid="7326" lane="6" entrytime="00:00:27.95" />
                <RESULT eventid="1320" points="525" reactiontime="+73" swimtime="00:01:02.30" resultid="4733" heatid="7390" lane="8" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="543" reactiontime="+73" swimtime="00:00:26.65" resultid="4734" heatid="7436" lane="8" />
                <RESULT eventid="1481" points="484" reactiontime="+70" swimtime="00:01:02.25" resultid="4735" heatid="7467" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="481" reactiontime="+75" swimtime="00:01:01.35" resultid="4736" heatid="7521" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="512" reactiontime="+69" swimtime="00:00:31.55" resultid="4737" heatid="7560" lane="0" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Miroslaw" gender="M" lastname="Warchol" nation="POL" athleteid="4596">
              <RESULTS>
                <RESULT eventid="1076" points="332" reactiontime="+94" swimtime="00:00:29.24" resultid="4597" heatid="7258" lane="5" entrytime="00:00:29.78" />
                <RESULT eventid="1108" points="278" reactiontime="+96" swimtime="00:02:47.83" resultid="4598" heatid="7281" lane="4" entrytime="00:02:44.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:02:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="329" reactiontime="+91" swimtime="00:01:05.09" resultid="4599" heatid="7356" lane="5" entrytime="00:01:09.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="282" reactiontime="+76" swimtime="00:01:14.52" resultid="4600" heatid="7464" lane="5" entrytime="00:01:15.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="280" reactiontime="+76" swimtime="00:02:41.43" resultid="4601" heatid="7534" lane="9" entrytime="00:02:42.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="zm męzczyzni I" number="6">
              <RESULTS>
                <RESULT eventid="1391" points="393" reactiontime="+76" swimtime="00:02:03.47" resultid="4756" heatid="7405" lane="5" entrytime="00:02:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:33.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4577" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4691" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4705" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4596" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="zm męzczyzni II" number="7">
              <RESULTS>
                <RESULT eventid="1391" points="519" reactiontime="+72" swimtime="00:01:52.50" resultid="4757" heatid="7406" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:00.55" />
                    <SPLIT distance="150" swimtime="00:01:27.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4730" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4712" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4629" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="4557" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="zm męzczyzni IV" number="8">
              <RESULTS>
                <RESULT eventid="1391" points="265" reactiontime="+69" swimtime="00:02:20.68" resultid="4758" heatid="7404" lane="2" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:01:49.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4666" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4634" number="2" />
                    <RELAYPOSITION athleteid="4681" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4551" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="dow męzczyzn I" number="9">
              <RESULTS>
                <RESULT eventid="1545" points="371" reactiontime="+78" swimtime="00:01:53.74" resultid="4759" heatid="7495" lane="8" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="100" swimtime="00:00:56.64" />
                    <SPLIT distance="150" swimtime="00:01:23.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4577" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4623" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="4705" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4596" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="dow męzczyzni II" number="10">
              <RESULTS>
                <RESULT eventid="1545" points="562" reactiontime="+71" swimtime="00:01:39.09" resultid="4760" heatid="7496" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.03" />
                    <SPLIT distance="100" swimtime="00:00:50.49" />
                    <SPLIT distance="150" swimtime="00:01:16.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4730" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4557" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="4673" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4629" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="zm męzczyzni III" number="12">
              <RESULTS>
                <RESULT eventid="1391" points="403" reactiontime="+62" swimtime="00:02:02.43" resultid="4762" heatid="7406" lane="9" entrytime="00:01:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:34.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4586" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4746" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4673" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4623" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="dow męzczyzni III" number="13">
              <RESULTS>
                <RESULT eventid="1545" points="478" reactiontime="+90" swimtime="00:01:44.56" resultid="4763" heatid="7496" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.40" />
                    <SPLIT distance="100" swimtime="00:00:51.56" />
                    <SPLIT distance="150" swimtime="00:01:18.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4746" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="4666" number="2" reactiontime="+9" />
                    <RELAYPOSITION athleteid="4586" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4712" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="dow kobiety" number="1">
              <RESULTS>
                <RESULT eventid="1529" points="451" reactiontime="+77" swimtime="00:02:02.38" resultid="4751" heatid="7491" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:01:01.08" />
                    <SPLIT distance="150" swimtime="00:01:33.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4684" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4641" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4659" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="4741" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="zm kobiety" number="11">
              <RESULTS>
                <RESULT eventid="1368" points="405" reactiontime="+71" swimtime="00:02:18.30" resultid="4761" heatid="7401" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:45.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4684" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4741" number="2" />
                    <RELAYPOSITION athleteid="4716" number="3" />
                    <RELAYPOSITION athleteid="4659" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="dow mix" number="2">
              <RESULTS>
                <RESULT eventid="1124" points="429" reactiontime="+74" swimtime="00:01:56.46" resultid="4752" heatid="7289" lane="3" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.58" />
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="150" swimtime="00:01:27.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4730" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4659" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4596" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="4684" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="zm mix I" number="3">
              <RESULTS>
                <RESULT eventid="1705" points="453" reactiontime="+70" swimtime="00:02:05.44" resultid="4753" heatid="7565" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="100" swimtime="00:01:01.68" />
                    <SPLIT distance="150" swimtime="00:01:32.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4730" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4712" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="4684" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4659" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="zm mix II" number="4">
              <RESULTS>
                <RESULT eventid="1705" points="389" reactiontime="+84" swimtime="00:02:12.05" resultid="4754" heatid="7564" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:01:46.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4716" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="4608" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4666" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="4673" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="zm mix III" number="5">
              <RESULTS>
                <RESULT eventid="1705" points="214" reactiontime="+73" swimtime="00:02:41.04" resultid="4755" heatid="7563" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:02:08.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4691" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4592" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4634" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4700" number="4" reactiontime="+81" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="2602" name="Warta Masters Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502 499 565" state="WIE" street="Osiedle Dębina 19 m 34" zip="661-450" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" license="500115600525" athleteid="5946">
              <RESULTS>
                <RESULT eventid="1059" points="75" swimtime="00:00:54.33" resultid="5947" heatid="7235" lane="2" entrytime="00:00:56.00" />
                <RESULT eventid="1240" points="107" swimtime="00:04:43.12" resultid="5948" heatid="7328" lane="0" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.63" />
                    <SPLIT distance="100" swimtime="00:02:14.21" />
                    <SPLIT distance="150" swimtime="00:03:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="109" swimtime="00:02:10.37" resultid="5949" heatid="7409" lane="9" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="116" reactiontime="+97" swimtime="00:00:58.41" resultid="5950" heatid="7539" lane="7" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="5989">
              <RESULTS>
                <RESULT eventid="1076" points="385" reactiontime="+75" swimtime="00:00:27.83" resultid="5990" heatid="7262" lane="7" entrytime="00:00:27.93" />
                <RESULT eventid="1156" points="348" reactiontime="+94" swimtime="00:10:30.29" resultid="5991" heatid="7294" lane="2" entrytime="00:09:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:48.02" />
                    <SPLIT distance="200" swimtime="00:02:26.10" />
                    <SPLIT distance="250" swimtime="00:03:04.51" />
                    <SPLIT distance="300" swimtime="00:03:43.07" />
                    <SPLIT distance="350" swimtime="00:04:22.74" />
                    <SPLIT distance="400" swimtime="00:05:02.74" />
                    <SPLIT distance="450" swimtime="00:05:42.95" />
                    <SPLIT distance="500" swimtime="00:06:23.35" />
                    <SPLIT distance="550" swimtime="00:07:03.79" />
                    <SPLIT distance="600" swimtime="00:07:44.96" />
                    <SPLIT distance="650" swimtime="00:08:26.38" />
                    <SPLIT distance="700" swimtime="00:09:08.11" />
                    <SPLIT distance="750" swimtime="00:09:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="341" reactiontime="+69" swimtime="00:00:31.79" resultid="5992" heatid="7324" lane="3" entrytime="00:00:31.71" />
                <RESULT eventid="1481" points="367" reactiontime="+67" swimtime="00:01:08.24" resultid="5993" heatid="7465" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="379" reactiontime="+81" swimtime="00:02:17.28" resultid="5994" heatid="7483" lane="2" entrytime="00:02:18.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="150" swimtime="00:01:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="335" reactiontime="+63" swimtime="00:02:32.01" resultid="5995" heatid="7534" lane="4" entrytime="00:02:34.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="364" reactiontime="+76" swimtime="00:04:57.02" resultid="5996" heatid="7575" lane="9" entrytime="00:04:54.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                    <SPLIT distance="200" swimtime="00:02:25.04" />
                    <SPLIT distance="250" swimtime="00:03:03.13" />
                    <SPLIT distance="300" swimtime="00:03:41.62" />
                    <SPLIT distance="350" swimtime="00:04:20.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="5951">
              <RESULTS>
                <RESULT eventid="1140" points="236" swimtime="00:12:55.20" resultid="5952" heatid="7292" lane="4" entrytime="00:13:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                    <SPLIT distance="150" swimtime="00:02:17.08" />
                    <SPLIT distance="200" swimtime="00:03:05.44" />
                    <SPLIT distance="250" swimtime="00:03:54.06" />
                    <SPLIT distance="300" swimtime="00:04:42.41" />
                    <SPLIT distance="350" swimtime="00:05:30.81" />
                    <SPLIT distance="400" swimtime="00:06:19.82" />
                    <SPLIT distance="450" swimtime="00:07:09.10" />
                    <SPLIT distance="500" swimtime="00:07:58.06" />
                    <SPLIT distance="550" swimtime="00:08:47.42" />
                    <SPLIT distance="600" swimtime="00:09:36.45" />
                    <SPLIT distance="650" swimtime="00:10:26.28" />
                    <SPLIT distance="700" swimtime="00:11:16.54" />
                    <SPLIT distance="750" swimtime="00:12:06.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" points="156" reactiontime="+91" swimtime="00:00:47.62" resultid="5953" heatid="7309" lane="1" entrytime="00:00:49.00" />
                <RESULT eventid="1272" points="192" swimtime="00:01:27.06" resultid="5954" heatid="7342" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="165" reactiontime="+76" swimtime="00:01:40.16" resultid="5955" heatid="7454" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="219" swimtime="00:03:02.94" resultid="5956" heatid="7470" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:28.99" />
                    <SPLIT distance="150" swimtime="00:02:16.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="188" reactiontime="+74" swimtime="00:03:27.79" resultid="5957" heatid="7525" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                    <SPLIT distance="100" swimtime="00:01:42.75" />
                    <SPLIT distance="150" swimtime="00:02:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="226" swimtime="00:06:23.67" resultid="5958" heatid="7569" lane="9" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                    <SPLIT distance="150" swimtime="00:02:15.98" />
                    <SPLIT distance="200" swimtime="00:03:05.58" />
                    <SPLIT distance="250" swimtime="00:03:55.77" />
                    <SPLIT distance="300" swimtime="00:04:45.77" />
                    <SPLIT distance="350" swimtime="00:05:35.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" license="500115600520" athleteid="5959">
              <RESULTS>
                <RESULT eventid="1059" points="134" swimtime="00:00:44.74" resultid="5960" heatid="7236" lane="6" entrytime="00:00:46.00" />
                <RESULT eventid="1240" points="167" swimtime="00:04:04.04" resultid="5961" heatid="7328" lane="3" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                    <SPLIT distance="100" swimtime="00:01:56.40" />
                    <SPLIT distance="150" swimtime="00:03:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="105" swimtime="00:01:46.34" resultid="5962" heatid="7341" lane="5" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="173" reactiontime="+98" swimtime="00:01:51.86" resultid="5963" heatid="7409" lane="5" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="104" swimtime="00:03:54.72" resultid="5964" heatid="7469" lane="9" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                    <SPLIT distance="100" swimtime="00:01:53.59" />
                    <SPLIT distance="150" swimtime="00:02:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="179" swimtime="00:00:50.67" resultid="5965" heatid="7539" lane="2" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-26" firstname="Oleksandr" gender="M" lastname="Kuchuk" nation="POL" athleteid="5997">
              <RESULTS>
                <RESULT eventid="1417" points="502" reactiontime="+78" swimtime="00:01:09.97" resultid="5998" heatid="7424" lane="5" entrytime="00:01:12.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="540" reactiontime="+73" swimtime="00:00:30.99" resultid="5999" heatid="7560" lane="2" entrytime="00:00:32.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-07-13" firstname="Paulina" gender="F" lastname="Mendowska" nation="POL" license="100115600340" athleteid="5966">
              <RESULTS>
                <RESULT eventid="1433" points="440" reactiontime="+73" swimtime="00:00:32.05" resultid="5967" heatid="7433" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1465" points="399" reactiontime="+76" swimtime="00:01:14.73" resultid="5968" heatid="7458" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="406" reactiontime="+73" swimtime="00:01:13.74" resultid="5969" heatid="7511" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="5970" heatid="7528" lane="2" entrytime="00:02:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" athleteid="6000">
              <RESULTS>
                <RESULT eventid="1288" points="388" reactiontime="+80" swimtime="00:01:01.57" resultid="6001" heatid="7360" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="362" reactiontime="+78" swimtime="00:02:19.32" resultid="6002" heatid="7483" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="330" reactiontime="+76" swimtime="00:05:06.94" resultid="6003" heatid="7576" lane="0" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:50.13" />
                    <SPLIT distance="200" swimtime="00:02:30.84" />
                    <SPLIT distance="250" swimtime="00:03:11.47" />
                    <SPLIT distance="300" swimtime="00:03:51.76" />
                    <SPLIT distance="350" swimtime="00:04:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-05" firstname="Filip" gender="M" lastname="Piotrowski" nation="POL" license="500115700522" athleteid="6004">
              <RESULTS>
                <RESULT eventid="1076" points="452" reactiontime="+82" swimtime="00:00:26.39" resultid="6005" heatid="7268" lane="9" entrytime="00:00:25.69" />
                <RESULT eventid="1156" points="370" reactiontime="+72" swimtime="00:10:17.54" resultid="6006" heatid="7294" lane="6" entrytime="00:09:54.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:46.80" />
                    <SPLIT distance="200" swimtime="00:02:24.53" />
                    <SPLIT distance="250" swimtime="00:03:03.01" />
                    <SPLIT distance="300" swimtime="00:03:42.03" />
                    <SPLIT distance="350" swimtime="00:04:21.00" />
                    <SPLIT distance="400" swimtime="00:04:59.60" />
                    <SPLIT distance="450" swimtime="00:05:38.71" />
                    <SPLIT distance="500" swimtime="00:06:18.26" />
                    <SPLIT distance="550" swimtime="00:06:58.18" />
                    <SPLIT distance="600" swimtime="00:07:38.02" />
                    <SPLIT distance="650" swimtime="00:08:18.54" />
                    <SPLIT distance="700" swimtime="00:08:59.72" />
                    <SPLIT distance="750" swimtime="00:09:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="458" reactiontime="+67" swimtime="00:00:58.26" resultid="6007" heatid="7365" lane="7" entrytime="00:00:57.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="377" reactiontime="+70" swimtime="00:02:29.79" resultid="6008" heatid="7398" lane="9" entrytime="00:02:30.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:52.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="6009" heatid="7448" lane="6" entrytime="00:00:28.30" />
                <RESULT eventid="1513" points="446" reactiontime="+70" swimtime="00:02:09.98" resultid="6010" heatid="7485" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="401" reactiontime="+65" swimtime="00:01:05.15" resultid="6011" heatid="7520" lane="4" entrytime="00:01:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="408" reactiontime="+69" swimtime="00:04:46.13" resultid="6012" heatid="7573" lane="1" entrytime="00:04:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="150" swimtime="00:01:46.23" />
                    <SPLIT distance="200" swimtime="00:02:23.45" />
                    <SPLIT distance="250" swimtime="00:02:59.63" />
                    <SPLIT distance="300" swimtime="00:03:36.15" />
                    <SPLIT distance="350" swimtime="00:04:12.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" license="500115600462" athleteid="5971">
              <RESULTS>
                <RESULT eventid="1092" points="129" reactiontime="+90" swimtime="00:04:00.80" resultid="5972" heatid="7271" lane="5" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                    <SPLIT distance="100" swimtime="00:01:56.69" />
                    <SPLIT distance="150" swimtime="00:03:00.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="128" reactiontime="+99" swimtime="00:30:24.89" resultid="5973" heatid="7301" lane="6" entrytime="00:31:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="100" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:42.09" />
                    <SPLIT distance="200" swimtime="00:03:41.43" />
                    <SPLIT distance="250" swimtime="00:04:40.80" />
                    <SPLIT distance="300" swimtime="00:05:41.51" />
                    <SPLIT distance="350" swimtime="00:06:43.37" />
                    <SPLIT distance="400" swimtime="00:07:44.27" />
                    <SPLIT distance="450" swimtime="00:08:45.19" />
                    <SPLIT distance="500" swimtime="00:09:46.93" />
                    <SPLIT distance="550" swimtime="00:10:47.50" />
                    <SPLIT distance="600" swimtime="00:11:49.58" />
                    <SPLIT distance="650" swimtime="00:12:50.60" />
                    <SPLIT distance="700" swimtime="00:13:52.51" />
                    <SPLIT distance="750" swimtime="00:14:54.04" />
                    <SPLIT distance="800" swimtime="00:15:56.49" />
                    <SPLIT distance="850" swimtime="00:16:58.35" />
                    <SPLIT distance="900" swimtime="00:18:00.89" />
                    <SPLIT distance="950" swimtime="00:19:03.71" />
                    <SPLIT distance="1000" swimtime="00:20:06.88" />
                    <SPLIT distance="1050" swimtime="00:21:08.77" />
                    <SPLIT distance="1100" swimtime="00:22:11.00" />
                    <SPLIT distance="1150" swimtime="00:23:14.23" />
                    <SPLIT distance="1200" swimtime="00:24:16.25" />
                    <SPLIT distance="1250" swimtime="00:25:17.78" />
                    <SPLIT distance="1300" swimtime="00:26:20.04" />
                    <SPLIT distance="1350" swimtime="00:27:22.40" />
                    <SPLIT distance="1400" swimtime="00:28:24.76" />
                    <SPLIT distance="1450" swimtime="00:29:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="177" reactiontime="+97" swimtime="00:03:59.62" resultid="5974" heatid="7328" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                    <SPLIT distance="100" swimtime="00:01:53.96" />
                    <SPLIT distance="150" swimtime="00:02:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="83" reactiontime="+90" swimtime="00:04:33.29" resultid="5975" heatid="7392" lane="9" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.64" />
                    <SPLIT distance="100" swimtime="00:02:06.68" />
                    <SPLIT distance="150" swimtime="00:03:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" status="DNS" swimtime="00:00:00.00" resultid="5976" heatid="7409" lane="3" entrytime="00:01:54.00" />
                <RESULT eventid="1561" points="140" reactiontime="+81" swimtime="00:08:18.09" resultid="5977" heatid="8149" lane="3" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:02:00.39" />
                    <SPLIT distance="150" swimtime="00:03:03.41" />
                    <SPLIT distance="200" swimtime="00:04:06.65" />
                    <SPLIT distance="250" swimtime="00:05:09.88" />
                    <SPLIT distance="300" swimtime="00:06:15.52" />
                    <SPLIT distance="350" swimtime="00:07:16.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="120" reactiontime="+92" swimtime="00:04:01.30" resultid="5978" heatid="7525" lane="7" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.21" />
                    <SPLIT distance="100" swimtime="00:01:56.91" />
                    <SPLIT distance="150" swimtime="00:03:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="201" reactiontime="+86" swimtime="00:00:48.73" resultid="5979" heatid="7540" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-12" firstname="Marcin" gender="M" lastname="Szymkowiak" nation="POL" license="500115700523" athleteid="6013">
              <RESULTS>
                <RESULT eventid="1076" points="518" reactiontime="+76" swimtime="00:00:25.22" resultid="6014" heatid="7268" lane="6" entrytime="00:00:25.36" />
                <RESULT eventid="1108" points="488" reactiontime="+73" swimtime="00:02:19.24" resultid="6015" heatid="7285" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="541" reactiontime="+73" swimtime="00:02:27.38" resultid="6016" heatid="7339" lane="6" entrytime="00:02:30.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="531" reactiontime="+68" swimtime="00:00:55.48" resultid="6017" heatid="7366" lane="2" entrytime="00:00:55.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="615" reactiontime="+73" swimtime="00:01:05.37" resultid="6018" heatid="7425" lane="7" entrytime="00:01:07.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="530" reactiontime="+71" swimtime="00:00:26.87" resultid="6019" heatid="7449" lane="9" entrytime="00:00:27.98" />
                <RESULT eventid="1689" points="647" reactiontime="+70" swimtime="00:00:29.19" resultid="6020" heatid="7561" lane="8" entrytime="00:00:29.90" />
                <RESULT eventid="1737" points="439" reactiontime="+75" swimtime="00:04:39.13" resultid="6021" heatid="7573" lane="7" entrytime="00:04:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:42.50" />
                    <SPLIT distance="200" swimtime="00:02:18.65" />
                    <SPLIT distance="250" swimtime="00:02:54.58" />
                    <SPLIT distance="300" swimtime="00:03:30.09" />
                    <SPLIT distance="350" swimtime="00:04:05.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700344" athleteid="6034">
              <RESULTS>
                <RESULT eventid="1156" points="184" swimtime="00:12:59.49" resultid="6035" heatid="7298" lane="8" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                    <SPLIT distance="150" swimtime="00:02:19.36" />
                    <SPLIT distance="200" swimtime="00:03:08.51" />
                    <SPLIT distance="250" swimtime="00:03:57.77" />
                    <SPLIT distance="300" swimtime="00:04:48.42" />
                    <SPLIT distance="350" swimtime="00:05:39.72" />
                    <SPLIT distance="450" swimtime="00:07:20.44" />
                    <SPLIT distance="500" swimtime="00:08:10.53" />
                    <SPLIT distance="550" swimtime="00:09:00.14" />
                    <SPLIT distance="600" swimtime="00:09:50.19" />
                    <SPLIT distance="650" swimtime="00:10:39.40" />
                    <SPLIT distance="700" swimtime="00:11:27.80" />
                    <SPLIT distance="750" swimtime="00:12:15.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="165" swimtime="00:03:16.99" resultid="6036" heatid="7396" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:37.63" />
                    <SPLIT distance="150" swimtime="00:02:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="171" swimtime="00:00:39.12" resultid="6037" heatid="7439" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1577" points="142" swimtime="00:07:30.91" resultid="6038" heatid="8155" lane="2" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                    <SPLIT distance="100" swimtime="00:01:43.89" />
                    <SPLIT distance="150" swimtime="00:02:47.61" />
                    <SPLIT distance="200" swimtime="00:03:48.16" />
                    <SPLIT distance="250" swimtime="00:04:50.79" />
                    <SPLIT distance="300" swimtime="00:05:54.60" />
                    <SPLIT distance="350" swimtime="00:06:44.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="147" swimtime="00:01:31.04" resultid="6039" heatid="7516" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="115" reactiontime="+88" swimtime="00:03:37.03" resultid="6040" heatid="7531" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:49.98" />
                    <SPLIT distance="150" swimtime="00:02:46.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-08" firstname="Błażej" gender="M" lastname="Wachowski" nation="POL" license="100115700545" athleteid="6022">
              <RESULTS>
                <RESULT eventid="1076" points="333" reactiontime="+94" swimtime="00:00:29.21" resultid="6023" heatid="7260" lane="4" entrytime="00:00:28.30" />
                <RESULT eventid="1156" points="340" swimtime="00:10:35.11" resultid="6024" heatid="7294" lane="8" entrytime="00:10:14.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:52.75" />
                    <SPLIT distance="200" swimtime="00:02:32.32" />
                    <SPLIT distance="250" swimtime="00:03:12.00" />
                    <SPLIT distance="300" swimtime="00:03:51.81" />
                    <SPLIT distance="350" swimtime="00:04:31.64" />
                    <SPLIT distance="400" swimtime="00:05:12.46" />
                    <SPLIT distance="450" swimtime="00:05:52.88" />
                    <SPLIT distance="500" swimtime="00:06:33.09" />
                    <SPLIT distance="550" swimtime="00:07:14.27" />
                    <SPLIT distance="600" swimtime="00:07:55.16" />
                    <SPLIT distance="650" swimtime="00:08:35.88" />
                    <SPLIT distance="700" swimtime="00:09:16.17" />
                    <SPLIT distance="750" swimtime="00:09:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="268" swimtime="00:02:47.80" resultid="6025" heatid="7397" lane="3" entrytime="00:02:44.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:02:00.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="345" reactiontime="+98" swimtime="00:02:21.61" resultid="6026" heatid="7483" lane="7" entrytime="00:02:18.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="277" reactiontime="+58" swimtime="00:01:13.71" resultid="6027" heatid="7517" lane="4" entrytime="00:01:11.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="332" reactiontime="+93" swimtime="00:05:06.26" resultid="6028" heatid="7576" lane="7" entrytime="00:05:04.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:52.86" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="250" swimtime="00:03:10.98" />
                    <SPLIT distance="300" swimtime="00:03:49.84" />
                    <SPLIT distance="350" swimtime="00:04:28.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="6029">
              <RESULTS>
                <RESULT eventid="1108" points="217" swimtime="00:03:02.41" resultid="6030" heatid="7281" lane="0" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                    <SPLIT distance="150" swimtime="00:02:17.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="259" reactiontime="+91" swimtime="00:03:08.35" resultid="6031" heatid="7336" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:27.78" />
                    <SPLIT distance="150" swimtime="00:02:17.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="289" reactiontime="+88" swimtime="00:01:24.03" resultid="6032" heatid="7420" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="291" reactiontime="+89" swimtime="00:00:38.06" resultid="6033" heatid="7552" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-12" firstname="Włodzimierz" gender="M" lastname="Wiatr " nation="POL" athleteid="2601">
              <RESULTS>
                <RESULT eventid="1108" points="118" swimtime="00:03:43.35" resultid="2603" heatid="7279" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                    <SPLIT distance="100" swimtime="00:01:50.95" />
                    <SPLIT distance="150" swimtime="00:02:53.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="145" swimtime="00:14:03.98" resultid="2604" heatid="7299" lane="5" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:35.74" />
                    <SPLIT distance="150" swimtime="00:02:28.07" />
                    <SPLIT distance="200" swimtime="00:03:22.91" />
                    <SPLIT distance="250" swimtime="00:04:16.57" />
                    <SPLIT distance="300" swimtime="00:05:11.27" />
                    <SPLIT distance="350" swimtime="00:06:06.14" />
                    <SPLIT distance="400" swimtime="00:07:00.47" />
                    <SPLIT distance="450" swimtime="00:07:54.21" />
                    <SPLIT distance="500" swimtime="00:08:47.99" />
                    <SPLIT distance="550" swimtime="00:09:40.94" />
                    <SPLIT distance="600" swimtime="00:10:34.05" />
                    <SPLIT distance="650" swimtime="00:11:27.49" />
                    <SPLIT distance="700" swimtime="00:12:21.12" />
                    <SPLIT distance="750" swimtime="00:13:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="113" swimtime="00:01:43.80" resultid="2605" heatid="7378" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="118" swimtime="00:08:00.04" resultid="2606" heatid="8153" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                    <SPLIT distance="100" swimtime="00:02:00.72" />
                    <SPLIT distance="150" swimtime="00:03:04.04" />
                    <SPLIT distance="200" swimtime="00:04:08.45" />
                    <SPLIT distance="250" swimtime="00:05:12.92" />
                    <SPLIT distance="300" swimtime="00:06:16.29" />
                    <SPLIT distance="350" swimtime="00:07:08.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Szymon" gender="M" lastname="Wieja" nation="POL" license="500115700467" athleteid="6041">
              <RESULTS>
                <RESULT eventid="1076" points="492" reactiontime="+67" swimtime="00:00:25.65" resultid="6042" heatid="7268" lane="2" entrytime="00:00:25.49" />
                <RESULT eventid="1108" points="481" reactiontime="+68" swimtime="00:02:19.83" resultid="6043" heatid="7285" lane="5" entrytime="00:02:16.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="416" reactiontime="+56" swimtime="00:00:29.75" resultid="6044" heatid="7326" lane="8" entrytime="00:00:29.60" />
                <RESULT eventid="1288" points="508" reactiontime="+66" swimtime="00:00:56.32" resultid="6045" heatid="7366" lane="6" entrytime="00:00:55.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="439" reactiontime="+66" swimtime="00:00:28.61" resultid="6046" heatid="7448" lane="7" entrytime="00:00:28.49" />
                <RESULT eventid="1481" points="423" reactiontime="+61" swimtime="00:01:05.08" resultid="6047" heatid="7466" lane="2" entrytime="00:01:06.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="389" reactiontime="+66" swimtime="00:02:24.60" resultid="6048" heatid="7536" lane="0" entrytime="00:02:24.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="424" reactiontime="+65" swimtime="00:00:33.59" resultid="6049" heatid="7559" lane="0" entrytime="00:00:33.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-11" firstname="Piotr" gender="M" lastname="Witt" nation="POL" license="500115700548" athleteid="6050">
              <RESULTS>
                <RESULT eventid="1076" points="538" swimtime="00:00:24.91" resultid="6051" heatid="7270" lane="0" entrytime="00:00:24.41" />
                <RESULT eventid="1224" points="413" reactiontime="+67" swimtime="00:00:29.83" resultid="6052" heatid="7326" lane="0" entrytime="00:00:29.78" />
                <RESULT eventid="1288" points="585" reactiontime="+68" swimtime="00:00:53.71" resultid="6053" heatid="7367" lane="8" entrytime="00:00:54.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="473" reactiontime="+73" swimtime="00:00:27.91" resultid="6054" heatid="7449" lane="2" entrytime="00:00:27.49" />
                <RESULT eventid="1513" points="497" reactiontime="+70" swimtime="00:02:05.41" resultid="6055" heatid="7486" lane="2" entrytime="00:02:08.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="100" swimtime="00:00:58.92" />
                    <SPLIT distance="150" swimtime="00:01:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="428" reactiontime="+74" swimtime="00:01:03.75" resultid="6056" heatid="7519" lane="7" entrytime="00:01:06.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="428" reactiontime="+76" swimtime="00:04:41.62" resultid="6057" heatid="7575" lane="8" entrytime="00:04:52.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:05.64" />
                    <SPLIT distance="150" swimtime="00:01:41.59" />
                    <SPLIT distance="200" swimtime="00:02:17.56" />
                    <SPLIT distance="250" swimtime="00:02:54.07" />
                    <SPLIT distance="300" swimtime="00:03:30.59" />
                    <SPLIT distance="350" swimtime="00:04:07.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-01" firstname="Natalia" gender="F" lastname="Wiśniewska" nation="POL" license="500115600544" athleteid="5980">
              <RESULTS>
                <RESULT eventid="1092" points="526" reactiontime="+76" swimtime="00:02:30.88" resultid="5981" heatid="7275" lane="5" entrytime="00:02:29.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="475" reactiontime="+80" swimtime="00:10:13.96" resultid="5982" heatid="7290" lane="5" entrytime="00:09:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:47.54" />
                    <SPLIT distance="200" swimtime="00:02:25.73" />
                    <SPLIT distance="250" swimtime="00:03:04.06" />
                    <SPLIT distance="300" swimtime="00:03:42.16" />
                    <SPLIT distance="350" swimtime="00:04:20.77" />
                    <SPLIT distance="400" swimtime="00:04:59.60" />
                    <SPLIT distance="450" swimtime="00:05:38.57" />
                    <SPLIT distance="500" swimtime="00:06:18.10" />
                    <SPLIT distance="550" swimtime="00:06:57.87" />
                    <SPLIT distance="600" swimtime="00:07:37.23" />
                    <SPLIT distance="650" swimtime="00:08:16.59" />
                    <SPLIT distance="700" swimtime="00:08:55.89" />
                    <SPLIT distance="750" swimtime="00:09:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="577" reactiontime="+72" swimtime="00:02:41.59" resultid="5983" heatid="7331" lane="4" entrytime="00:02:41.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:01:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="535" reactiontime="+74" swimtime="00:01:09.58" resultid="5984" heatid="7376" lane="7" entrytime="00:01:09.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="585" reactiontime="+72" swimtime="00:01:14.56" resultid="5985" heatid="7413" lane="4" entrytime="00:01:14.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1561" points="528" reactiontime="+72" swimtime="00:05:20.27" resultid="5986" heatid="8151" lane="5" entrytime="00:05:23.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:02:34.67" />
                    <SPLIT distance="250" swimtime="00:03:18.19" />
                    <SPLIT distance="300" swimtime="00:04:02.40" />
                    <SPLIT distance="350" swimtime="00:04:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="601" reactiontime="+72" swimtime="00:00:33.83" resultid="5987" heatid="7545" lane="4" entrytime="00:00:33.69" />
                <RESULT eventid="1721" points="488" reactiontime="+70" swimtime="00:04:56.94" resultid="5988" heatid="7566" lane="6" entrytime="00:04:54.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:47.01" />
                    <SPLIT distance="200" swimtime="00:02:25.76" />
                    <SPLIT distance="250" swimtime="00:03:04.15" />
                    <SPLIT distance="300" swimtime="00:03:42.38" />
                    <SPLIT distance="350" swimtime="00:04:19.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 1" number="1">
              <RESULTS>
                <RESULT eventid="1391" points="484" reactiontime="+65" swimtime="00:01:55.14" resultid="6058" heatid="7406" lane="7" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:00:58.85" />
                    <SPLIT distance="150" swimtime="00:01:27.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6041" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="6013" number="2" reactiontime="+2" />
                    <RELAYPOSITION athleteid="6004" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="5989" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 7" number="2">
              <RESULTS>
                <RESULT eventid="1545" points="499" reactiontime="+68" swimtime="00:01:43.13" resultid="6059" heatid="7496" lane="1" entrytime="00:01:43.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                    <SPLIT distance="100" swimtime="00:00:52.93" />
                    <SPLIT distance="150" swimtime="00:01:19.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6041" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="5989" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="6004" number="3" reactiontime="+20" />
                    <RELAYPOSITION athleteid="6013" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WARTA 5" number="5">
              <RESULTS>
                <RESULT eventid="1545" points="435" reactiontime="+70" swimtime="00:01:47.95" resultid="6062" heatid="7495" lane="3" entrytime="00:01:48.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.68" />
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="150" swimtime="00:01:20.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6050" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5997" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="6022" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="6000" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WARTA 6" number="6">
              <RESULTS>
                <RESULT eventid="1391" points="383" reactiontime="+95" swimtime="00:02:04.53" resultid="6063" heatid="7405" lane="3" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:32.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6000" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="5997" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="6050" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="6029" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="WARTA 4" number="4">
              <RESULTS>
                <RESULT eventid="1368" points="129" swimtime="00:03:22.50" resultid="6061" heatid="7400" lane="8" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:45.76" />
                    <SPLIT distance="150" swimtime="00:02:07.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5951" number="1" />
                    <RELAYPOSITION athleteid="5946" number="2" />
                    <RELAYPOSITION athleteid="5971" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5959" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="WARTA 7" number="7">
              <RESULTS>
                <RESULT eventid="1529" points="128" swimtime="00:03:06.23" resultid="6064" heatid="7490" lane="8" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:19.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5951" number="1" />
                    <RELAYPOSITION athleteid="5971" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="5946" number="3" />
                    <RELAYPOSITION athleteid="5959" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="WARTA 3" number="3">
              <RESULTS>
                <RESULT eventid="1705" points="225" reactiontime="+93" swimtime="00:02:38.41" resultid="6060" heatid="7563" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5951" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="5997" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="5971" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="6029" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="WARTA 8" number="8">
              <RESULTS>
                <RESULT eventid="1124" points="237" reactiontime="+71" swimtime="00:02:21.89" resultid="6065" heatid="7287" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:48.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6050" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5959" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="5971" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="6029" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02611" nation="POL" region="11" clubid="3762" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="102611600021" athleteid="3763">
              <RESULTS>
                <RESULT eventid="1076" points="260" reactiontime="+81" swimtime="00:00:31.74" resultid="3764" heatid="7256" lane="9" entrytime="00:00:31.80" />
                <RESULT eventid="1224" points="170" reactiontime="+74" swimtime="00:00:40.11" resultid="3765" heatid="7320" lane="8" entrytime="00:00:40.24" />
                <RESULT eventid="1288" points="247" reactiontime="+96" swimtime="00:01:11.56" resultid="3766" heatid="7356" lane="0" entrytime="00:01:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="213" reactiontime="+85" swimtime="00:00:36.37" resultid="3767" heatid="7440" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1481" points="173" reactiontime="+83" swimtime="00:01:27.66" resultid="3768" heatid="7463" lane="7" entrytime="00:01:24.85" />
                <RESULT eventid="1657" points="160" reactiontime="+75" swimtime="00:03:14.33" resultid="3769" heatid="7532" lane="8" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="102611600023" athleteid="3776">
              <RESULTS>
                <RESULT eventid="1059" points="201" swimtime="00:00:39.11" resultid="3777" heatid="7238" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1207" points="143" reactiontime="+72" swimtime="00:00:49.05" resultid="3778" heatid="7309" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="1465" points="130" reactiontime="+68" swimtime="00:01:48.51" resultid="3780" heatid="7453" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="125" reactiontime="+85" swimtime="00:00:57.01" resultid="3781" heatid="7538" lane="8" entrytime="00:01:05.00" />
                <RESULT eventid="1304" points="147" reactiontime="+92" swimtime="00:01:47.04" resultid="5192" heatid="7369" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="102611600014" athleteid="3813">
              <RESULTS>
                <RESULT eventid="1076" points="96" reactiontime="+95" swimtime="00:00:44.16" resultid="3814" heatid="7249" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="3815" heatid="7437" lane="3" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="3770">
              <RESULTS>
                <RESULT eventid="1059" points="70" swimtime="00:00:55.62" resultid="3771" heatid="7235" lane="8" entrytime="00:01:05.00" />
                <RESULT eventid="1207" points="70" reactiontime="+78" swimtime="00:01:02.02" resultid="3772" heatid="7307" lane="6" entrytime="00:01:08.00" />
                <RESULT eventid="1240" points="81" reactiontime="+99" swimtime="00:05:10.24" resultid="3773" heatid="7328" lane="1" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.21" />
                    <SPLIT distance="100" swimtime="00:02:29.42" />
                    <SPLIT distance="150" swimtime="00:03:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="76" swimtime="00:02:26.60" resultid="3774" heatid="7408" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="110" swimtime="00:00:59.44" resultid="3775" heatid="7538" lane="0" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-02-18" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" license="502611100006" athleteid="3786">
              <RESULTS>
                <RESULT eventid="1059" points="197" swimtime="00:00:39.36" resultid="3787" heatid="7237" lane="3" entrytime="00:00:40.80" />
                <RESULT eventid="1207" points="221" reactiontime="+73" swimtime="00:00:42.45" resultid="3788" heatid="7310" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1304" points="181" reactiontime="+86" swimtime="00:01:39.80" resultid="3789" heatid="7371" lane="8" entrytime="00:01:35.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="162" reactiontime="+85" swimtime="00:00:44.72" resultid="3790" heatid="7428" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1465" points="197" reactiontime="+78" swimtime="00:01:34.46" resultid="3791" heatid="7455" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="204" reactiontime="+76" swimtime="00:03:22.49" resultid="3792" heatid="7526" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:38.38" />
                    <SPLIT distance="150" swimtime="00:02:30.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="102611600015" athleteid="3793">
              <RESULTS>
                <RESULT eventid="1076" points="224" swimtime="00:00:33.35" resultid="3794" heatid="7255" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1288" points="183" reactiontime="+94" swimtime="00:01:19.05" resultid="3795" heatid="7353" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="140" reactiontime="+97" swimtime="00:01:36.63" resultid="3796" heatid="7380" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="191" reactiontime="+93" swimtime="00:00:37.75" resultid="3797" heatid="7440" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1689" points="166" reactiontime="+90" swimtime="00:00:45.93" resultid="3798" heatid="7549" lane="5" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-04-14" firstname="Gabriela" gender="F" lastname="Molenda" nation="POL" athleteid="3806">
              <RESULTS>
                <RESULT eventid="1059" points="163" swimtime="00:00:41.90" resultid="3807" heatid="7237" lane="7" entrytime="00:00:42.60" />
                <RESULT eventid="1207" points="111" reactiontime="+93" swimtime="00:00:53.37" resultid="3808" heatid="7308" lane="3" entrytime="00:00:54.29" />
                <RESULT eventid="1272" points="152" reactiontime="+96" swimtime="00:01:34.15" resultid="3809" heatid="7342" lane="1" entrytime="00:01:33.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1465" points="118" reactiontime="+79" swimtime="00:01:52.11" resultid="3810" heatid="7453" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="141" reactiontime="+99" swimtime="00:03:32.14" resultid="3811" heatid="7469" lane="6" entrytime="00:03:29.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                    <SPLIT distance="100" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="126" reactiontime="+89" swimtime="00:03:57.68" resultid="3812" heatid="7525" lane="2" entrytime="00:03:56.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.25" />
                    <SPLIT distance="100" swimtime="00:01:56.10" />
                    <SPLIT distance="150" swimtime="00:02:57.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611100004" athleteid="3782">
              <RESULTS>
                <RESULT eventid="1224" points="132" reactiontime="+73" swimtime="00:00:43.54" resultid="3783" heatid="7319" lane="0" entrytime="00:00:43.89" />
                <RESULT eventid="1481" points="120" reactiontime="+71" swimtime="00:01:39.09" resultid="3784" heatid="7462" lane="1" entrytime="00:01:39.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="107" reactiontime="+74" swimtime="00:03:41.81" resultid="3785" heatid="7531" lane="0" entrytime="00:03:48.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                    <SPLIT distance="100" swimtime="00:01:44.87" />
                    <SPLIT distance="150" swimtime="00:02:43.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="102611600016" athleteid="3799">
              <RESULTS>
                <RESULT eventid="1140" points="441" reactiontime="+74" swimtime="00:10:29.42" resultid="3800" heatid="7290" lane="3" entrytime="00:10:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                    <SPLIT distance="200" swimtime="00:02:32.92" />
                    <SPLIT distance="250" swimtime="00:03:12.63" />
                    <SPLIT distance="300" swimtime="00:03:52.44" />
                    <SPLIT distance="350" swimtime="00:04:32.62" />
                    <SPLIT distance="400" swimtime="00:05:12.49" />
                    <SPLIT distance="450" swimtime="00:05:52.50" />
                    <SPLIT distance="500" swimtime="00:06:32.31" />
                    <SPLIT distance="550" swimtime="00:07:11.85" />
                    <SPLIT distance="600" swimtime="00:07:51.45" />
                    <SPLIT distance="650" swimtime="00:08:31.07" />
                    <SPLIT distance="700" swimtime="00:09:11.07" />
                    <SPLIT distance="750" swimtime="00:09:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="390" reactiontime="+73" swimtime="00:03:04.08" resultid="3801" heatid="7331" lane="3" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="404" reactiontime="+86" swimtime="00:01:24.35" resultid="3802" heatid="7413" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="432" reactiontime="+86" swimtime="00:02:25.98" resultid="3803" heatid="7473" lane="4" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="394" reactiontime="+82" swimtime="00:00:38.93" resultid="3804" heatid="7543" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1721" points="444" reactiontime="+94" swimtime="00:05:06.46" resultid="3805" heatid="7566" lane="1" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:14.11" />
                    <SPLIT distance="150" swimtime="00:01:52.77" />
                    <SPLIT distance="200" swimtime="00:02:31.84" />
                    <SPLIT distance="250" swimtime="00:03:10.85" />
                    <SPLIT distance="300" swimtime="00:03:49.94" />
                    <SPLIT distance="350" swimtime="00:04:28.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utraciły kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 13:30)" eventid="1368" reactiontime="+89" status="DSQ" swimtime="00:02:56.33" resultid="3816" heatid="7400" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3786" number="1" reactiontime="+89" status="DSQ" />
                    <RELAYPOSITION athleteid="3799" number="2" reactiontime="-81" status="DSQ" />
                    <RELAYPOSITION athleteid="3776" number="3" reactiontime="+57" status="DSQ" />
                    <RELAYPOSITION athleteid="3806" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1529" points="221" reactiontime="+87" swimtime="00:02:35.28" resultid="3818" heatid="7490" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3776" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3806" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3786" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3799" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1705" points="177" reactiontime="+71" swimtime="00:02:51.52" resultid="3817" heatid="7563" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:34.43" />
                    <SPLIT distance="150" swimtime="00:02:12.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3782" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3786" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3793" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3776" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1124" points="160" swimtime="00:02:41.77" resultid="3819" heatid="7287" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                    <SPLIT distance="150" swimtime="00:02:06.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3813" number="1" />
                    <RELAYPOSITION athleteid="3776" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3786" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3793" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00601" nation="POL" region="01" clubid="4920" name="WKS Śląsk Wrocław" shortname="Śląsk Wrocław">
          <CONTACT email="marrot68@wp.pl" name="Rother Marek" phone="785209045" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="4921">
              <RESULTS>
                <RESULT eventid="1224" points="397" reactiontime="+64" swimtime="00:00:30.21" resultid="4922" heatid="7324" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1320" points="390" reactiontime="+75" swimtime="00:01:08.76" resultid="4923" heatid="7387" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="410" reactiontime="+67" swimtime="00:01:05.75" resultid="4924" heatid="7465" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="397" reactiontime="+72" swimtime="00:02:23.68" resultid="4925" heatid="7535" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:47.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKIY" nation="UKR" clubid="2844" name="Wolfpack SC Kyiv">
          <ATHLETES>
            <ATHLETE birthdate="1983-11-15" firstname="Nadia" gender="F" lastname="Fedorovska" nation="UKR" athleteid="2861">
              <RESULTS>
                <RESULT eventid="1092" reactiontime="+74" status="DNF" swimtime="00:00:00.00" resultid="2862" heatid="7272" lane="6" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="300" reactiontime="+82" swimtime="00:01:14.99" resultid="2863" heatid="7343" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="256" reactiontime="+81" swimtime="00:01:28.93" resultid="2864" heatid="7372" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="256" reactiontime="+87" swimtime="00:00:38.38" resultid="2865" heatid="7429" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1497" points="271" reactiontime="+82" swimtime="00:02:50.59" resultid="2866" heatid="7471" lane="0" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                    <SPLIT distance="150" swimtime="00:02:08.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1608" points="209" reactiontime="+88" swimtime="00:01:31.99" resultid="2867" heatid="7509" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-06-01" firstname="Oleksandr" gender="M" lastname="Linyvyi" nation="UKR" athleteid="2843">
              <RESULTS>
                <RESULT eventid="1076" points="260" reactiontime="+79" swimtime="00:00:31.72" resultid="2845" heatid="7254" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1288" points="224" reactiontime="+81" swimtime="00:01:13.99" resultid="2846" heatid="7353" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="185" reactiontime="+87" swimtime="00:01:28.08" resultid="2847" heatid="7380" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="194" reactiontime="+78" swimtime="00:00:37.53" resultid="2848" heatid="7440" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="1513" points="168" reactiontime="+94" swimtime="00:02:59.95" resultid="2849" heatid="7478" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="154" reactiontime="+77" swimtime="00:01:29.54" resultid="2850" heatid="7515" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="144" reactiontime="+95" swimtime="00:06:44.21" resultid="2851" heatid="7582" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:34.97" />
                    <SPLIT distance="150" swimtime="00:02:27.54" />
                    <SPLIT distance="200" swimtime="00:03:20.62" />
                    <SPLIT distance="250" swimtime="00:04:12.14" />
                    <SPLIT distance="300" swimtime="00:05:04.03" />
                    <SPLIT distance="350" swimtime="00:05:55.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-17" firstname="Yevhen " gender="M" lastname="Samoilenko" nation="UKR" athleteid="2852">
              <RESULTS>
                <RESULT eventid="1076" points="568" reactiontime="+81" swimtime="00:00:24.45" resultid="2853" heatid="7270" lane="9" entrytime="00:00:24.50" />
                <RESULT eventid="1108" points="474" reactiontime="+87" swimtime="00:02:20.58" resultid="2854" heatid="7283" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="580" reactiontime="+72" swimtime="00:00:53.87" resultid="2855" heatid="7366" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="546" reactiontime="+68" swimtime="00:01:01.49" resultid="2856" heatid="7388" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="594" reactiontime="+72" swimtime="00:00:25.87" resultid="2857" heatid="7451" lane="9" entrytime="00:00:26.00" />
                <RESULT eventid="1513" points="498" reactiontime="+68" swimtime="00:02:05.33" resultid="2858" heatid="7486" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1625" points="497" reactiontime="+75" swimtime="00:01:00.68" resultid="2859" heatid="7520" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1737" points="441" reactiontime="+76" swimtime="00:04:38.67" resultid="2860" heatid="7574" lane="8" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                    <SPLIT distance="150" swimtime="00:01:43.12" />
                    <SPLIT distance="200" swimtime="00:02:19.76" />
                    <SPLIT distance="250" swimtime="00:02:56.56" />
                    <SPLIT distance="300" swimtime="00:03:32.17" />
                    <SPLIT distance="350" swimtime="00:04:05.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00000" nation="POL" clubid="2016" name="Zawodnik Niezrzeszomy">
          <CONTACT city="ŚWIECIE" name="KLONOWSKI" phone="6061229393" street="RZEPAKOWA 3" zip="86-100" />
          <ATHLETES>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="3395">
              <RESULTS>
                <RESULT eventid="1076" points="373" reactiontime="+92" swimtime="00:00:28.13" resultid="3396" heatid="7262" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1188" points="339" reactiontime="+98" swimtime="00:20:15.44" resultid="3397" heatid="7302" lane="8" entrytime="00:19:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                    <SPLIT distance="200" swimtime="00:02:26.66" />
                    <SPLIT distance="250" swimtime="00:03:05.48" />
                    <SPLIT distance="300" swimtime="00:03:44.60" />
                    <SPLIT distance="350" swimtime="00:04:24.52" />
                    <SPLIT distance="450" swimtime="00:05:44.38" />
                    <SPLIT distance="500" swimtime="00:06:24.82" />
                    <SPLIT distance="550" swimtime="00:07:05.15" />
                    <SPLIT distance="600" swimtime="00:07:46.21" />
                    <SPLIT distance="650" swimtime="00:08:27.29" />
                    <SPLIT distance="700" swimtime="00:09:08.71" />
                    <SPLIT distance="750" swimtime="00:09:50.88" />
                    <SPLIT distance="800" swimtime="00:10:32.47" />
                    <SPLIT distance="850" swimtime="00:11:14.36" />
                    <SPLIT distance="900" swimtime="00:11:56.39" />
                    <SPLIT distance="950" swimtime="00:12:37.51" />
                    <SPLIT distance="1000" swimtime="00:13:19.71" />
                    <SPLIT distance="1050" swimtime="00:14:02.00" />
                    <SPLIT distance="1100" swimtime="00:14:43.96" />
                    <SPLIT distance="1150" swimtime="00:15:26.37" />
                    <SPLIT distance="1200" swimtime="00:16:08.24" />
                    <SPLIT distance="1250" swimtime="00:16:49.54" />
                    <SPLIT distance="1300" swimtime="00:17:30.88" />
                    <SPLIT distance="1350" swimtime="00:18:13.12" />
                    <SPLIT distance="1400" swimtime="00:18:55.13" />
                    <SPLIT distance="1450" swimtime="00:19:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="390" reactiontime="+83" swimtime="00:01:01.46" resultid="3398" heatid="7361" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="338" reactiontime="+96" swimtime="00:01:12.11" resultid="3399" heatid="7386" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="290" reactiontime="+81" swimtime="00:01:13.82" resultid="3400" heatid="7465" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="382" reactiontime="+95" swimtime="00:02:16.86" resultid="3401" heatid="7484" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="150" swimtime="00:01:41.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="3402" heatid="7535" lane="8" entrytime="00:02:30.00" />
                <RESULT eventid="1737" points="372" reactiontime="+89" swimtime="00:04:55.12" resultid="3403" heatid="7576" lane="4" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:46.50" />
                    <SPLIT distance="200" swimtime="00:02:24.84" />
                    <SPLIT distance="250" swimtime="00:03:03.29" />
                    <SPLIT distance="300" swimtime="00:03:42.07" />
                    <SPLIT distance="350" swimtime="00:04:19.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-12-02" firstname="Krzysztof" gender="M" lastname="Drózd" nation="POL" athleteid="2334">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2335" heatid="7261" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2336" heatid="7322" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="2337" heatid="7381" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="1417" status="DNS" swimtime="00:00:00.00" resultid="2338" heatid="7414" lane="4" />
                <RESULT eventid="1481" status="DNS" swimtime="00:00:00.00" resultid="2339" heatid="7464" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="2340" heatid="7533" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="2341" heatid="7546" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-03" firstname="Jarosław" gender="M" lastname="Klonowski" nation="POL" athleteid="4907">
              <RESULTS>
                <RESULT eventid="1076" points="242" reactiontime="+59" swimtime="00:00:32.51" resultid="4908" heatid="7255" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1288" points="234" reactiontime="+76" swimtime="00:01:12.90" resultid="4909" heatid="7355" lane="2" entrytime="00:01:12.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="167" swimtime="00:03:00.30" resultid="4910" heatid="7479" lane="2" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:17.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Krzysztof" gender="M" lastname="Kolibczyński" nation="POL" athleteid="2023">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2024" heatid="7260" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="2025" heatid="7361" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="1449" status="DNS" swimtime="00:00:00.00" resultid="2026" heatid="7445" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-21" firstname="Małgorzata" gender="F" lastname="Osmola" nation="POL" athleteid="3327">
              <RESULTS>
                <RESULT eventid="1059" points="387" reactiontime="+93" swimtime="00:00:31.45" resultid="3328" heatid="7241" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1140" points="321" reactiontime="+90" swimtime="00:11:39.61" resultid="3329" heatid="7291" lane="3" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                    <SPLIT distance="200" swimtime="00:02:41.31" />
                    <SPLIT distance="250" swimtime="00:03:24.72" />
                    <SPLIT distance="300" swimtime="00:04:09.05" />
                    <SPLIT distance="350" swimtime="00:04:53.34" />
                    <SPLIT distance="400" swimtime="00:05:38.20" />
                    <SPLIT distance="450" swimtime="00:06:23.78" />
                    <SPLIT distance="500" swimtime="00:07:09.48" />
                    <SPLIT distance="550" swimtime="00:07:54.79" />
                    <SPLIT distance="600" swimtime="00:08:40.15" />
                    <SPLIT distance="650" swimtime="00:09:25.65" />
                    <SPLIT distance="700" swimtime="00:10:11.85" />
                    <SPLIT distance="750" swimtime="00:10:56.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1207" status="DNS" swimtime="00:00:00.00" resultid="3330" heatid="7312" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1272" points="373" reactiontime="+89" swimtime="00:01:09.79" resultid="3331" heatid="7347" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="3332" heatid="7430" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1497" status="DNS" swimtime="00:00:00.00" resultid="3333" heatid="7473" lane="6" entrytime="00:02:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-05" firstname="Przemysław" gender="M" lastname="Pilarski" nation="POL" athleteid="5825">
              <RESULTS>
                <RESULT eventid="1076" points="112" reactiontime="+99" swimtime="00:00:42.00" resultid="5826" heatid="7260" lane="1" entrytime="00:00:28.58" />
                <RESULT eventid="1108" points="70" swimtime="00:04:25.68" resultid="5827" heatid="7282" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.08" />
                    <SPLIT distance="100" swimtime="00:02:17.38" />
                    <SPLIT distance="150" swimtime="00:03:22.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="77" reactiontime="+98" swimtime="00:00:52.16" resultid="5828" heatid="7323" lane="3" entrytime="00:00:33.40" />
                <RESULT eventid="1256" points="100" swimtime="00:04:18.14" resultid="5829" heatid="7335" lane="6" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.88" />
                    <SPLIT distance="100" swimtime="00:02:06.33" />
                    <SPLIT distance="150" swimtime="00:03:14.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="98" reactiontime="+93" swimtime="00:02:00.23" resultid="5830" heatid="7418" lane="2" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1481" points="56" reactiontime="+93" swimtime="00:02:07.75" resultid="5831" heatid="7463" lane="3" entrytime="00:01:21.00" />
                <RESULT eventid="1657" status="DNS" swimtime="00:00:00.00" resultid="5832" heatid="7533" lane="3" entrytime="00:02:46.00" />
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5833" heatid="7557" lane="2" entrytime="00:00:35.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-14" firstname="Mateusz" gender="M" lastname="Szot" nation="POL" athleteid="5741">
              <RESULTS>
                <RESULT eventid="1256" points="441" reactiontime="+72" swimtime="00:02:37.79" resultid="5742" heatid="7338" lane="6" entrytime="00:02:45.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="527" reactiontime="+77" swimtime="00:01:08.83" resultid="5743" heatid="7425" lane="8" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" status="DNS" swimtime="00:00:00.00" resultid="5744" heatid="7561" lane="0" entrytime="00:00:30.22" />
                <RESULT eventid="1737" status="DNS" swimtime="00:00:00.00" resultid="5745" heatid="7577" lane="4" entrytime="00:05:10.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-04-28" firstname="Andrzej" gender="M" lastname="Wiśniewski" nation="POL" athleteid="6495">
              <RESULTS>
                <RESULT eventid="1188" status="WDR" swimtime="00:00:00.00" resultid="6496" heatid="7305" lane="3" entrytime="00:40:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka " nation="POL" athleteid="6483">
              <RESULTS>
                <RESULT eventid="1092" points="212" reactiontime="+87" swimtime="00:03:24.16" resultid="6484" heatid="7272" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                    <SPLIT distance="100" swimtime="00:01:37.40" />
                    <SPLIT distance="150" swimtime="00:02:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="240" reactiontime="+90" swimtime="00:01:30.90" resultid="6485" heatid="7371" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1400" points="248" reactiontime="+84" swimtime="00:01:39.16" resultid="6486" heatid="7411" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="228" reactiontime="+83" swimtime="00:00:39.87" resultid="6487" heatid="7428" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1673" points="259" reactiontime="+84" swimtime="00:00:44.80" resultid="6488" heatid="7541" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KUPI" nation="SVK" region="BAO" clubid="2791" name="ŠPK Kúpele Piešťany ">
          <ATHLETES>
            <ATHLETE birthdate="1972-04-03" firstname="Juraj" gender="M" lastname="Horii" nation="SVK" license="SVK14912" athleteid="2807">
              <RESULTS>
                <RESULT eventid="1513" points="244" reactiontime="+78" swimtime="00:02:38.95" resultid="2808" heatid="7479" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="215" reactiontime="+81" swimtime="00:12:19.80" resultid="2809" heatid="7297" lane="1" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:58.95" />
                    <SPLIT distance="200" swimtime="00:02:43.86" />
                    <SPLIT distance="250" swimtime="00:03:29.66" />
                    <SPLIT distance="300" swimtime="00:04:16.47" />
                    <SPLIT distance="350" swimtime="00:05:03.47" />
                    <SPLIT distance="400" swimtime="00:05:51.04" />
                    <SPLIT distance="450" swimtime="00:06:38.16" />
                    <SPLIT distance="500" swimtime="00:07:26.19" />
                    <SPLIT distance="550" swimtime="00:08:15.50" />
                    <SPLIT distance="600" swimtime="00:09:04.08" />
                    <SPLIT distance="650" swimtime="00:09:52.51" />
                    <SPLIT distance="700" swimtime="00:10:41.95" />
                    <SPLIT distance="750" swimtime="00:11:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1689" points="341" reactiontime="+81" swimtime="00:00:36.12" resultid="2810" heatid="7556" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="1417" points="327" reactiontime="+78" swimtime="00:01:20.64" resultid="2811" heatid="7421" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="289" reactiontime="+78" swimtime="00:03:01.68" resultid="2812" heatid="7337" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:13.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="256" reactiontime="+84" swimtime="00:01:19.10" resultid="2813" heatid="7382" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-15" firstname="Lucia" gender="F" lastname="Ivicová" nation="SVK" license="SVK10033" athleteid="2823">
              <RESULTS>
                <RESULT eventid="1207" points="396" reactiontime="+78" swimtime="00:00:34.93" resultid="2824" heatid="7312" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1465" points="372" reactiontime="+78" swimtime="00:01:16.49" resultid="2825" heatid="7457" lane="8" entrytime="00:01:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="383" reactiontime="+72" swimtime="00:02:44.16" resultid="2826" heatid="7527" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="428" swimtime="00:00:30.41" resultid="2827" heatid="7243" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1272" points="428" reactiontime="+78" swimtime="00:01:06.67" resultid="2828" heatid="7346" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1497" points="436" reactiontime="+76" swimtime="00:02:25.60" resultid="2829" heatid="7472" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="410" reactiontime="+80" swimtime="00:05:14.71" resultid="2830" heatid="7567" lane="1" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:52.45" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="250" swimtime="00:03:12.43" />
                    <SPLIT distance="300" swimtime="00:03:53.56" />
                    <SPLIT distance="350" swimtime="00:04:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="379" swimtime="00:11:02.06" resultid="2831" heatid="7290" lane="0" entrytime="00:11:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:13.33" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                    <SPLIT distance="200" swimtime="00:02:34.41" />
                    <SPLIT distance="250" swimtime="00:03:16.17" />
                    <SPLIT distance="300" swimtime="00:03:58.52" />
                    <SPLIT distance="350" swimtime="00:04:40.67" />
                    <SPLIT distance="400" swimtime="00:05:23.03" />
                    <SPLIT distance="450" swimtime="00:06:05.63" />
                    <SPLIT distance="500" swimtime="00:06:48.12" />
                    <SPLIT distance="550" swimtime="00:07:30.50" />
                    <SPLIT distance="600" swimtime="00:08:13.37" />
                    <SPLIT distance="650" swimtime="00:08:55.89" />
                    <SPLIT distance="700" swimtime="00:09:38.59" />
                    <SPLIT distance="750" swimtime="00:10:20.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-20" firstname="Anna" gender="F" lastname="Kičínová" nation="SVK" license="SVK13974" athleteid="2790">
              <RESULTS>
                <RESULT eventid="1673" points="294" reactiontime="+77" swimtime="00:00:42.94" resultid="2792" heatid="7542" lane="1" entrytime="00:00:43.70" />
                <RESULT eventid="1400" points="298" reactiontime="+89" swimtime="00:01:33.28" resultid="2793" heatid="7411" lane="4" entrytime="00:01:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="267" reactiontime="+95" swimtime="00:03:28.92" resultid="2794" heatid="7330" lane="6" entrytime="00:03:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:36.19" />
                    <SPLIT distance="150" swimtime="00:02:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="235" reactiontime="+80" swimtime="00:00:39.48" resultid="2795" heatid="7429" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1608" points="248" reactiontime="+83" swimtime="00:01:26.87" resultid="2796" heatid="7509" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="203" reactiontime="+95" swimtime="00:03:23.39" resultid="2797" heatid="7393" lane="8" entrytime="00:03:13.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="150" swimtime="00:02:23.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="242" reactiontime="+96" swimtime="00:03:15.36" resultid="2798" heatid="7273" lane="0" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:34.22" />
                    <SPLIT distance="150" swimtime="00:02:26.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-12" firstname="Zuzanna" gender="F" lastname="Matúšová" nation="SVK" license="SVK21695" athleteid="2814">
              <RESULTS>
                <RESULT eventid="1059" points="446" swimtime="00:00:30.01" resultid="2815" heatid="7244" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1272" points="439" reactiontime="+82" swimtime="00:01:06.08" resultid="2816" heatid="7347" lane="9" entrytime="00:01:07.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="415" reactiontime="+79" swimtime="00:00:32.66" resultid="2817" heatid="7433" lane="2" entrytime="00:00:31.10" />
                <RESULT eventid="1608" points="406" reactiontime="+83" swimtime="00:01:13.70" resultid="2818" heatid="7510" lane="5" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1673" points="474" reactiontime="+81" swimtime="00:00:36.62" resultid="2819" heatid="7544" lane="6" entrytime="00:00:37.60" />
                <RESULT eventid="1400" points="420" reactiontime="+81" swimtime="00:01:23.27" resultid="2820" heatid="7413" lane="9" entrytime="00:01:26.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="427" reactiontime="+81" swimtime="00:01:14.99" resultid="2821" heatid="7375" lane="9" entrytime="00:01:15.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="414" reactiontime="+80" swimtime="00:02:43.47" resultid="2822" heatid="7275" lane="8" entrytime="00:02:43.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:06.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol" gender="M" lastname="Škodný" nation="SVK" license="SVK12519" athleteid="2799">
              <RESULTS>
                <RESULT eventid="1224" points="277" reactiontime="+78" swimtime="00:00:34.06" resultid="2800" heatid="7323" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1481" points="294" reactiontime="+78" swimtime="00:01:13.49" resultid="2801" heatid="7465" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1657" points="312" reactiontime="+75" swimtime="00:02:35.68" resultid="2802" heatid="7534" lane="6" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="368" reactiontime="+86" swimtime="00:02:32.90" resultid="2803" heatid="7282" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1577" points="336" reactiontime="+94" swimtime="00:05:38.43" resultid="2804" heatid="8157" lane="3" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                    <SPLIT distance="150" swimtime="00:02:01.04" />
                    <SPLIT distance="200" swimtime="00:02:43.23" />
                    <SPLIT distance="250" swimtime="00:03:31.98" />
                    <SPLIT distance="300" swimtime="00:04:21.58" />
                    <SPLIT distance="350" swimtime="00:05:01.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1352" points="265" swimtime="00:02:48.51" resultid="2805" heatid="7397" lane="0" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="343" reactiontime="+95" swimtime="00:10:33.39" resultid="2806" heatid="7296" lane="5" entrytime="00:11:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="150" swimtime="00:01:51.53" />
                    <SPLIT distance="200" swimtime="00:02:31.20" />
                    <SPLIT distance="250" swimtime="00:03:11.68" />
                    <SPLIT distance="300" swimtime="00:03:52.26" />
                    <SPLIT distance="350" swimtime="00:04:33.73" />
                    <SPLIT distance="400" swimtime="00:05:15.01" />
                    <SPLIT distance="450" swimtime="00:05:55.96" />
                    <SPLIT distance="500" swimtime="00:06:36.89" />
                    <SPLIT distance="550" swimtime="00:07:17.53" />
                    <SPLIT distance="600" swimtime="00:07:57.99" />
                    <SPLIT distance="650" swimtime="00:08:37.24" />
                    <SPLIT distance="700" swimtime="00:09:17.69" />
                    <SPLIT distance="750" swimtime="00:09:56.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1124" points="413" reactiontime="+80" swimtime="00:01:58.00" resultid="2832" heatid="7288" lane="5" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:00.42" />
                    <SPLIT distance="150" swimtime="00:01:30.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2814" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2823" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2807" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2799" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1705" points="398" reactiontime="+81" swimtime="00:02:11.00" resultid="2833" heatid="7564" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:10.94" />
                    <SPLIT distance="150" swimtime="00:01:43.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2823" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2807" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2814" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2799" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1884" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria A" type="MINIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:45.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1886" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria A" type="MINIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:22:15.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1890" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria B" type="MINIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:15.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1892" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria B" type="MINIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1896" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria C" type="MINIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:21:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1898" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria C" type="MINIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:24:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1902" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria D" type="MINIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:22:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1904" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria D" type="MINIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:26:15.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1908" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria E" type="MINIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:24:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1910" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria E" type="MINIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:28:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1914" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria F" type="MINIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:25:15.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1916" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria F" type="MINIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:30:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1920" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria G" type="MINIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:26:45.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1922" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria G" type="MINIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:33:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1926" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria H" type="MINIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:28:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1928" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria H" type="MINIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:35:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1932" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria I" type="MINIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:29:45.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1934" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria I" type="MINIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:32:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1938" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria J" type="MINIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:32:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1940" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria J" type="MINIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:41:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1944" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria K" type="MINIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:36:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1946" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria K" type="MINIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:44:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1950" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria L" type="MINIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:48:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1952" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria L" type="MINIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:45:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1956" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria M" type="MINIMUM">
      <AGEGROUP agemax="90" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:50:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1958" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria M" type="MINIMUM">
      <AGEGROUP agemax="90" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:45:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1962" course="SCM" gender="M" name="Minikum Startowe 1500m Kategoria N" type="MINIMUM">
      <AGEGROUP agemax="94" agemin="91" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:50:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1964" course="SCM" gender="F" name="Minikum Startowe 1500m Kategoria N" type="MINIMUM">
      <AGEGROUP agemax="94" agemin="91" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:45:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1761" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria A" type="MINIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:10:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1763" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria A" type="MINIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:12:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1773" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria B" type="MINIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:11:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1775" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria B" type="MINIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1779" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria C" type="MINIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:11:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1781" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria C" type="MINIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1785" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria D" type="MINIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1787" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria D" type="MINIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1791" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria E" type="MINIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:13:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1793" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria E" type="MINIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1797" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria F" type="MINIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1799" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria F" type="MINIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1803" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria G" type="MINIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:14:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1805" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria G" type="MINIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1809" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria H" type="MINIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:15:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1811" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria H" type="MINIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1815" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria I" type="MINIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:16:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1817" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria I" type="MINIMUM">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:18:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1821" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria J" type="MINIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:18:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1823" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria J" type="MINIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1827" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria K" type="MINIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:19:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1829" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria K" type="MINIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:22:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1833" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria L" type="MINIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:22:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1835" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria L" type="MINIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:25:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1839" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria M" type="MINIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:23:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1841" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria M" type="MINIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:28:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1845" course="SCM" gender="M" name="Minikum Startowe 800m Kategoria N" type="MINIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:25:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1847" course="SCM" gender="F" name="Minikum Startowe 800m Kategoria N" type="MINIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:30:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>

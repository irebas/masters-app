<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Miejski Klub Plywacki" version="11.56278">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Olsztyn" name="Zimowe Mistrzostwa Polski w Pływaniu w kategoriach Masters, Puchar Polski" course="SCM" deadline="2018-11-07" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2018-11-16" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Olsztyn" nation="POL" />
      <POINTTABLE pointtableid="1122" name="DSV Master Performance Table" version="2016" />
      <SESSIONS>
        <SESSION date="2018-11-16" daytime="14:00" endtime="20:27" name="I Blok" number="1" warmupfrom="12:40" warmupuntil="13:40">
          <EVENTS>
            <EVENT eventid="1150" daytime="17:13" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15091" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15092" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10378" />
                    <RANKING order="2" place="2" resultid="12850" />
                    <RANKING order="3" place="3" resultid="11140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15093" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9170" />
                    <RANKING order="2" place="2" resultid="12089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15094" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10722" />
                    <RANKING order="2" place="2" resultid="12024" />
                    <RANKING order="3" place="3" resultid="10556" />
                    <RANKING order="4" place="-1" resultid="10010" />
                    <RANKING order="5" place="-1" resultid="12002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15095" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12834" />
                    <RANKING order="2" place="2" resultid="11338" />
                    <RANKING order="3" place="3" resultid="10566" />
                    <RANKING order="4" place="4" resultid="9619" />
                    <RANKING order="5" place="5" resultid="10994" />
                    <RANKING order="6" place="6" resultid="11896" />
                    <RANKING order="7" place="7" resultid="10048" />
                    <RANKING order="8" place="8" resultid="12871" />
                    <RANKING order="9" place="9" resultid="11148" />
                    <RANKING order="10" place="-1" resultid="10924" />
                    <RANKING order="11" place="-1" resultid="11870" />
                    <RANKING order="12" place="-1" resultid="12448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15096" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8943" />
                    <RANKING order="2" place="2" resultid="9057" />
                    <RANKING order="3" place="3" resultid="12842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15097" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8936" />
                    <RANKING order="2" place="2" resultid="11926" />
                    <RANKING order="3" place="3" resultid="11209" />
                    <RANKING order="4" place="4" resultid="11774" />
                    <RANKING order="5" place="5" resultid="11909" />
                    <RANKING order="6" place="6" resultid="10641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15098" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12863" />
                    <RANKING order="2" place="2" resultid="11766" />
                    <RANKING order="3" place="3" resultid="9088" />
                    <RANKING order="4" place="4" resultid="11955" />
                    <RANKING order="5" place="5" resultid="11292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15099" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9885" />
                    <RANKING order="2" place="2" resultid="10634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15100" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10353" />
                    <RANKING order="2" place="2" resultid="10627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15101" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9708" />
                    <RANKING order="2" place="2" resultid="12790" />
                    <RANKING order="3" place="3" resultid="10251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15102" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11156" />
                    <RANKING order="2" place="-1" resultid="8882" />
                    <RANKING order="3" place="-1" resultid="11811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15103" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15104" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15105" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14182" daytime="17:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14183" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14184" daytime="17:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14185" daytime="17:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14186" daytime="18:06" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1090" daytime="14:49" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15046" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11916" />
                    <RANKING order="2" place="2" resultid="12082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15047" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9337" />
                    <RANKING order="2" place="2" resultid="9193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15048" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9208" />
                    <RANKING order="2" place="2" resultid="10400" />
                    <RANKING order="3" place="3" resultid="8950" />
                    <RANKING order="4" place="4" resultid="11829" />
                    <RANKING order="5" place="5" resultid="11309" />
                    <RANKING order="6" place="6" resultid="10392" />
                    <RANKING order="7" place="-1" resultid="12438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15049" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9065" />
                    <RANKING order="2" place="2" resultid="12825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15050" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11033" />
                    <RANKING order="2" place="2" resultid="11003" />
                    <RANKING order="3" place="3" resultid="9261" />
                    <RANKING order="4" place="4" resultid="10466" />
                    <RANKING order="5" place="-1" resultid="12464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15051" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9897" />
                    <RANKING order="2" place="2" resultid="9586" />
                    <RANKING order="3" place="3" resultid="13283" />
                    <RANKING order="4" place="4" resultid="11226" />
                    <RANKING order="5" place="5" resultid="11843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15052" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9603" />
                    <RANKING order="2" place="2" resultid="11705" />
                    <RANKING order="3" place="3" resultid="12780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15053" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12045" />
                    <RANKING order="2" place="2" resultid="9049" />
                    <RANKING order="3" place="3" resultid="11981" />
                    <RANKING order="4" place="-1" resultid="11054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15054" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11410" />
                    <RANKING order="2" place="2" resultid="9329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15055" agemax="69" agemin="65" name="65-69" />
                <AGEGROUP agegroupid="15056" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15057" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15058" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15059" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15060" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14162" daytime="14:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14163" daytime="14:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14164" daytime="15:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14165" daytime="15:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="14:16" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15031" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10322" />
                    <RANKING order="2" place="2" resultid="8973" />
                    <RANKING order="3" place="3" resultid="10792" />
                    <RANKING order="4" place="4" resultid="10592" />
                    <RANKING order="5" place="5" resultid="10772" />
                    <RANKING order="6" place="6" resultid="10942" />
                    <RANKING order="7" place="7" resultid="9655" />
                    <RANKING order="8" place="8" resultid="8985" />
                    <RANKING order="9" place="9" resultid="9358" />
                    <RANKING order="10" place="10" resultid="8921" />
                    <RANKING order="11" place="11" resultid="12883" />
                    <RANKING order="12" place="12" resultid="10342" />
                    <RANKING order="13" place="13" resultid="8967" />
                    <RANKING order="14" place="14" resultid="10751" />
                    <RANKING order="15" place="15" resultid="10763" />
                    <RANKING order="16" place="16" resultid="9115" />
                    <RANKING order="17" place="17" resultid="10736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15032" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9474" />
                    <RANKING order="2" place="2" resultid="9027" />
                    <RANKING order="3" place="3" resultid="9151" />
                    <RANKING order="4" place="4" resultid="12919" />
                    <RANKING order="5" place="5" resultid="9145" />
                    <RANKING order="6" place="6" resultid="10947" />
                    <RANKING order="7" place="7" resultid="12017" />
                    <RANKING order="8" place="8" resultid="9105" />
                    <RANKING order="9" place="9" resultid="11321" />
                    <RANKING order="10" place="10" resultid="10798" />
                    <RANKING order="11" place="11" resultid="10803" />
                    <RANKING order="12" place="12" resultid="9368" />
                    <RANKING order="13" place="13" resultid="10755" />
                    <RANKING order="14" place="14" resultid="10759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15033" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9824" />
                    <RANKING order="2" place="2" resultid="9418" />
                    <RANKING order="3" place="3" resultid="9142" />
                    <RANKING order="4" place="4" resultid="10286" />
                    <RANKING order="5" place="5" resultid="9133" />
                    <RANKING order="6" place="6" resultid="10295" />
                    <RANKING order="7" place="7" resultid="9176" />
                    <RANKING order="8" place="8" resultid="10281" />
                    <RANKING order="9" place="9" resultid="9917" />
                    <RANKING order="10" place="10" resultid="9479" />
                    <RANKING order="11" place="11" resultid="10728" />
                    <RANKING order="12" place="12" resultid="9313" />
                    <RANKING order="13" place="13" resultid="10069" />
                    <RANKING order="14" place="14" resultid="9169" />
                    <RANKING order="15" place="15" resultid="10931" />
                    <RANKING order="16" place="16" resultid="10373" />
                    <RANKING order="17" place="17" resultid="11075" />
                    <RANKING order="18" place="18" resultid="9180" />
                    <RANKING order="19" place="19" resultid="9819" />
                    <RANKING order="20" place="20" resultid="9272" />
                    <RANKING order="21" place="21" resultid="12088" />
                    <RANKING order="22" place="-1" resultid="9178" />
                    <RANKING order="23" place="-1" resultid="9569" />
                    <RANKING order="24" place="-1" resultid="9955" />
                    <RANKING order="25" place="-1" resultid="10548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15034" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10302" />
                    <RANKING order="2" place="2" resultid="11303" />
                    <RANKING order="3" place="3" resultid="11046" />
                    <RANKING order="4" place="4" resultid="9902" />
                    <RANKING order="5" place="5" resultid="12075" />
                    <RANKING order="6" place="6" resultid="11942" />
                    <RANKING order="7" place="7" resultid="9751" />
                    <RANKING order="8" place="8" resultid="9138" />
                    <RANKING order="9" place="9" resultid="9973" />
                    <RANKING order="10" place="10" resultid="10365" />
                    <RANKING order="11" place="11" resultid="11249" />
                    <RANKING order="12" place="11" resultid="12857" />
                    <RANKING order="13" place="13" resultid="10039" />
                    <RANKING order="14" place="14" resultid="11118" />
                    <RANKING order="15" place="15" resultid="10009" />
                    <RANKING order="16" place="16" resultid="10062" />
                    <RANKING order="17" place="17" resultid="10016" />
                    <RANKING order="18" place="18" resultid="12805" />
                    <RANKING order="19" place="19" resultid="10969" />
                    <RANKING order="20" place="19" resultid="11235" />
                    <RANKING order="21" place="21" resultid="10937" />
                    <RANKING order="22" place="22" resultid="10424" />
                    <RANKING order="23" place="23" resultid="10024" />
                    <RANKING order="24" place="24" resultid="9424" />
                    <RANKING order="25" place="25" resultid="10076" />
                    <RANKING order="26" place="26" resultid="9965" />
                    <RANKING order="27" place="27" resultid="9015" />
                    <RANKING order="28" place="-1" resultid="11136" />
                    <RANKING order="29" place="-1" resultid="8867" />
                    <RANKING order="30" place="-1" resultid="9186" />
                    <RANKING order="31" place="-1" resultid="10054" />
                    <RANKING order="32" place="-1" resultid="10555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15035" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9155" />
                    <RANKING order="2" place="2" resultid="10565" />
                    <RANKING order="3" place="3" resultid="11933" />
                    <RANKING order="4" place="4" resultid="10988" />
                    <RANKING order="5" place="5" resultid="10242" />
                    <RANKING order="6" place="6" resultid="9611" />
                    <RANKING order="7" place="7" resultid="9987" />
                    <RANKING order="8" place="8" resultid="9795" />
                    <RANKING order="9" place="9" resultid="11950" />
                    <RANKING order="10" place="10" resultid="9444" />
                    <RANKING order="11" place="11" resultid="11337" />
                    <RANKING order="12" place="12" resultid="12844" />
                    <RANKING order="13" place="13" resultid="11895" />
                    <RANKING order="14" place="14" resultid="11869" />
                    <RANKING order="15" place="15" resultid="11112" />
                    <RANKING order="16" place="16" resultid="12447" />
                    <RANKING order="17" place="17" resultid="10047" />
                    <RANKING order="18" place="18" resultid="12102" />
                    <RANKING order="19" place="19" resultid="10993" />
                    <RANKING order="20" place="20" resultid="11278" />
                    <RANKING order="21" place="21" resultid="9815" />
                    <RANKING order="22" place="22" resultid="8784" />
                    <RANKING order="23" place="23" resultid="10918" />
                    <RANKING order="24" place="24" resultid="9188" />
                    <RANKING order="25" place="25" resultid="12870" />
                    <RANKING order="26" place="26" resultid="10923" />
                    <RANKING order="27" place="27" resultid="9319" />
                    <RANKING order="28" place="-1" resultid="9996" />
                    <RANKING order="29" place="-1" resultid="9184" />
                    <RANKING order="30" place="-1" resultid="9268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15036" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11387" />
                    <RANKING order="2" place="2" resultid="10572" />
                    <RANKING order="3" place="3" resultid="8913" />
                    <RANKING order="4" place="4" resultid="10472" />
                    <RANKING order="5" place="5" resultid="10831" />
                    <RANKING order="6" place="6" resultid="10823" />
                    <RANKING order="7" place="7" resultid="8897" />
                    <RANKING order="8" place="8" resultid="11884" />
                    <RANKING order="9" place="9" resultid="11364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15037" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10726" />
                    <RANKING order="2" place="2" resultid="12423" />
                    <RANKING order="3" place="3" resultid="11282" />
                    <RANKING order="4" place="4" resultid="11784" />
                    <RANKING order="5" place="5" resultid="11925" />
                    <RANKING order="6" place="6" resultid="9949" />
                    <RANKING order="7" place="7" resultid="11208" />
                    <RANKING order="8" place="8" resultid="11805" />
                    <RANKING order="9" place="9" resultid="8844" />
                    <RANKING order="10" place="10" resultid="11773" />
                    <RANKING order="11" place="11" resultid="11072" />
                    <RANKING order="12" place="12" resultid="9392" />
                    <RANKING order="13" place="13" resultid="9428" />
                    <RANKING order="14" place="14" resultid="11890" />
                    <RANKING order="15" place="-1" resultid="9845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15038" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9034" />
                    <RANKING order="2" place="2" resultid="9802" />
                    <RANKING order="3" place="3" resultid="11078" />
                    <RANKING order="4" place="4" resultid="11765" />
                    <RANKING order="5" place="5" resultid="11197" />
                    <RANKING order="6" place="6" resultid="9399" />
                    <RANKING order="7" place="7" resultid="9087" />
                    <RANKING order="8" place="8" resultid="11291" />
                    <RANKING order="9" place="-1" resultid="11759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15039" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12815" />
                    <RANKING order="2" place="2" resultid="10542" />
                    <RANKING order="3" place="3" resultid="11202" />
                    <RANKING order="4" place="4" resultid="9123" />
                    <RANKING order="5" place="5" resultid="11754" />
                    <RANKING order="6" place="6" resultid="10347" />
                    <RANKING order="7" place="7" resultid="10877" />
                    <RANKING order="8" place="8" resultid="9851" />
                    <RANKING order="9" place="9" resultid="9411" />
                    <RANKING order="10" place="10" resultid="9690" />
                    <RANKING order="11" place="11" resultid="9839" />
                    <RANKING order="12" place="-1" resultid="12387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15040" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11257" />
                    <RANKING order="2" place="2" resultid="11746" />
                    <RANKING order="3" place="3" resultid="11393" />
                    <RANKING order="4" place="4" resultid="9531" />
                    <RANKING order="5" place="4" resultid="10352" />
                    <RANKING order="6" place="6" resultid="11741" />
                    <RANKING order="7" place="7" resultid="10448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15041" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9920" />
                    <RANKING order="2" place="2" resultid="8792" />
                    <RANKING order="3" place="3" resultid="10500" />
                    <RANKING order="4" place="4" resultid="12789" />
                    <RANKING order="5" place="5" resultid="9535" />
                    <RANKING order="6" place="6" resultid="8818" />
                    <RANKING order="7" place="-1" resultid="8862" />
                    <RANKING order="8" place="-1" resultid="10441" />
                    <RANKING order="9" place="-1" resultid="11735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15042" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10889" />
                    <RANKING order="2" place="2" resultid="11155" />
                    <RANKING order="3" place="3" resultid="10435" />
                    <RANKING order="4" place="4" resultid="10528" />
                    <RANKING order="5" place="5" resultid="9745" />
                    <RANKING order="6" place="6" resultid="11810" />
                    <RANKING order="7" place="7" resultid="8827" />
                    <RANKING order="8" place="8" resultid="8810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15043" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11380" />
                    <RANKING order="2" place="2" resultid="10430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15044" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9305" />
                    <RANKING order="2" place="2" resultid="9302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15045" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14142" daytime="14:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14143" daytime="14:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14144" daytime="14:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14145" daytime="14:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14146" daytime="14:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14147" daytime="14:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14148" daytime="14:27" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14149" daytime="14:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14150" daytime="14:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14151" daytime="14:31" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14152" daytime="14:33" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14153" daytime="14:34" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14154" daytime="14:36" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14155" daytime="14:37" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14156" daytime="14:39" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14157" daytime="14:40" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="14158" daytime="14:42" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="14159" daytime="14:43" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="14160" daytime="14:44" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="14161" daytime="14:46" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="15:11" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15061" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15062" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12764" />
                    <RANKING order="2" place="2" resultid="9648" />
                    <RANKING order="3" place="3" resultid="12849" />
                    <RANKING order="4" place="-1" resultid="11191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15063" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9825" />
                    <RANKING order="2" place="2" resultid="9926" />
                    <RANKING order="3" place="3" resultid="10287" />
                    <RANKING order="4" place="4" resultid="9314" />
                    <RANKING order="5" place="5" resultid="9480" />
                    <RANKING order="6" place="6" resultid="12756" />
                    <RANKING order="7" place="-1" resultid="9372" />
                    <RANKING order="8" place="-1" resultid="10549" />
                    <RANKING order="9" place="-1" resultid="10964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15064" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10303" />
                    <RANKING order="2" place="2" resultid="11943" />
                    <RANKING order="3" place="3" resultid="9979" />
                    <RANKING order="4" place="4" resultid="9903" />
                    <RANKING order="5" place="5" resultid="11250" />
                    <RANKING order="6" place="6" resultid="10366" />
                    <RANKING order="7" place="7" resultid="10385" />
                    <RANKING order="8" place="8" resultid="11236" />
                    <RANKING order="9" place="9" resultid="10360" />
                    <RANKING order="10" place="10" resultid="10017" />
                    <RANKING order="11" place="11" resultid="10036" />
                    <RANKING order="12" place="-1" resultid="10040" />
                    <RANKING order="13" place="-1" resultid="12001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15065" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12833" />
                    <RANKING order="2" place="2" resultid="11934" />
                    <RANKING order="3" place="3" resultid="9988" />
                    <RANKING order="4" place="4" resultid="9161" />
                    <RANKING order="5" place="5" resultid="9618" />
                    <RANKING order="6" place="6" resultid="11862" />
                    <RANKING order="7" place="7" resultid="11122" />
                    <RANKING order="8" place="8" resultid="8785" />
                    <RANKING order="9" place="9" resultid="9320" />
                    <RANKING order="10" place="-1" resultid="11316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15066" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10578" />
                    <RANKING order="2" place="2" resultid="9634" />
                    <RANKING order="3" place="3" resultid="10473" />
                    <RANKING order="4" place="4" resultid="8914" />
                    <RANKING order="5" place="5" resultid="9054" />
                    <RANKING order="6" place="6" resultid="10832" />
                    <RANKING order="7" place="7" resultid="11017" />
                    <RANKING order="8" place="8" resultid="11365" />
                    <RANKING order="9" place="-1" resultid="11011" />
                    <RANKING order="10" place="-1" resultid="8942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15067" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11283" />
                    <RANKING order="2" place="2" resultid="12424" />
                    <RANKING order="3" place="3" resultid="12396" />
                    <RANKING order="4" place="4" resultid="8845" />
                    <RANKING order="5" place="5" resultid="9465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15068" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9035" />
                    <RANKING order="2" place="2" resultid="9963" />
                    <RANKING order="3" place="3" resultid="9803" />
                    <RANKING order="4" place="4" resultid="9594" />
                    <RANKING order="5" place="5" resultid="9737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15069" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12816" />
                    <RANKING order="2" place="2" resultid="8778" />
                    <RANKING order="3" place="3" resultid="9662" />
                    <RANKING order="4" place="4" resultid="9124" />
                    <RANKING order="5" place="5" resultid="10633" />
                    <RANKING order="6" place="6" resultid="11264" />
                    <RANKING order="7" place="7" resultid="9404" />
                    <RANKING order="8" place="8" resultid="9852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15070" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11747" />
                    <RANKING order="2" place="2" resultid="11373" />
                    <RANKING order="3" place="3" resultid="9571" />
                    <RANKING order="4" place="4" resultid="11727" />
                    <RANKING order="5" place="5" resultid="10449" />
                    <RANKING order="6" place="-1" resultid="8835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15071" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10621" />
                    <RANKING order="2" place="2" resultid="9707" />
                    <RANKING order="3" place="3" resultid="11819" />
                    <RANKING order="4" place="4" resultid="10250" />
                    <RANKING order="5" place="5" resultid="8819" />
                    <RANKING order="6" place="6" resultid="8872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15072" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10529" />
                    <RANKING order="2" place="2" resultid="8828" />
                    <RANKING order="3" place="-1" resultid="8881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15073" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15074" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15075" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14166" daytime="15:11" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14167" daytime="15:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14168" daytime="15:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14169" daytime="15:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14170" daytime="15:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14171" daytime="15:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14172" daytime="15:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14173" daytime="15:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14174" daytime="15:47" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="15:53" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="14960" agemax="99" agemin="80" name="80-99" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14961" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12923" />
                    <RANKING order="2" place="2" resultid="11177" />
                    <RANKING order="3" place="-1" resultid="9215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14962" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9216" />
                    <RANKING order="2" place="2" resultid="10312" />
                    <RANKING order="3" place="3" resultid="10080" />
                    <RANKING order="4" place="4" resultid="12112" />
                    <RANKING order="5" place="5" resultid="10456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14963" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9936" />
                    <RANKING order="2" place="2" resultid="9773" />
                    <RANKING order="3" place="3" resultid="12921" />
                    <RANKING order="4" place="4" resultid="11900" />
                    <RANKING order="5" place="5" resultid="11029" />
                    <RANKING order="6" place="6" resultid="12453" />
                    <RANKING order="7" place="7" resultid="11901" />
                    <RANKING order="8" place="8" resultid="12036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14964" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11792" />
                    <RANKING order="2" place="2" resultid="9070" />
                    <RANKING order="3" place="3" resultid="12035" />
                    <RANKING order="4" place="4" resultid="10457" />
                    <RANKING order="5" place="-1" resultid="9938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14965" agemax="279" agemin="240" name="240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9775" />
                    <RANKING order="2" place="2" resultid="10893" />
                    <RANKING order="3" place="-1" resultid="11789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14966" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9554" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14175" daytime="15:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14176" daytime="15:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14177" daytime="16:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1058" daytime="14:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1062" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9382" />
                    <RANKING order="2" place="2" resultid="8980" />
                    <RANKING order="3" place="3" resultid="10739" />
                    <RANKING order="4" place="-1" resultid="10788" />
                    <RANKING order="5" place="-1" resultid="10808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10958" />
                    <RANKING order="2" place="2" resultid="12794" />
                    <RANKING order="3" place="3" resultid="9488" />
                    <RANKING order="4" place="4" resultid="10778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11722" />
                    <RANKING order="2" place="2" resultid="10260" />
                    <RANKING order="3" place="3" resultid="9207" />
                    <RANKING order="4" place="4" resultid="10399" />
                    <RANKING order="5" place="5" resultid="9200" />
                    <RANKING order="6" place="6" resultid="10747" />
                    <RANKING order="7" place="7" resultid="10272" />
                    <RANKING order="8" place="8" resultid="10265" />
                    <RANKING order="9" place="9" resultid="11048" />
                    <RANKING order="10" place="-1" resultid="12110" />
                    <RANKING order="11" place="-1" resultid="12404" />
                    <RANKING order="12" place="-1" resultid="13297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9059" />
                    <RANKING order="2" place="2" resultid="10033" />
                    <RANKING order="3" place="3" resultid="12432" />
                    <RANKING order="4" place="4" resultid="12824" />
                    <RANKING order="5" place="5" resultid="9810" />
                    <RANKING order="6" place="6" resultid="12915" />
                    <RANKING order="7" place="7" resultid="12812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10058" />
                    <RANKING order="2" place="2" resultid="10980" />
                    <RANKING order="3" place="3" resultid="11836" />
                    <RANKING order="4" place="4" resultid="11345" />
                    <RANKING order="5" place="5" resultid="13208" />
                    <RANKING order="6" place="6" resultid="11002" />
                    <RANKING order="7" place="7" resultid="11848" />
                    <RANKING order="8" place="8" resultid="11799" />
                    <RANKING order="9" place="9" resultid="12799" />
                    <RANKING order="10" place="10" resultid="10733" />
                    <RANKING order="11" place="11" resultid="11990" />
                    <RANKING order="12" place="12" resultid="12030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9678" />
                    <RANKING order="2" place="2" resultid="9911" />
                    <RANKING order="3" place="3" resultid="11711" />
                    <RANKING order="4" place="4" resultid="9585" />
                    <RANKING order="5" place="5" resultid="13282" />
                    <RANKING order="6" place="6" resultid="10417" />
                    <RANKING order="7" place="7" resultid="12888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9671" />
                    <RANKING order="2" place="2" resultid="10678" />
                    <RANKING order="3" place="3" resultid="10586" />
                    <RANKING order="4" place="4" resultid="9602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9866" />
                    <RANKING order="2" place="2" resultid="9698" />
                    <RANKING order="3" place="3" resultid="11699" />
                    <RANKING order="4" place="4" resultid="10859" />
                    <RANKING order="5" place="5" resultid="13291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11995" />
                    <RANKING order="2" place="2" resultid="9759" />
                    <RANKING order="3" place="3" resultid="10868" />
                    <RANKING order="4" place="4" resultid="9328" />
                    <RANKING order="5" place="5" resultid="10408" />
                    <RANKING order="6" place="6" resultid="12457" />
                    <RANKING order="7" place="-1" resultid="11693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9499" />
                    <RANKING order="2" place="2" resultid="10523" />
                    <RANKING order="3" place="3" resultid="10646" />
                    <RANKING order="4" place="4" resultid="12010" />
                    <RANKING order="5" place="5" resultid="10884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11360" />
                    <RANKING order="2" place="2" resultid="9550" />
                    <RANKING order="3" place="3" resultid="9716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="2243" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1059" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14134" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14135" daytime="14:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14136" daytime="14:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14137" daytime="14:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14138" daytime="14:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14139" daytime="14:09" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14140" daytime="14:11" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14141" daytime="14:12" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="16:05" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15076" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11917" />
                    <RANKING order="2" place="2" resultid="9383" />
                    <RANKING order="3" place="3" resultid="8995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15077" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15078" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8951" />
                    <RANKING order="2" place="2" resultid="10273" />
                    <RANKING order="3" place="3" resultid="11310" />
                    <RANKING order="4" place="4" resultid="12439" />
                    <RANKING order="5" place="5" resultid="12405" />
                    <RANKING order="6" place="-1" resultid="11049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15079" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15080" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11034" />
                    <RANKING order="2" place="2" resultid="9969" />
                    <RANKING order="3" place="3" resultid="12465" />
                    <RANKING order="4" place="4" resultid="11144" />
                    <RANKING order="5" place="-1" resultid="10027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15081" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9543" />
                    <RANKING order="2" place="2" resultid="11227" />
                    <RANKING order="3" place="3" resultid="10418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15082" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15083" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9699" />
                    <RANKING order="2" place="2" resultid="10860" />
                    <RANKING order="3" place="3" resultid="11982" />
                    <RANKING order="4" place="-1" resultid="11055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15084" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9760" />
                    <RANKING order="2" place="2" resultid="10869" />
                    <RANKING order="3" place="3" resultid="10409" />
                    <RANKING order="4" place="4" resultid="11970" />
                    <RANKING order="5" place="-1" resultid="11062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15085" agemax="69" agemin="65" name="65-69" />
                <AGEGROUP agegroupid="15086" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15087" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15088" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15089" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15090" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14178" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14179" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14180" daytime="16:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14181" daytime="16:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="18:32" gender="F" number="8" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15106" agemax="24" agemin="20" name="20-24" />
                <AGEGROUP agegroupid="15107" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9194" />
                    <RANKING order="2" place="2" resultid="9338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15108" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12895" />
                    <RANKING order="2" place="2" resultid="12068" />
                    <RANKING order="3" place="-1" resultid="10393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15109" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9460" />
                    <RANKING order="2" place="2" resultid="9073" />
                    <RANKING order="3" place="-1" resultid="11129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15110" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10702" />
                    <RANKING order="2" place="-1" resultid="8963" />
                    <RANKING order="3" place="-1" resultid="9768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15111" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15112" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15113" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11854" />
                    <RANKING order="2" place="2" resultid="9725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15114" agemax="64" agemin="60" name="60-64" />
                <AGEGROUP agegroupid="15115" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10647" />
                    <RANKING order="2" place="2" resultid="11298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15116" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15117" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15118" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15119" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15120" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14187" daytime="18:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14188" daytime="18:59" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8179" daytime="19:36" gender="M" number="9" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15121" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9021" />
                    <RANKING order="2" place="2" resultid="9656" />
                    <RANKING order="3" place="3" resultid="9627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15122" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12765" />
                    <RANKING order="2" place="-1" resultid="9493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15123" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9373" />
                    <RANKING order="2" place="2" resultid="10238" />
                    <RANKING order="3" place="-1" resultid="10717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15124" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13279" />
                    <RANKING order="2" place="-1" resultid="12806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15125" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12903" />
                    <RANKING order="2" place="2" resultid="8930" />
                    <RANKING order="3" place="3" resultid="9796" />
                    <RANKING order="4" place="4" resultid="9643" />
                    <RANKING order="5" place="5" resultid="11863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15126" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10697" />
                    <RANKING order="2" place="2" resultid="10824" />
                    <RANKING order="3" place="-1" resultid="11104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15127" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11782" />
                    <RANKING order="2" place="2" resultid="11073" />
                    <RANKING order="3" place="3" resultid="13205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15128" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15129" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12388" />
                    <RANKING order="2" place="2" resultid="12053" />
                    <RANKING order="3" place="3" resultid="9001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15130" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11728" />
                    <RANKING order="2" place="2" resultid="8836" />
                    <RANKING order="3" place="3" resultid="10518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15131" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11820" />
                    <RANKING order="2" place="2" resultid="8793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15132" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15133" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15134" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15135" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14189" daytime="19:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14190" daytime="19:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14191" daytime="20:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14192" daytime="20:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-11-17" daytime="09:00" endtime="13:04" name="II Blok" number="2" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="8245" daytime="09:58" gender="M" number="13" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15181" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9022" />
                    <RANKING order="2" place="2" resultid="8986" />
                    <RANKING order="3" place="3" resultid="10329" />
                    <RANKING order="4" place="4" resultid="10607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15182" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10379" />
                    <RANKING order="2" place="2" resultid="10781" />
                    <RANKING order="3" place="3" resultid="12742" />
                    <RANKING order="4" place="-1" resultid="9452" />
                    <RANKING order="5" place="-1" resultid="9942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15183" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11354" />
                    <RANKING order="2" place="2" resultid="10282" />
                    <RANKING order="3" place="3" resultid="12360" />
                    <RANKING order="4" place="4" resultid="12757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15184" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11944" />
                    <RANKING order="2" place="2" resultid="12858" />
                    <RANKING order="3" place="3" resultid="10041" />
                    <RANKING order="4" place="4" resultid="11877" />
                    <RANKING order="5" place="5" resultid="12417" />
                    <RANKING order="6" place="-1" resultid="10011" />
                    <RANKING order="7" place="-1" resultid="10063" />
                    <RANKING order="8" place="-1" resultid="12003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15185" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9006" />
                    <RANKING order="2" place="2" resultid="11123" />
                    <RANKING order="3" place="-1" resultid="10661" />
                    <RANKING order="4" place="-1" resultid="11978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15186" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11012" />
                    <RANKING order="2" place="2" resultid="8944" />
                    <RANKING order="3" place="3" resultid="11366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15187" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12397" />
                    <RANKING order="2" place="2" resultid="11910" />
                    <RANKING order="3" place="3" resultid="10642" />
                    <RANKING order="4" place="4" resultid="9466" />
                    <RANKING order="5" place="5" resultid="8905" />
                    <RANKING order="6" place="6" resultid="9393" />
                    <RANKING order="7" place="7" resultid="11271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15188" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11198" />
                    <RANKING order="2" place="2" resultid="11767" />
                    <RANKING order="3" place="3" resultid="12864" />
                    <RANKING order="4" place="4" resultid="9738" />
                    <RANKING order="5" place="5" resultid="9881" />
                    <RANKING order="6" place="-1" resultid="12413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15189" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8779" />
                    <RANKING order="2" place="2" resultid="9125" />
                    <RANKING order="3" place="3" resultid="9663" />
                    <RANKING order="4" place="4" resultid="11265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15190" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11748" />
                    <RANKING order="2" place="2" resultid="11374" />
                    <RANKING order="3" place="3" resultid="10513" />
                    <RANKING order="4" place="4" resultid="9572" />
                    <RANKING order="5" place="5" resultid="11742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15191" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9833" />
                    <RANKING order="2" place="2" resultid="11821" />
                    <RANKING order="3" place="3" resultid="10443" />
                    <RANKING order="4" place="4" resultid="10252" />
                    <RANKING order="5" place="5" resultid="8820" />
                    <RANKING order="6" place="6" resultid="8873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15192" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9503" />
                    <RANKING order="2" place="2" resultid="8854" />
                    <RANKING order="3" place="-1" resultid="8883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15193" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15194" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15195" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14212" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14213" daytime="10:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14214" daytime="10:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14215" daytime="10:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14216" daytime="10:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14217" daytime="10:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8277" daytime="10:47" gender="M" number="15" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15211" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10794" />
                    <RANKING order="2" place="2" resultid="8974" />
                    <RANKING order="3" place="3" resultid="10773" />
                    <RANKING order="4" place="4" resultid="9657" />
                    <RANKING order="5" place="5" resultid="10943" />
                    <RANKING order="6" place="6" resultid="8923" />
                    <RANKING order="7" place="7" resultid="9361" />
                    <RANKING order="8" place="8" resultid="12884" />
                    <RANKING order="9" place="9" resultid="10600" />
                    <RANKING order="10" place="10" resultid="10752" />
                    <RANKING order="11" place="11" resultid="10764" />
                    <RANKING order="12" place="12" resultid="10343" />
                    <RANKING order="13" place="13" resultid="8968" />
                    <RANKING order="14" place="14" resultid="9116" />
                    <RANKING order="15" place="-1" resultid="10330" />
                    <RANKING order="16" place="-1" resultid="10594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15212" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9475" />
                    <RANKING order="2" place="2" resultid="12019" />
                    <RANKING order="3" place="3" resultid="11398" />
                    <RANKING order="4" place="4" resultid="9106" />
                    <RANKING order="5" place="5" resultid="12851" />
                    <RANKING order="6" place="6" resultid="9369" />
                    <RANKING order="7" place="7" resultid="11141" />
                    <RANKING order="8" place="8" resultid="10756" />
                    <RANKING order="9" place="9" resultid="10760" />
                    <RANKING order="10" place="-1" resultid="11192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15213" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9826" />
                    <RANKING order="2" place="2" resultid="9134" />
                    <RANKING order="3" place="3" resultid="12365" />
                    <RANKING order="4" place="4" resultid="10296" />
                    <RANKING order="5" place="5" resultid="9481" />
                    <RANKING order="6" place="6" resultid="9172" />
                    <RANKING order="7" place="7" resultid="9315" />
                    <RANKING order="8" place="8" resultid="10718" />
                    <RANKING order="9" place="9" resultid="10932" />
                    <RANKING order="10" place="10" resultid="10070" />
                    <RANKING order="11" place="11" resultid="9821" />
                    <RANKING order="12" place="12" resultid="12090" />
                    <RANKING order="13" place="-1" resultid="9956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15214" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12076" />
                    <RANKING order="2" place="2" resultid="9904" />
                    <RANKING order="3" place="3" resultid="9974" />
                    <RANKING order="4" place="4" resultid="9139" />
                    <RANKING order="5" place="5" resultid="11252" />
                    <RANKING order="6" place="6" resultid="9752" />
                    <RANKING order="7" place="7" resultid="11137" />
                    <RANKING order="8" place="8" resultid="12807" />
                    <RANKING order="9" place="9" resultid="10558" />
                    <RANKING order="10" place="10" resultid="11878" />
                    <RANKING order="11" place="11" resultid="10970" />
                    <RANKING order="12" place="12" resultid="10938" />
                    <RANKING order="13" place="13" resultid="10425" />
                    <RANKING order="14" place="14" resultid="9425" />
                    <RANKING order="15" place="15" resultid="12418" />
                    <RANKING order="16" place="16" resultid="9966" />
                    <RANKING order="17" place="17" resultid="9016" />
                    <RANKING order="18" place="-1" resultid="8868" />
                    <RANKING order="19" place="-1" resultid="10953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15215" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12835" />
                    <RANKING order="2" place="2" resultid="11936" />
                    <RANKING order="3" place="3" resultid="10567" />
                    <RANKING order="4" place="4" resultid="10989" />
                    <RANKING order="5" place="5" resultid="9613" />
                    <RANKING order="6" place="6" resultid="12904" />
                    <RANKING order="7" place="7" resultid="11951" />
                    <RANKING order="8" place="8" resultid="9797" />
                    <RANKING order="9" place="9" resultid="11340" />
                    <RANKING order="10" place="10" resultid="9445" />
                    <RANKING order="11" place="11" resultid="11898" />
                    <RANKING order="12" place="12" resultid="11871" />
                    <RANKING order="13" place="13" resultid="9998" />
                    <RANKING order="14" place="14" resultid="10995" />
                    <RANKING order="15" place="15" resultid="12449" />
                    <RANKING order="16" place="16" resultid="11279" />
                    <RANKING order="17" place="17" resultid="10050" />
                    <RANKING order="18" place="18" resultid="11113" />
                    <RANKING order="19" place="19" resultid="12103" />
                    <RANKING order="20" place="20" resultid="9816" />
                    <RANKING order="21" place="21" resultid="12873" />
                    <RANKING order="22" place="22" resultid="8786" />
                    <RANKING order="23" place="23" resultid="11149" />
                    <RANKING order="24" place="24" resultid="10925" />
                    <RANKING order="25" place="25" resultid="10919" />
                    <RANKING order="26" place="26" resultid="9440" />
                    <RANKING order="27" place="-1" resultid="9989" />
                    <RANKING order="28" place="-1" resultid="11317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15216" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11388" />
                    <RANKING order="2" place="2" resultid="9635" />
                    <RANKING order="3" place="3" resultid="10573" />
                    <RANKING order="4" place="4" resultid="8916" />
                    <RANKING order="5" place="5" resultid="10833" />
                    <RANKING order="6" place="6" resultid="10698" />
                    <RANKING order="7" place="7" resultid="10825" />
                    <RANKING order="8" place="8" resultid="8898" />
                    <RANKING order="9" place="9" resultid="11885" />
                    <RANKING order="10" place="10" resultid="9346" />
                    <RANKING order="11" place="11" resultid="9434" />
                    <RANKING order="12" place="-1" resultid="11105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15217" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8937" />
                    <RANKING order="2" place="2" resultid="12425" />
                    <RANKING order="3" place="3" resultid="11806" />
                    <RANKING order="4" place="4" resultid="11210" />
                    <RANKING order="5" place="5" resultid="11775" />
                    <RANKING order="6" place="6" resultid="8846" />
                    <RANKING order="7" place="7" resultid="12911" />
                    <RANKING order="8" place="8" resultid="9394" />
                    <RANKING order="9" place="9" resultid="11892" />
                    <RANKING order="10" place="-1" resultid="9846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15218" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9961" />
                    <RANKING order="2" place="2" resultid="9036" />
                    <RANKING order="3" place="3" resultid="9805" />
                    <RANKING order="4" place="4" resultid="9595" />
                    <RANKING order="5" place="5" resultid="9527" />
                    <RANKING order="6" place="6" resultid="9400" />
                    <RANKING order="7" place="7" resultid="11293" />
                    <RANKING order="8" place="-1" resultid="11761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15219" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10544" />
                    <RANKING order="2" place="2" resultid="11203" />
                    <RANKING order="3" place="3" resultid="12389" />
                    <RANKING order="4" place="4" resultid="10879" />
                    <RANKING order="5" place="5" resultid="9002" />
                    <RANKING order="6" place="6" resultid="9692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15220" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11259" />
                    <RANKING order="2" place="2" resultid="10354" />
                    <RANKING order="3" place="3" resultid="9351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15221" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9709" />
                    <RANKING order="2" place="2" resultid="9922" />
                    <RANKING order="3" place="3" resultid="8794" />
                    <RANKING order="4" place="-1" resultid="11737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15222" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11158" />
                    <RANKING order="2" place="2" resultid="10890" />
                    <RANKING order="3" place="3" resultid="9747" />
                    <RANKING order="4" place="4" resultid="10437" />
                    <RANKING order="5" place="5" resultid="11813" />
                    <RANKING order="6" place="6" resultid="8812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15223" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15224" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9308" />
                    <RANKING order="2" place="2" resultid="9098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15225" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14224" daytime="10:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14225" daytime="10:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14226" daytime="10:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14227" daytime="10:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14228" daytime="11:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14229" daytime="11:03" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14230" daytime="11:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14231" daytime="11:07" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14232" daytime="11:09" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14233" daytime="11:11" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14234" daytime="11:13" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14235" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14236" daytime="11:17" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14237" daytime="11:19" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8213" daytime="09:12" gender="M" number="11" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15151" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10793" />
                    <RANKING order="2" place="2" resultid="10323" />
                    <RANKING order="3" place="3" resultid="10593" />
                    <RANKING order="4" place="4" resultid="10315" />
                    <RANKING order="5" place="5" resultid="9360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15152" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10948" />
                    <RANKING order="2" place="2" resultid="9494" />
                    <RANKING order="3" place="3" resultid="12018" />
                    <RANKING order="4" place="4" resultid="11322" />
                    <RANKING order="5" place="5" resultid="12741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15153" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10288" />
                    <RANKING order="2" place="2" resultid="11327" />
                    <RANKING order="3" place="3" resultid="12359" />
                    <RANKING order="4" place="4" resultid="10672" />
                    <RANKING order="5" place="5" resultid="9171" />
                    <RANKING order="6" place="6" resultid="9273" />
                    <RANKING order="7" place="7" resultid="9820" />
                    <RANKING order="8" place="-1" resultid="10550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15154" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10304" />
                    <RANKING order="2" place="2" resultid="11304" />
                    <RANKING order="3" place="3" resultid="9874" />
                    <RANKING order="4" place="4" resultid="9980" />
                    <RANKING order="5" place="5" resultid="11251" />
                    <RANKING order="6" place="6" resultid="10367" />
                    <RANKING order="7" place="7" resultid="10386" />
                    <RANKING order="8" place="8" resultid="10557" />
                    <RANKING order="9" place="9" resultid="10025" />
                    <RANKING order="10" place="-1" resultid="10055" />
                    <RANKING order="11" place="-1" resultid="11237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15155" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9156" />
                    <RANKING order="2" place="2" resultid="9612" />
                    <RANKING order="3" place="3" resultid="11935" />
                    <RANKING order="4" place="4" resultid="9280" />
                    <RANKING order="5" place="5" resultid="10243" />
                    <RANKING order="6" place="6" resultid="11897" />
                    <RANKING order="7" place="7" resultid="11864" />
                    <RANKING order="8" place="8" resultid="11339" />
                    <RANKING order="9" place="9" resultid="9997" />
                    <RANKING order="10" place="10" resultid="9162" />
                    <RANKING order="11" place="11" resultid="10049" />
                    <RANKING order="12" place="12" resultid="9269" />
                    <RANKING order="13" place="13" resultid="12872" />
                    <RANKING order="14" place="14" resultid="9439" />
                    <RANKING order="15" place="15" resultid="9321" />
                    <RANKING order="16" place="-1" resultid="9620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15156" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10474" />
                    <RANKING order="2" place="2" resultid="10579" />
                    <RANKING order="3" place="3" resultid="11331" />
                    <RANKING order="4" place="4" resultid="8915" />
                    <RANKING order="5" place="5" resultid="11125" />
                    <RANKING order="6" place="6" resultid="9051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15157" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13223" />
                    <RANKING order="2" place="2" resultid="11284" />
                    <RANKING order="3" place="3" resultid="11927" />
                    <RANKING order="4" place="4" resultid="11891" />
                    <RANKING order="5" place="-1" resultid="11785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15158" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11079" />
                    <RANKING order="2" place="2" resultid="9804" />
                    <RANKING order="3" place="3" resultid="9526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15159" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12817" />
                    <RANKING order="2" place="2" resultid="10543" />
                    <RANKING order="3" place="3" resultid="9886" />
                    <RANKING order="4" place="4" resultid="10635" />
                    <RANKING order="5" place="5" resultid="10878" />
                    <RANKING order="6" place="6" resultid="11755" />
                    <RANKING order="7" place="7" resultid="9405" />
                    <RANKING order="8" place="8" resultid="9412" />
                    <RANKING order="9" place="9" resultid="9691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15160" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11258" />
                    <RANKING order="2" place="2" resultid="11394" />
                    <RANKING order="3" place="3" resultid="8837" />
                    <RANKING order="4" place="4" resultid="10628" />
                    <RANKING order="5" place="5" resultid="10450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15161" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8863" />
                    <RANKING order="2" place="2" resultid="9539" />
                    <RANKING order="3" place="3" resultid="9832" />
                    <RANKING order="4" place="4" resultid="10622" />
                    <RANKING order="5" place="5" resultid="10442" />
                    <RANKING order="6" place="6" resultid="10501" />
                    <RANKING order="7" place="7" resultid="9733" />
                    <RANKING order="8" place="-1" resultid="9921" />
                    <RANKING order="9" place="-1" resultid="11736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15162" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10530" />
                    <RANKING order="2" place="2" resultid="11157" />
                    <RANKING order="3" place="3" resultid="10436" />
                    <RANKING order="4" place="4" resultid="8829" />
                    <RANKING order="5" place="5" resultid="11812" />
                    <RANKING order="6" place="6" resultid="8811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15163" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11381" />
                    <RANKING order="2" place="2" resultid="10431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15164" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15165" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14198" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14199" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14200" daytime="09:17" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14201" daytime="09:19" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14202" daytime="09:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14203" daytime="09:23" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14204" daytime="09:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14205" daytime="09:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14206" daytime="09:27" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14207" daytime="09:29" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8341" daytime="12:31" gender="M" number="19" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15271" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11133" />
                    <RANKING order="2" place="2" resultid="9628" />
                    <RANKING order="3" place="3" resultid="10331" />
                    <RANKING order="4" place="-1" resultid="10316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15272" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12767" />
                    <RANKING order="2" place="2" resultid="9649" />
                    <RANKING order="3" place="-1" resultid="9453" />
                    <RANKING order="4" place="-1" resultid="9943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15273" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12366" />
                    <RANKING order="2" place="2" resultid="12758" />
                    <RANKING order="3" place="3" resultid="9375" />
                    <RANKING order="4" place="-1" resultid="10239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15274" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9975" />
                    <RANKING order="2" place="2" resultid="9981" />
                    <RANKING order="3" place="3" resultid="10723" />
                    <RANKING order="4" place="4" resultid="12025" />
                    <RANKING order="5" place="-1" resultid="12004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15275" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9644" />
                    <RANKING order="2" place="2" resultid="8931" />
                    <RANKING order="3" place="3" resultid="9163" />
                    <RANKING order="4" place="4" resultid="10996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15276" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10574" />
                    <RANKING order="2" place="2" resultid="8945" />
                    <RANKING order="3" place="3" resultid="9056" />
                    <RANKING order="4" place="4" resultid="11018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15277" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8938" />
                    <RANKING order="2" place="2" resultid="11211" />
                    <RANKING order="3" place="3" resultid="12398" />
                    <RANKING order="4" place="4" resultid="8847" />
                    <RANKING order="5" place="5" resultid="8906" />
                    <RANKING order="6" place="-1" resultid="9467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15278" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9596" />
                    <RANKING order="2" place="2" resultid="11956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15279" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12818" />
                    <RANKING order="2" place="2" resultid="11204" />
                    <RANKING order="3" place="3" resultid="9664" />
                    <RANKING order="4" place="4" resultid="9854" />
                    <RANKING order="5" place="5" resultid="9840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15280" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11730" />
                    <RANKING order="2" place="2" resultid="8838" />
                    <RANKING order="3" place="3" resultid="10519" />
                    <RANKING order="4" place="4" resultid="10451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15281" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10253" />
                    <RANKING order="2" place="2" resultid="11822" />
                    <RANKING order="3" place="3" resultid="8874" />
                    <RANKING order="4" place="-1" resultid="9710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15282" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8855" />
                    <RANKING order="2" place="2" resultid="8830" />
                    <RANKING order="3" place="-1" resultid="8884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15283" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15284" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15285" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14258" daytime="12:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14259" daytime="12:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14260" daytime="12:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14261" daytime="12:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14262" daytime="12:52" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8261" daytime="10:29" gender="F" number="14" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15196" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9385" />
                    <RANKING order="2" place="2" resultid="10789" />
                    <RANKING order="3" place="-1" resultid="10809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15197" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9339" />
                    <RANKING order="2" place="2" resultid="10959" />
                    <RANKING order="3" place="3" resultid="9196" />
                    <RANKING order="4" place="4" resultid="10779" />
                    <RANKING order="5" place="-1" resultid="9489" />
                    <RANKING order="6" place="-1" resultid="12795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15198" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11724" />
                    <RANKING order="2" place="2" resultid="10261" />
                    <RANKING order="3" place="3" resultid="10748" />
                    <RANKING order="4" place="4" resultid="12441" />
                    <RANKING order="5" place="5" resultid="13298" />
                    <RANKING order="6" place="6" resultid="12406" />
                    <RANKING order="7" place="7" resultid="10267" />
                    <RANKING order="8" place="8" resultid="11050" />
                    <RANKING order="9" place="9" resultid="12097" />
                    <RANKING order="10" place="-1" resultid="9202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15199" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9461" />
                    <RANKING order="2" place="2" resultid="9060" />
                    <RANKING order="3" place="3" resultid="12827" />
                    <RANKING order="4" place="4" resultid="9811" />
                    <RANKING order="5" place="5" resultid="12434" />
                    <RANKING order="6" place="6" resultid="10690" />
                    <RANKING order="7" place="7" resultid="9074" />
                    <RANKING order="8" place="-1" resultid="12379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15200" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8799" />
                    <RANKING order="2" place="2" resultid="10059" />
                    <RANKING order="3" place="3" resultid="10981" />
                    <RANKING order="4" place="4" resultid="13209" />
                    <RANKING order="5" place="5" resultid="11837" />
                    <RANKING order="6" place="6" resultid="11850" />
                    <RANKING order="7" place="7" resultid="11800" />
                    <RANKING order="8" place="8" resultid="10734" />
                    <RANKING order="9" place="9" resultid="12032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15201" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9679" />
                    <RANKING order="2" place="2" resultid="9588" />
                    <RANKING order="3" place="3" resultid="11713" />
                    <RANKING order="4" place="4" resultid="13284" />
                    <RANKING order="5" place="5" resultid="12890" />
                    <RANKING order="6" place="-1" resultid="9684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15202" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12783" />
                    <RANKING order="2" place="2" resultid="10587" />
                    <RANKING order="3" place="3" resultid="11964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15203" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11701" />
                    <RANKING order="2" place="2" resultid="9700" />
                    <RANKING order="3" place="3" resultid="10862" />
                    <RANKING order="4" place="4" resultid="10507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15204" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9563" />
                    <RANKING order="2" place="2" resultid="11972" />
                    <RANKING order="3" place="3" resultid="9331" />
                    <RANKING order="4" place="4" resultid="10411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15205" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10649" />
                    <RANKING order="2" place="2" resultid="12012" />
                    <RANKING order="3" place="3" resultid="10886" />
                    <RANKING order="4" place="4" resultid="11299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15206" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15207" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15208" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15209" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15210" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14218" daytime="10:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14219" daytime="10:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14220" daytime="10:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14221" daytime="10:37" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14222" daytime="10:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14223" daytime="10:42" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8373" daytime="13:09" gender="M" number="21" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15600" agemax="99" agemin="80" name="80-99" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15601" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9222" />
                    <RANKING order="2" place="2" resultid="12920" />
                    <RANKING order="3" place="3" resultid="11184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15602" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10310" />
                    <RANKING order="2" place="2" resultid="9221" />
                    <RANKING order="3" place="3" resultid="10082" />
                    <RANKING order="4" place="4" resultid="11404" />
                    <RANKING order="5" place="5" resultid="10459" />
                    <RANKING order="6" place="6" resultid="10975" />
                    <RANKING order="7" place="7" resultid="11182" />
                    <RANKING order="8" place="8" resultid="10083" />
                    <RANKING order="9" place="9" resultid="9285" />
                    <RANKING order="10" place="10" resultid="10977" />
                    <RANKING order="11" place="11" resultid="10084" />
                    <RANKING order="12" place="12" resultid="9220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15603" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12038" />
                    <RANKING order="2" place="2" resultid="9932" />
                    <RANKING order="3" place="3" resultid="11151" />
                    <RANKING order="4" place="4" resultid="11031" />
                    <RANKING order="5" place="5" resultid="11903" />
                    <RANKING order="6" place="6" resultid="12455" />
                    <RANKING order="7" place="7" resultid="9449" />
                    <RANKING order="8" place="-1" resultid="10837" />
                    <RANKING order="9" place="-1" resultid="12039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15604" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11405" />
                    <RANKING order="2" place="2" resultid="12924" />
                    <RANKING order="3" place="3" resultid="10460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15605" agemax="279" agemin="240" name="240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9934" />
                    <RANKING order="2" place="2" resultid="11795" />
                    <RANKING order="3" place="3" resultid="9780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15606" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9556" />
                    <RANKING order="2" place="2" resultid="10539" />
                    <RANKING order="3" place="3" resultid="12726" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14265" daytime="13:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14266" daytime="13:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14267" daytime="13:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14268" daytime="13:21" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8293" daytime="11:24" gender="F" number="16" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15226" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11919" />
                    <RANKING order="2" place="2" resultid="9110" />
                    <RANKING order="3" place="3" resultid="12083" />
                    <RANKING order="4" place="4" resultid="8981" />
                    <RANKING order="5" place="5" resultid="10614" />
                    <RANKING order="6" place="6" resultid="10740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15227" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9340" />
                    <RANKING order="2" place="2" resultid="10960" />
                    <RANKING order="3" place="3" resultid="10742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15228" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9210" />
                    <RANKING order="2" place="2" resultid="10402" />
                    <RANKING order="3" place="3" resultid="11831" />
                    <RANKING order="4" place="4" resultid="8953" />
                    <RANKING order="5" place="5" resultid="11311" />
                    <RANKING order="6" place="6" resultid="10767" />
                    <RANKING order="7" place="7" resultid="10395" />
                    <RANKING order="8" place="8" resultid="12098" />
                    <RANKING order="9" place="-1" resultid="9203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15229" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11244" />
                    <RANKING order="2" place="2" resultid="9064" />
                    <RANKING order="3" place="3" resultid="9075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15230" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9579" />
                    <RANKING order="2" place="2" resultid="8800" />
                    <RANKING order="3" place="3" resultid="9861" />
                    <RANKING order="4" place="4" resultid="9263" />
                    <RANKING order="5" place="5" resultid="11035" />
                    <RANKING order="6" place="6" resultid="10982" />
                    <RANKING order="7" place="7" resultid="11005" />
                    <RANKING order="8" place="8" resultid="12801" />
                    <RANKING order="9" place="9" resultid="12467" />
                    <RANKING order="10" place="10" resultid="9769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15231" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9913" />
                    <RANKING order="2" place="2" resultid="12372" />
                    <RANKING order="3" place="3" resultid="13285" />
                    <RANKING order="4" place="4" resultid="11229" />
                    <RANKING order="5" place="5" resultid="13289" />
                    <RANKING order="6" place="6" resultid="11844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15232" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9673" />
                    <RANKING order="2" place="2" resultid="10680" />
                    <RANKING order="3" place="3" resultid="9605" />
                    <RANKING order="4" place="4" resultid="11706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15233" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9868" />
                    <RANKING order="2" place="2" resultid="12047" />
                    <RANKING order="3" place="3" resultid="11856" />
                    <RANKING order="4" place="4" resultid="13293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15234" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11997" />
                    <RANKING order="2" place="2" resultid="11411" />
                    <RANKING order="3" place="3" resultid="12459" />
                    <RANKING order="4" place="-1" resultid="11695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15235" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10524" />
                    <RANKING order="2" place="2" resultid="8768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15236" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13220" />
                    <RANKING order="2" place="2" resultid="9719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15237" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15238" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15239" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15240" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14238" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14239" daytime="11:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14240" daytime="11:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14241" daytime="11:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14242" daytime="11:37" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14243" daytime="11:39" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8309" daytime="11:44" gender="M" number="17" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15241" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10324" />
                    <RANKING order="2" place="2" resultid="8987" />
                    <RANKING order="3" place="3" resultid="10595" />
                    <RANKING order="4" place="4" resultid="8924" />
                    <RANKING order="5" place="5" resultid="10608" />
                    <RANKING order="6" place="6" resultid="10601" />
                    <RANKING order="7" place="-1" resultid="10774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15242" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9028" />
                    <RANKING order="2" place="2" resultid="9152" />
                    <RANKING order="3" place="3" resultid="12766" />
                    <RANKING order="4" place="4" resultid="9146" />
                    <RANKING order="5" place="5" resultid="11323" />
                    <RANKING order="6" place="-1" resultid="11399" />
                    <RANKING order="7" place="-1" resultid="10799" />
                    <RANKING order="8" place="-1" resultid="10804" />
                    <RANKING order="9" place="-1" resultid="10949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15243" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9827" />
                    <RANKING order="2" place="2" resultid="9419" />
                    <RANKING order="3" place="3" resultid="10289" />
                    <RANKING order="4" place="4" resultid="10965" />
                    <RANKING order="5" place="5" resultid="10297" />
                    <RANKING order="6" place="6" resultid="9135" />
                    <RANKING order="7" place="7" resultid="10673" />
                    <RANKING order="8" place="8" resultid="10729" />
                    <RANKING order="9" place="9" resultid="9374" />
                    <RANKING order="10" place="10" resultid="10933" />
                    <RANKING order="11" place="11" resultid="9274" />
                    <RANKING order="12" place="12" resultid="12091" />
                    <RANKING order="13" place="-1" resultid="9482" />
                    <RANKING order="14" place="-1" resultid="9927" />
                    <RANKING order="15" place="-1" resultid="10551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15244" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11305" />
                    <RANKING order="2" place="2" resultid="10042" />
                    <RANKING order="3" place="3" resultid="9905" />
                    <RANKING order="4" place="4" resultid="10368" />
                    <RANKING order="5" place="5" resultid="12077" />
                    <RANKING order="6" place="6" resultid="9753" />
                    <RANKING order="7" place="7" resultid="10387" />
                    <RANKING order="8" place="8" resultid="10064" />
                    <RANKING order="9" place="9" resultid="10361" />
                    <RANKING order="10" place="10" resultid="10012" />
                    <RANKING order="11" place="11" resultid="10939" />
                    <RANKING order="12" place="12" resultid="10018" />
                    <RANKING order="13" place="13" resultid="10971" />
                    <RANKING order="14" place="14" resultid="10037" />
                    <RANKING order="15" place="-1" resultid="10305" />
                    <RANKING order="16" place="-1" resultid="9875" />
                    <RANKING order="17" place="-1" resultid="10077" />
                    <RANKING order="18" place="-1" resultid="11238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15245" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12836" />
                    <RANKING order="2" place="2" resultid="9990" />
                    <RANKING order="3" place="3" resultid="10244" />
                    <RANKING order="4" place="4" resultid="9281" />
                    <RANKING order="5" place="5" resultid="9798" />
                    <RANKING order="6" place="6" resultid="9621" />
                    <RANKING order="7" place="7" resultid="11865" />
                    <RANKING order="8" place="8" resultid="9446" />
                    <RANKING order="9" place="9" resultid="9257" />
                    <RANKING order="10" place="10" resultid="12104" />
                    <RANKING order="11" place="11" resultid="8787" />
                    <RANKING order="12" place="12" resultid="10926" />
                    <RANKING order="13" place="13" resultid="9441" />
                    <RANKING order="14" place="14" resultid="10920" />
                    <RANKING order="15" place="15" resultid="9322" />
                    <RANKING order="16" place="-1" resultid="10662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15246" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10580" />
                    <RANKING order="2" place="2" resultid="9636" />
                    <RANKING order="3" place="3" resultid="10475" />
                    <RANKING order="4" place="4" resultid="11332" />
                    <RANKING order="5" place="5" resultid="10826" />
                    <RANKING order="6" place="6" resultid="10834" />
                    <RANKING order="7" place="7" resultid="11886" />
                    <RANKING order="8" place="8" resultid="12879" />
                    <RANKING order="9" place="9" resultid="11367" />
                    <RANKING order="10" place="10" resultid="9435" />
                    <RANKING order="11" place="-1" resultid="11106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15247" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13224" />
                    <RANKING order="2" place="2" resultid="11285" />
                    <RANKING order="3" place="3" resultid="12426" />
                    <RANKING order="4" place="4" resultid="11786" />
                    <RANKING order="5" place="5" resultid="9950" />
                    <RANKING order="6" place="6" resultid="11776" />
                    <RANKING order="7" place="7" resultid="9429" />
                    <RANKING order="8" place="-1" resultid="11272" />
                    <RANKING order="9" place="-1" resultid="9847" />
                    <RANKING order="10" place="-1" resultid="11911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15248" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9037" />
                    <RANKING order="2" place="2" resultid="11080" />
                    <RANKING order="3" place="3" resultid="12865" />
                    <RANKING order="4" place="4" resultid="9089" />
                    <RANKING order="5" place="5" resultid="9739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15249" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9887" />
                    <RANKING order="2" place="2" resultid="9126" />
                    <RANKING order="3" place="3" resultid="10636" />
                    <RANKING order="4" place="4" resultid="10348" />
                    <RANKING order="5" place="5" resultid="11266" />
                    <RANKING order="6" place="6" resultid="9413" />
                    <RANKING order="7" place="7" resultid="9853" />
                    <RANKING order="8" place="-1" resultid="12390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15250" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11749" />
                    <RANKING order="2" place="2" resultid="11395" />
                    <RANKING order="3" place="3" resultid="11375" />
                    <RANKING order="4" place="4" resultid="11729" />
                    <RANKING order="5" place="5" resultid="9532" />
                    <RANKING order="6" place="6" resultid="9352" />
                    <RANKING order="7" place="-1" resultid="10514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15251" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10623" />
                    <RANKING order="2" place="2" resultid="9536" />
                    <RANKING order="3" place="3" resultid="10502" />
                    <RANKING order="4" place="4" resultid="8821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15252" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15253" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15254" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15255" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14244" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14245" daytime="11:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14246" daytime="11:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14247" daytime="11:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14248" daytime="11:58" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14249" daytime="12:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14250" daytime="12:02" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14251" daytime="12:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14252" daytime="12:07" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14253" daytime="12:09" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14254" daytime="12:11" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14255" daytime="12:13" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8229" daytime="09:33" gender="F" number="12" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15166" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11918" />
                    <RANKING order="2" place="2" resultid="12749" />
                    <RANKING order="3" place="3" resultid="10613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15167" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11350" />
                    <RANKING order="2" place="2" resultid="9190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15168" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10401" />
                    <RANKING order="2" place="2" resultid="10274" />
                    <RANKING order="3" place="3" resultid="8952" />
                    <RANKING order="4" place="4" resultid="12069" />
                    <RANKING order="5" place="5" resultid="11830" />
                    <RANKING order="6" place="6" resultid="10394" />
                    <RANKING order="7" place="-1" resultid="9201" />
                    <RANKING order="8" place="-1" resultid="10266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15169" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15170" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9578" />
                    <RANKING order="2" place="2" resultid="8958" />
                    <RANKING order="3" place="3" resultid="11004" />
                    <RANKING order="4" place="4" resultid="11346" />
                    <RANKING order="5" place="5" resultid="9970" />
                    <RANKING order="6" place="6" resultid="10028" />
                    <RANKING order="7" place="7" resultid="11991" />
                    <RANKING order="8" place="8" resultid="12031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15171" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9544" />
                    <RANKING order="2" place="2" resultid="11228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15172" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9604" />
                    <RANKING order="2" place="2" resultid="12782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15173" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9045" />
                    <RANKING order="2" place="2" resultid="13292" />
                    <RANKING order="3" place="3" resultid="11983" />
                    <RANKING order="4" place="4" resultid="9726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15174" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11996" />
                    <RANKING order="2" place="2" resultid="10870" />
                    <RANKING order="3" place="3" resultid="11971" />
                    <RANKING order="4" place="4" resultid="11063" />
                    <RANKING order="5" place="-1" resultid="11694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15175" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12011" />
                    <RANKING order="2" place="2" resultid="9514" />
                    <RANKING order="3" place="3" resultid="8767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15176" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15177" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15178" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15179" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15180" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14208" daytime="09:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14209" daytime="09:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14210" daytime="09:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14211" daytime="09:51" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8196" daytime="09:00" gender="F" number="10" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15136" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10335" />
                    <RANKING order="2" place="2" resultid="9892" />
                    <RANKING order="3" place="3" resultid="8996" />
                    <RANKING order="4" place="4" resultid="9384" />
                    <RANKING order="5" place="5" resultid="12748" />
                    <RANKING order="6" place="6" resultid="10785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15137" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9195" />
                    <RANKING order="2" place="2" resultid="10668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15138" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9209" />
                    <RANKING order="2" place="2" resultid="11723" />
                    <RANKING order="3" place="3" resultid="12440" />
                    <RANKING order="4" place="4" resultid="12896" />
                    <RANKING order="5" place="-1" resultid="10684" />
                    <RANKING order="6" place="-1" resultid="12111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15139" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9062" />
                    <RANKING order="2" place="2" resultid="12826" />
                    <RANKING order="3" place="3" resultid="10034" />
                    <RANKING order="4" place="4" resultid="12813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15140" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9262" />
                    <RANKING order="2" place="2" resultid="9860" />
                    <RANKING order="3" place="3" resultid="12800" />
                    <RANKING order="4" place="4" resultid="11849" />
                    <RANKING order="5" place="5" resultid="12466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15141" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9912" />
                    <RANKING order="2" place="2" resultid="11712" />
                    <RANKING order="3" place="3" resultid="9587" />
                    <RANKING order="4" place="4" resultid="10419" />
                    <RANKING order="5" place="5" resultid="12889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15142" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9672" />
                    <RANKING order="2" place="2" resultid="10679" />
                    <RANKING order="3" place="3" resultid="11963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15143" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9867" />
                    <RANKING order="2" place="2" resultid="12046" />
                    <RANKING order="3" place="3" resultid="11700" />
                    <RANKING order="4" place="4" resultid="10506" />
                    <RANKING order="5" place="5" resultid="10861" />
                    <RANKING order="6" place="-1" resultid="11855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15144" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9562" />
                    <RANKING order="2" place="2" resultid="9761" />
                    <RANKING order="3" place="3" resultid="9330" />
                    <RANKING order="4" place="4" resultid="10410" />
                    <RANKING order="5" place="5" resultid="12458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15145" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9500" />
                    <RANKING order="2" place="2" resultid="10648" />
                    <RANKING order="3" place="3" resultid="10885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15146" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11361" />
                    <RANKING order="2" place="2" resultid="9551" />
                    <RANKING order="3" place="3" resultid="8803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15147" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15148" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15149" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15150" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14193" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14194" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14195" daytime="09:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14196" daytime="09:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14197" daytime="09:08" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8325" daytime="12:18" gender="F" number="18" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15256" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15257" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15258" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12897" />
                    <RANKING order="2" place="2" resultid="10275" />
                    <RANKING order="3" place="3" resultid="12407" />
                    <RANKING order="4" place="4" resultid="11312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15259" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10073" />
                    <RANKING order="2" place="2" resultid="11130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15260" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10467" />
                    <RANKING order="2" place="2" resultid="10703" />
                    <RANKING order="3" place="3" resultid="11145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15261" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15262" agemax="54" agemin="50" name="50-54" />
                <AGEGROUP agegroupid="15263" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9701" />
                    <RANKING order="2" place="2" resultid="9048" />
                    <RANKING order="3" place="3" resultid="11984" />
                    <RANKING order="4" place="4" resultid="9727" />
                    <RANKING order="5" place="-1" resultid="11056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15264" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9762" />
                    <RANKING order="2" place="2" resultid="10871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15265" agemax="69" agemin="65" name="65-69" />
                <AGEGROUP agegroupid="15266" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15267" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15268" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15269" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15270" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14256" daytime="12:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14257" daytime="12:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8357" daytime="12:59" gender="F" number="20" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15593" agemax="99" agemin="80" name="80-99" calculate="TOTAL" />
                <AGEGROUP agegroupid="15594" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12922" />
                    <RANKING order="2" place="-1" resultid="11178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15595" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9224" />
                    <RANKING order="2" place="2" resultid="11180" />
                    <RANKING order="3" place="-1" resultid="10081" />
                    <RANKING order="4" place="-1" resultid="10693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15596" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9930" />
                    <RANKING order="2" place="2" resultid="10458" />
                    <RANKING order="3" place="-1" resultid="11902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15597" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9778" />
                    <RANKING order="2" place="2" resultid="12037" />
                    <RANKING order="3" place="-1" resultid="11793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15598" agemax="279" agemin="240" name="240-279" calculate="TOTAL" />
                <AGEGROUP agegroupid="15599" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9555" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14263" daytime="12:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14264" daytime="13:03" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-11-17" daytime="16:00" endtime="21:27" name="III Blok" number="3" warmupfrom="15:00" warmupuntil="15:00">
          <EVENTS>
            <EVENT eventid="8518" daytime="18:41" gender="M" number="29" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15391" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10333" />
                    <RANKING order="2" place="2" resultid="9658" />
                    <RANKING order="3" place="3" resultid="9629" />
                    <RANKING order="4" place="4" resultid="9363" />
                    <RANKING order="5" place="-1" resultid="9023" />
                    <RANKING order="6" place="-1" resultid="10603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15392" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9476" />
                    <RANKING order="2" place="2" resultid="11401" />
                    <RANKING order="3" place="3" resultid="9107" />
                    <RANKING order="4" place="4" resultid="12853" />
                    <RANKING order="5" place="5" resultid="12021" />
                    <RANKING order="6" place="-1" resultid="11142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15393" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9928" />
                    <RANKING order="2" place="2" resultid="11328" />
                    <RANKING order="3" place="3" resultid="9174" />
                    <RANKING order="4" place="4" resultid="9316" />
                    <RANKING order="5" place="5" resultid="10299" />
                    <RANKING order="6" place="6" resultid="9376" />
                    <RANKING order="7" place="7" resultid="9484" />
                    <RANKING order="8" place="8" resultid="10719" />
                    <RANKING order="9" place="9" resultid="10375" />
                    <RANKING order="10" place="10" resultid="12093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15394" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11253" />
                    <RANKING order="2" place="2" resultid="12026" />
                    <RANKING order="3" place="3" resultid="10560" />
                    <RANKING order="4" place="4" resultid="11880" />
                    <RANKING order="5" place="5" resultid="12809" />
                    <RANKING order="6" place="6" resultid="10427" />
                    <RANKING order="7" place="7" resultid="10972" />
                    <RANKING order="8" place="8" resultid="9967" />
                    <RANKING order="9" place="9" resultid="9426" />
                    <RANKING order="10" place="10" resultid="9017" />
                    <RANKING order="11" place="-1" resultid="8869" />
                    <RANKING order="12" place="-1" resultid="10014" />
                    <RANKING order="13" place="-1" resultid="10955" />
                    <RANKING order="14" place="-1" resultid="11240" />
                    <RANKING order="15" place="-1" resultid="12005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15395" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12837" />
                    <RANKING order="2" place="2" resultid="10991" />
                    <RANKING order="3" place="3" resultid="8932" />
                    <RANKING order="4" place="4" resultid="12905" />
                    <RANKING order="5" place="5" resultid="9992" />
                    <RANKING order="6" place="6" resultid="11342" />
                    <RANKING order="7" place="7" resultid="9800" />
                    <RANKING order="8" place="8" resultid="9448" />
                    <RANKING order="9" place="9" resultid="11873" />
                    <RANKING order="10" place="10" resultid="10997" />
                    <RANKING order="11" place="11" resultid="10051" />
                    <RANKING order="12" place="12" resultid="12450" />
                    <RANKING order="13" place="13" resultid="9258" />
                    <RANKING order="14" place="14" resultid="12875" />
                    <RANKING order="15" place="15" resultid="9008" />
                    <RANKING order="16" place="16" resultid="8789" />
                    <RANKING order="17" place="17" resultid="11150" />
                    <RANKING order="18" place="18" resultid="10928" />
                    <RANKING order="19" place="-1" resultid="11318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15396" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10582" />
                    <RANKING order="2" place="2" resultid="11390" />
                    <RANKING order="3" place="3" resultid="9637" />
                    <RANKING order="4" place="4" resultid="10699" />
                    <RANKING order="5" place="5" resultid="10836" />
                    <RANKING order="6" place="6" resultid="11334" />
                    <RANKING order="7" place="7" resultid="8900" />
                    <RANKING order="8" place="8" resultid="9348" />
                    <RANKING order="9" place="9" resultid="9437" />
                    <RANKING order="10" place="10" resultid="11369" />
                    <RANKING order="11" place="-1" resultid="10827" />
                    <RANKING order="12" place="-1" resultid="11108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15397" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8939" />
                    <RANKING order="2" place="2" resultid="12427" />
                    <RANKING order="3" place="3" resultid="11807" />
                    <RANKING order="4" place="4" resultid="11929" />
                    <RANKING order="5" place="5" resultid="11213" />
                    <RANKING order="6" place="6" resultid="11778" />
                    <RANKING order="7" place="7" resultid="12912" />
                    <RANKING order="8" place="8" resultid="9396" />
                    <RANKING order="9" place="9" resultid="9431" />
                    <RANKING order="10" place="10" resultid="11274" />
                    <RANKING order="11" place="-1" resultid="9849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15398" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9962" />
                    <RANKING order="2" place="2" resultid="9082" />
                    <RANKING order="3" place="3" resultid="9807" />
                    <RANKING order="4" place="4" resultid="9597" />
                    <RANKING order="5" place="5" resultid="11958" />
                    <RANKING order="6" place="6" resultid="9401" />
                    <RANKING order="7" place="7" resultid="11295" />
                    <RANKING order="8" place="-1" resultid="11762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15399" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12820" />
                    <RANKING order="2" place="2" resultid="8780" />
                    <RANKING order="3" place="3" resultid="12392" />
                    <RANKING order="4" place="4" resultid="12054" />
                    <RANKING order="5" place="5" resultid="10881" />
                    <RANKING order="6" place="6" resultid="9841" />
                    <RANKING order="7" place="7" resultid="9694" />
                    <RANKING order="8" place="-1" resultid="9004" />
                    <RANKING order="9" place="-1" resultid="10546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15400" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11261" />
                    <RANKING order="2" place="2" resultid="10356" />
                    <RANKING order="3" place="3" resultid="11732" />
                    <RANKING order="4" place="4" resultid="9354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15401" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9711" />
                    <RANKING order="2" place="2" resultid="11823" />
                    <RANKING order="3" place="3" resultid="8795" />
                    <RANKING order="4" place="4" resultid="12791" />
                    <RANKING order="5" place="5" resultid="8876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15402" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10892" />
                    <RANKING order="2" place="2" resultid="9748" />
                    <RANKING order="3" place="3" resultid="8814" />
                    <RANKING order="4" place="-1" resultid="8885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15403" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15404" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9310" />
                    <RANKING order="2" place="2" resultid="9100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15405" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14322" daytime="18:41" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14323" daytime="18:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14324" daytime="18:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14325" daytime="18:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14326" daytime="19:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14327" daytime="19:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14328" daytime="19:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14329" daytime="19:13" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14330" daytime="19:17" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14331" daytime="19:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14332" daytime="19:23" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14333" daytime="19:27" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8486" daytime="17:46" gender="M" number="27" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15361" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10795" />
                    <RANKING order="2" place="2" resultid="10597" />
                    <RANKING order="3" place="3" resultid="10318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15362" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9495" />
                    <RANKING order="2" place="2" resultid="12768" />
                    <RANKING order="3" place="3" resultid="11324" />
                    <RANKING order="4" place="4" resultid="12744" />
                    <RANKING order="5" place="-1" resultid="9944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15363" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10291" />
                    <RANKING order="2" place="2" resultid="12361" />
                    <RANKING order="3" place="3" resultid="10675" />
                    <RANKING order="4" place="4" resultid="9276" />
                    <RANKING order="5" place="-1" resultid="10553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15364" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10307" />
                    <RANKING order="2" place="2" resultid="9983" />
                    <RANKING order="3" place="3" resultid="9877" />
                    <RANKING order="4" place="4" resultid="10369" />
                    <RANKING order="5" place="5" resultid="10388" />
                    <RANKING order="6" place="6" resultid="9754" />
                    <RANKING order="7" place="7" resultid="10559" />
                    <RANKING order="8" place="8" resultid="10019" />
                    <RANKING order="9" place="-1" resultid="11307" />
                    <RANKING order="10" place="-1" resultid="12420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15365" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9158" />
                    <RANKING order="2" place="2" resultid="9614" />
                    <RANKING order="3" place="3" resultid="11937" />
                    <RANKING order="4" place="4" resultid="9283" />
                    <RANKING order="5" place="5" resultid="9622" />
                    <RANKING order="6" place="6" resultid="11899" />
                    <RANKING order="7" place="7" resultid="11866" />
                    <RANKING order="8" place="8" resultid="9270" />
                    <RANKING order="9" place="9" resultid="9324" />
                    <RANKING order="10" place="-1" resultid="9164" />
                    <RANKING order="11" place="-1" resultid="9442" />
                    <RANKING order="12" place="-1" resultid="10000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15366" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10477" />
                    <RANKING order="2" place="2" resultid="8918" />
                    <RANKING order="3" place="3" resultid="9052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15367" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13225" />
                    <RANKING order="2" place="2" resultid="11287" />
                    <RANKING order="3" place="3" resultid="11928" />
                    <RANKING order="4" place="4" resultid="11787" />
                    <RANKING order="5" place="5" resultid="11212" />
                    <RANKING order="6" place="6" resultid="11893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15368" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9039" />
                    <RANKING order="2" place="2" resultid="11081" />
                    <RANKING order="3" place="3" resultid="9528" />
                    <RANKING order="4" place="4" resultid="9091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15369" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9888" />
                    <RANKING order="2" place="2" resultid="9128" />
                    <RANKING order="3" place="3" resultid="10637" />
                    <RANKING order="4" place="4" resultid="10880" />
                    <RANKING order="5" place="5" resultid="9406" />
                    <RANKING order="6" place="6" resultid="9855" />
                    <RANKING order="7" place="-1" resultid="9003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15370" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11260" />
                    <RANKING order="2" place="2" resultid="11396" />
                    <RANKING order="3" place="3" resultid="8840" />
                    <RANKING order="4" place="4" resultid="9353" />
                    <RANKING order="5" place="5" resultid="10452" />
                    <RANKING order="6" place="-1" resultid="10629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15371" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9835" />
                    <RANKING order="2" place="2" resultid="9540" />
                    <RANKING order="3" place="3" resultid="10624" />
                    <RANKING order="4" place="4" resultid="9734" />
                    <RANKING order="5" place="-1" resultid="10445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15372" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11160" />
                    <RANKING order="2" place="2" resultid="10533" />
                    <RANKING order="3" place="3" resultid="10438" />
                    <RANKING order="4" place="4" resultid="11815" />
                    <RANKING order="5" place="5" resultid="8813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15373" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15374" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15375" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14308" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14309" daytime="17:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14310" daytime="17:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14311" daytime="17:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14312" daytime="18:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14313" daytime="18:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14314" daytime="18:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14315" daytime="18:06" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8404" daytime="16:00" gender="F" number="22" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15286" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11920" />
                    <RANKING order="2" place="2" resultid="9111" />
                    <RANKING order="3" place="3" resultid="9300" />
                    <RANKING order="4" place="4" resultid="8982" />
                    <RANKING order="5" place="5" resultid="12750" />
                    <RANKING order="6" place="6" resultid="10615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15287" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9010" />
                    <RANKING order="2" place="2" resultid="10743" />
                    <RANKING order="3" place="3" resultid="9490" />
                    <RANKING order="4" place="4" resultid="11351" />
                    <RANKING order="5" place="5" resultid="10669" />
                    <RANKING order="6" place="-1" resultid="9191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15288" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10262" />
                    <RANKING order="2" place="2" resultid="10403" />
                    <RANKING order="3" place="3" resultid="10276" />
                    <RANKING order="4" place="4" resultid="12070" />
                    <RANKING order="5" place="5" resultid="11832" />
                    <RANKING order="6" place="6" resultid="10768" />
                    <RANKING order="7" place="-1" resultid="9204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15289" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11245" />
                    <RANKING order="2" place="-1" resultid="12380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15290" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9580" />
                    <RANKING order="2" place="2" resultid="9862" />
                    <RANKING order="3" place="3" resultid="8959" />
                    <RANKING order="4" place="4" resultid="11347" />
                    <RANKING order="5" place="5" resultid="11006" />
                    <RANKING order="6" place="6" resultid="13210" />
                    <RANKING order="7" place="7" resultid="11992" />
                    <RANKING order="8" place="8" resultid="12033" />
                    <RANKING order="9" place="-1" resultid="11838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15291" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9545" />
                    <RANKING order="2" place="2" resultid="9589" />
                    <RANKING order="3" place="3" resultid="11230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15292" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10655" />
                    <RANKING order="2" place="2" resultid="9606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15293" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9044" />
                    <RANKING order="2" place="2" resultid="13294" />
                    <RANKING order="3" place="3" resultid="11985" />
                    <RANKING order="4" place="4" resultid="10863" />
                    <RANKING order="5" place="5" resultid="9728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15294" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11998" />
                    <RANKING order="2" place="2" resultid="11412" />
                    <RANKING order="3" place="3" resultid="10872" />
                    <RANKING order="4" place="4" resultid="12460" />
                    <RANKING order="5" place="5" resultid="11064" />
                    <RANKING order="6" place="-1" resultid="11696" />
                    <RANKING order="7" place="-1" resultid="11973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15295" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12013" />
                    <RANKING order="2" place="2" resultid="9515" />
                    <RANKING order="3" place="3" resultid="8769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15296" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9720" />
                    <RANKING order="2" place="2" resultid="8805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15297" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15298" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15299" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15300" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14269" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14270" daytime="16:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14271" daytime="16:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14272" daytime="16:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14273" daytime="16:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14274" daytime="16:16" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8454" daytime="17:03" gender="M" number="25" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15331" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10325" />
                    <RANKING order="2" place="2" resultid="10944" />
                    <RANKING order="3" place="3" resultid="10775" />
                    <RANKING order="4" place="4" resultid="10596" />
                    <RANKING order="5" place="5" resultid="8976" />
                    <RANKING order="6" place="6" resultid="10317" />
                    <RANKING order="7" place="7" resultid="11134" />
                    <RANKING order="8" place="8" resultid="8926" />
                    <RANKING order="9" place="9" resultid="12885" />
                    <RANKING order="10" place="10" resultid="10765" />
                    <RANKING order="11" place="11" resultid="10344" />
                    <RANKING order="12" place="12" resultid="10610" />
                    <RANKING order="13" place="13" resultid="10602" />
                    <RANKING order="14" place="14" resultid="8969" />
                    <RANKING order="15" place="15" resultid="10753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15332" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10950" />
                    <RANKING order="2" place="2" resultid="9030" />
                    <RANKING order="3" place="3" resultid="12852" />
                    <RANKING order="4" place="4" resultid="9650" />
                    <RANKING order="5" place="5" resultid="11400" />
                    <RANKING order="6" place="6" resultid="9148" />
                    <RANKING order="7" place="7" resultid="12020" />
                    <RANKING order="8" place="8" resultid="10757" />
                    <RANKING order="9" place="9" resultid="10761" />
                    <RANKING order="10" place="-1" resultid="12917" />
                    <RANKING order="11" place="-1" resultid="9455" />
                    <RANKING order="12" place="-1" resultid="11193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15333" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9828" />
                    <RANKING order="2" place="2" resultid="9421" />
                    <RANKING order="3" place="3" resultid="9143" />
                    <RANKING order="4" place="4" resultid="9136" />
                    <RANKING order="5" place="5" resultid="9918" />
                    <RANKING order="6" place="6" resultid="10966" />
                    <RANKING order="7" place="7" resultid="9483" />
                    <RANKING order="8" place="8" resultid="10298" />
                    <RANKING order="9" place="9" resultid="9173" />
                    <RANKING order="10" place="10" resultid="10071" />
                    <RANKING order="11" place="11" resultid="10934" />
                    <RANKING order="12" place="12" resultid="10374" />
                    <RANKING order="13" place="13" resultid="11356" />
                    <RANKING order="14" place="14" resultid="12092" />
                    <RANKING order="15" place="-1" resultid="9957" />
                    <RANKING order="16" place="-1" resultid="10290" />
                    <RANKING order="17" place="-1" resultid="10552" />
                    <RANKING order="18" place="-1" resultid="12367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15334" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10306" />
                    <RANKING order="2" place="2" resultid="10536" />
                    <RANKING order="3" place="3" resultid="11946" />
                    <RANKING order="4" place="4" resultid="9876" />
                    <RANKING order="5" place="5" resultid="10044" />
                    <RANKING order="6" place="6" resultid="12078" />
                    <RANKING order="7" place="7" resultid="9976" />
                    <RANKING order="8" place="8" resultid="11119" />
                    <RANKING order="9" place="9" resultid="9140" />
                    <RANKING order="10" place="10" resultid="10066" />
                    <RANKING order="11" place="11" resultid="10362" />
                    <RANKING order="12" place="12" resultid="10013" />
                    <RANKING order="13" place="13" resultid="10426" />
                    <RANKING order="14" place="14" resultid="10940" />
                    <RANKING order="15" place="-1" resultid="11138" />
                    <RANKING order="16" place="-1" resultid="9907" />
                    <RANKING order="17" place="-1" resultid="10954" />
                    <RANKING order="18" place="-1" resultid="11239" />
                    <RANKING order="19" place="-1" resultid="11306" />
                    <RANKING order="20" place="-1" resultid="12808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15335" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9157" />
                    <RANKING order="2" place="2" resultid="10246" />
                    <RANKING order="3" place="3" resultid="10990" />
                    <RANKING order="4" place="4" resultid="9991" />
                    <RANKING order="5" place="5" resultid="9799" />
                    <RANKING order="6" place="6" resultid="11952" />
                    <RANKING order="7" place="7" resultid="11341" />
                    <RANKING order="8" place="8" resultid="9447" />
                    <RANKING order="9" place="9" resultid="12846" />
                    <RANKING order="10" place="10" resultid="12106" />
                    <RANKING order="11" place="11" resultid="9999" />
                    <RANKING order="12" place="12" resultid="11115" />
                    <RANKING order="13" place="13" resultid="10921" />
                    <RANKING order="14" place="14" resultid="8788" />
                    <RANKING order="15" place="15" resultid="12874" />
                    <RANKING order="16" place="16" resultid="10927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15336" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10575" />
                    <RANKING order="2" place="2" resultid="10476" />
                    <RANKING order="3" place="3" resultid="11389" />
                    <RANKING order="4" place="4" resultid="11333" />
                    <RANKING order="5" place="5" resultid="10835" />
                    <RANKING order="6" place="6" resultid="11019" />
                    <RANKING order="7" place="7" resultid="9347" />
                    <RANKING order="8" place="8" resultid="8899" />
                    <RANKING order="9" place="9" resultid="11887" />
                    <RANKING order="10" place="-1" resultid="11107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15337" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11286" />
                    <RANKING order="2" place="2" resultid="9952" />
                    <RANKING order="3" place="3" resultid="8848" />
                    <RANKING order="4" place="-1" resultid="9848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15338" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9038" />
                    <RANKING order="2" place="2" resultid="9806" />
                    <RANKING order="3" place="3" resultid="11957" />
                    <RANKING order="4" place="4" resultid="9090" />
                    <RANKING order="5" place="5" resultid="11294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15339" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10545" />
                    <RANKING order="2" place="2" resultid="12819" />
                    <RANKING order="3" place="3" resultid="11205" />
                    <RANKING order="4" place="4" resultid="12391" />
                    <RANKING order="5" place="5" resultid="9414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15340" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10355" />
                    <RANKING order="2" place="2" resultid="9574" />
                    <RANKING order="3" place="3" resultid="11731" />
                    <RANKING order="4" place="4" resultid="9533" />
                    <RANKING order="5" place="5" resultid="8839" />
                    <RANKING order="6" place="-1" resultid="10516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15341" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9923" />
                    <RANKING order="2" place="2" resultid="10503" />
                    <RANKING order="3" place="3" resultid="8875" />
                    <RANKING order="4" place="4" resultid="9537" />
                    <RANKING order="5" place="5" resultid="10254" />
                    <RANKING order="6" place="6" resultid="8823" />
                    <RANKING order="7" place="-1" resultid="8864" />
                    <RANKING order="8" place="-1" resultid="11738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15342" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11159" />
                    <RANKING order="2" place="2" resultid="8857" />
                    <RANKING order="3" place="3" resultid="10891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15343" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15344" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15345" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14290" daytime="17:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14291" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14292" daytime="17:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14293" daytime="17:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14294" daytime="17:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14295" daytime="17:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14296" daytime="17:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14297" daytime="17:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14298" daytime="17:17" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14299" daytime="17:18" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14300" daytime="17:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14301" daytime="17:21" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14302" daytime="17:23" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8550" daytime="19:43" gender="M" number="31" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15614" agemax="99" agemin="80" name="80-99" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15615" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12926" />
                    <RANKING order="2" place="2" resultid="9217" />
                    <RANKING order="3" place="3" resultid="11185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15616" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9218" />
                    <RANKING order="2" place="2" resultid="10309" />
                    <RANKING order="3" place="3" resultid="11406" />
                    <RANKING order="4" place="4" resultid="12042" />
                    <RANKING order="5" place="5" resultid="10086" />
                    <RANKING order="6" place="6" resultid="10461" />
                    <RANKING order="7" place="7" resultid="10974" />
                    <RANKING order="8" place="8" resultid="11153" />
                    <RANKING order="9" place="9" resultid="11183" />
                    <RANKING order="10" place="10" resultid="9286" />
                    <RANKING order="11" place="11" resultid="10976" />
                    <RANKING order="12" place="12" resultid="10088" />
                    <RANKING order="13" place="-1" resultid="10087" />
                    <RANKING order="14" place="-1" resultid="9450" />
                    <RANKING order="15" place="-1" resultid="9219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15617" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12927" />
                    <RANKING order="2" place="2" resultid="11407" />
                    <RANKING order="3" place="3" resultid="11032" />
                    <RANKING order="4" place="4" resultid="11905" />
                    <RANKING order="5" place="5" resultid="9933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15618" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12928" />
                    <RANKING order="2" place="2" resultid="10462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15619" agemax="279" agemin="240" name="240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11796" />
                    <RANKING order="2" place="2" resultid="9935" />
                    <RANKING order="3" place="3" resultid="9779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15620" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9558" />
                    <RANKING order="2" place="2" resultid="10538" />
                    <RANKING order="3" place="-1" resultid="12727" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14336" daytime="19:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14337" daytime="19:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14338" daytime="19:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14339" daytime="19:53" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8438" daytime="16:51" gender="F" number="24" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15316" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12084" />
                    <RANKING order="2" place="2" resultid="10616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15317" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10961" />
                    <RANKING order="2" place="2" resultid="9011" />
                    <RANKING order="3" place="3" resultid="10744" />
                    <RANKING order="4" place="4" resultid="12775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15318" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11725" />
                    <RANKING order="2" place="2" resultid="12898" />
                    <RANKING order="3" place="3" resultid="11313" />
                    <RANKING order="4" place="4" resultid="13299" />
                    <RANKING order="5" place="5" resultid="12408" />
                    <RANKING order="6" place="6" resultid="10769" />
                    <RANKING order="7" place="7" resultid="10396" />
                    <RANKING order="8" place="-1" resultid="10685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15319" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11246" />
                    <RANKING order="2" place="2" resultid="9061" />
                    <RANKING order="3" place="3" resultid="12828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15320" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9581" />
                    <RANKING order="2" place="2" resultid="10060" />
                    <RANKING order="3" place="3" resultid="10468" />
                    <RANKING order="4" place="4" resultid="10983" />
                    <RANKING order="5" place="5" resultid="13211" />
                    <RANKING order="6" place="6" resultid="10029" />
                    <RANKING order="7" place="7" resultid="9770" />
                    <RANKING order="8" place="-1" resultid="11801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15321" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9899" />
                    <RANKING order="2" place="2" resultid="9680" />
                    <RANKING order="3" place="3" resultid="13286" />
                    <RANKING order="4" place="4" resultid="9685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15322" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9674" />
                    <RANKING order="2" place="2" resultid="10681" />
                    <RANKING order="3" place="3" resultid="11707" />
                    <RANKING order="4" place="4" resultid="9607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15323" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9869" />
                    <RANKING order="2" place="2" resultid="9702" />
                    <RANKING order="3" place="3" resultid="9046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15324" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11413" />
                    <RANKING order="2" place="2" resultid="9763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15325" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9501" />
                    <RANKING order="2" place="2" resultid="10650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15326" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15327" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9522" />
                    <RANKING order="2" place="2" resultid="9510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15328" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15329" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15330" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14285" daytime="16:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14286" daytime="16:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14287" daytime="16:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14288" daytime="16:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14289" daytime="16:59" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8470" daytime="17:27" gender="F" number="26" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15346" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10337" />
                    <RANKING order="2" place="2" resultid="8997" />
                    <RANKING order="3" place="3" resultid="9893" />
                    <RANKING order="4" place="4" resultid="12085" />
                    <RANKING order="5" place="5" resultid="9386" />
                    <RANKING order="6" place="6" resultid="12751" />
                    <RANKING order="7" place="7" resultid="10786" />
                    <RANKING order="8" place="-1" resultid="10790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15347" agemax="29" agemin="25" name="25-29" />
                <AGEGROUP agegroupid="15348" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9211" />
                    <RANKING order="2" place="2" resultid="12442" />
                    <RANKING order="3" place="3" resultid="10268" />
                    <RANKING order="4" place="-1" resultid="10686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15349" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12829" />
                    <RANKING order="2" place="2" resultid="9076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15350" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9863" />
                    <RANKING order="2" place="2" resultid="9264" />
                    <RANKING order="3" place="3" resultid="12802" />
                    <RANKING order="4" place="4" resultid="11851" />
                    <RANKING order="5" place="5" resultid="12468" />
                    <RANKING order="6" place="-1" resultid="10704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15351" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9914" />
                    <RANKING order="2" place="2" resultid="12373" />
                    <RANKING order="3" place="3" resultid="11714" />
                    <RANKING order="4" place="4" resultid="12891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15352" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10682" />
                    <RANKING order="2" place="2" resultid="9675" />
                    <RANKING order="3" place="3" resultid="11965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15353" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12048" />
                    <RANKING order="2" place="2" resultid="9870" />
                    <RANKING order="3" place="3" resultid="11857" />
                    <RANKING order="4" place="4" resultid="10508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15354" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9564" />
                    <RANKING order="2" place="2" resultid="9332" />
                    <RANKING order="3" place="3" resultid="10412" />
                    <RANKING order="4" place="4" resultid="11065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15355" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10525" />
                    <RANKING order="2" place="2" resultid="10887" />
                    <RANKING order="3" place="3" resultid="8770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15356" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11362" />
                    <RANKING order="2" place="2" resultid="9552" />
                    <RANKING order="3" place="3" resultid="8806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15357" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15358" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15359" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15360" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14303" daytime="17:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14304" daytime="17:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14305" daytime="17:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14306" daytime="17:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14307" daytime="17:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8534" daytime="19:33" gender="F" number="30" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15607" agemax="99" agemin="80" name="80-99" calculate="TOTAL" />
                <AGEGROUP agegroupid="15608" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12925" />
                    <RANKING order="2" place="-1" resultid="12115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15609" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11181" />
                    <RANKING order="2" place="-1" resultid="10085" />
                    <RANKING order="3" place="-1" resultid="9223" />
                    <RANKING order="4" place="-1" resultid="10694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15610" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9931" />
                    <RANKING order="2" place="2" resultid="11904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15611" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9777" />
                    <RANKING order="2" place="-1" resultid="11794" />
                    <RANKING order="3" place="-1" resultid="12040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15612" agemax="279" agemin="240" name="240-279" calculate="TOTAL" />
                <AGEGROUP agegroupid="15613" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9557" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14334" daytime="19:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14335" daytime="19:37" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8566" daytime="19:59" gender="F" number="32" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15406" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11921" />
                    <RANKING order="2" place="-1" resultid="10339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15407" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15408" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10404" />
                    <RANKING order="2" place="2" resultid="10277" />
                    <RANKING order="3" place="-1" resultid="8954" />
                    <RANKING order="4" place="-1" resultid="9212" />
                    <RANKING order="5" place="-1" resultid="11314" />
                    <RANKING order="6" place="-1" resultid="11833" />
                    <RANKING order="7" place="-1" resultid="12071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15409" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11131" />
                    <RANKING order="2" place="-1" resultid="12382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15410" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11037" />
                    <RANKING order="2" place="2" resultid="11007" />
                    <RANKING order="3" place="-1" resultid="11802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15411" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12374" />
                    <RANKING order="2" place="2" resultid="9686" />
                    <RANKING order="3" place="3" resultid="11845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15412" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10656" />
                    <RANKING order="2" place="2" resultid="12785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15413" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12049" />
                    <RANKING order="2" place="2" resultid="11858" />
                    <RANKING order="3" place="3" resultid="11986" />
                    <RANKING order="4" place="4" resultid="9729" />
                    <RANKING order="5" place="-1" resultid="11058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15414" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9764" />
                    <RANKING order="2" place="2" resultid="10873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15415" agemax="69" agemin="65" name="65-69" />
                <AGEGROUP agegroupid="15416" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15417" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15418" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15419" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15420" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14340" daytime="19:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14341" daytime="20:09" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14342" daytime="20:17" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8406" daytime="16:21" gender="M" number="23" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15301" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10332" />
                    <RANKING order="2" place="2" resultid="8975" />
                    <RANKING order="3" place="3" resultid="8988" />
                    <RANKING order="4" place="4" resultid="8925" />
                    <RANKING order="5" place="5" resultid="9362" />
                    <RANKING order="6" place="6" resultid="9117" />
                    <RANKING order="7" place="7" resultid="10609" />
                    <RANKING order="8" place="8" resultid="10737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15302" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8991" />
                    <RANKING order="2" place="2" resultid="9029" />
                    <RANKING order="3" place="3" resultid="9147" />
                    <RANKING order="4" place="4" resultid="10380" />
                    <RANKING order="5" place="5" resultid="10782" />
                    <RANKING order="6" place="6" resultid="10805" />
                    <RANKING order="7" place="7" resultid="10800" />
                    <RANKING order="8" place="8" resultid="12743" />
                    <RANKING order="9" place="-1" resultid="9153" />
                    <RANKING order="10" place="-1" resultid="9454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15303" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9420" />
                    <RANKING order="2" place="2" resultid="10283" />
                    <RANKING order="3" place="3" resultid="11355" />
                    <RANKING order="4" place="4" resultid="10730" />
                    <RANKING order="5" place="5" resultid="12759" />
                    <RANKING order="6" place="6" resultid="9822" />
                    <RANKING order="7" place="7" resultid="9275" />
                    <RANKING order="8" place="-1" resultid="10674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15304" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11945" />
                    <RANKING order="2" place="2" resultid="9906" />
                    <RANKING order="3" place="3" resultid="10043" />
                    <RANKING order="4" place="4" resultid="12859" />
                    <RANKING order="5" place="5" resultid="9982" />
                    <RANKING order="6" place="6" resultid="10065" />
                    <RANKING order="7" place="7" resultid="11879" />
                    <RANKING order="8" place="8" resultid="12419" />
                    <RANKING order="9" place="-1" resultid="10078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15305" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11979" />
                    <RANKING order="2" place="2" resultid="10568" />
                    <RANKING order="3" place="3" resultid="9282" />
                    <RANKING order="4" place="4" resultid="10245" />
                    <RANKING order="5" place="5" resultid="12845" />
                    <RANKING order="6" place="6" resultid="9007" />
                    <RANKING order="7" place="7" resultid="11280" />
                    <RANKING order="8" place="8" resultid="12105" />
                    <RANKING order="9" place="9" resultid="11114" />
                    <RANKING order="10" place="10" resultid="9817" />
                    <RANKING order="11" place="11" resultid="9323" />
                    <RANKING order="12" place="-1" resultid="10663" />
                    <RANKING order="13" place="-1" resultid="11872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15306" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10581" />
                    <RANKING order="2" place="2" resultid="11013" />
                    <RANKING order="3" place="3" resultid="8917" />
                    <RANKING order="4" place="4" resultid="11368" />
                    <RANKING order="5" place="5" resultid="12880" />
                    <RANKING order="6" place="6" resultid="9436" />
                    <RANKING order="7" place="-1" resultid="11126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15307" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9951" />
                    <RANKING order="2" place="2" resultid="11912" />
                    <RANKING order="3" place="3" resultid="11777" />
                    <RANKING order="4" place="4" resultid="12399" />
                    <RANKING order="5" place="5" resultid="10643" />
                    <RANKING order="6" place="6" resultid="9756" />
                    <RANKING order="7" place="7" resultid="8907" />
                    <RANKING order="8" place="8" resultid="9395" />
                    <RANKING order="9" place="9" resultid="9430" />
                    <RANKING order="10" place="10" resultid="11273" />
                    <RANKING order="11" place="-1" resultid="9468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15308" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11199" />
                    <RANKING order="2" place="2" resultid="11768" />
                    <RANKING order="3" place="3" resultid="9882" />
                    <RANKING order="4" place="4" resultid="9740" />
                    <RANKING order="5" place="-1" resultid="12414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15309" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9665" />
                    <RANKING order="2" place="2" resultid="9127" />
                    <RANKING order="3" place="3" resultid="11267" />
                    <RANKING order="4" place="4" resultid="10349" />
                    <RANKING order="5" place="5" resultid="9693" />
                    <RANKING order="6" place="-1" resultid="11756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15310" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11750" />
                    <RANKING order="2" place="2" resultid="11376" />
                    <RANKING order="3" place="3" resultid="10515" />
                    <RANKING order="4" place="4" resultid="11743" />
                    <RANKING order="5" place="-1" resultid="9573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15311" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9834" />
                    <RANKING order="2" place="2" resultid="10444" />
                    <RANKING order="3" place="3" resultid="8822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15312" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9504" />
                    <RANKING order="2" place="2" resultid="8856" />
                    <RANKING order="3" place="3" resultid="10532" />
                    <RANKING order="4" place="4" resultid="11814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15313" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11383" />
                    <RANKING order="2" place="-1" resultid="10432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15314" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9309" />
                    <RANKING order="2" place="2" resultid="9099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15315" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14275" daytime="16:21" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14276" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14277" daytime="16:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14278" daytime="16:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14279" daytime="16:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14280" daytime="16:37" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14281" daytime="16:39" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14282" daytime="16:41" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14283" daytime="16:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14284" daytime="16:46" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8502" daytime="18:12" gender="F" number="28" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15376" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10338" />
                    <RANKING order="2" place="2" resultid="9387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15377" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9197" />
                    <RANKING order="2" place="2" resultid="9341" />
                    <RANKING order="3" place="3" resultid="12796" />
                    <RANKING order="4" place="4" resultid="12776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15378" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10749" />
                    <RANKING order="2" place="2" resultid="12443" />
                    <RANKING order="3" place="3" resultid="12899" />
                    <RANKING order="4" place="4" resultid="10269" />
                    <RANKING order="5" place="5" resultid="12409" />
                    <RANKING order="6" place="6" resultid="10397" />
                    <RANKING order="7" place="7" resultid="11051" />
                    <RANKING order="8" place="8" resultid="12099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15379" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9462" />
                    <RANKING order="2" place="2" resultid="12435" />
                    <RANKING order="3" place="3" resultid="9077" />
                    <RANKING order="4" place="4" resultid="10691" />
                    <RANKING order="5" place="-1" resultid="12381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15380" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11036" />
                    <RANKING order="2" place="2" resultid="10984" />
                    <RANKING order="3" place="3" resultid="11839" />
                    <RANKING order="4" place="4" resultid="10705" />
                    <RANKING order="5" place="5" resultid="11146" />
                    <RANKING order="6" place="6" resultid="12469" />
                    <RANKING order="7" place="7" resultid="10030" />
                    <RANKING order="8" place="8" resultid="9771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15381" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9546" />
                    <RANKING order="2" place="2" resultid="9590" />
                    <RANKING order="3" place="3" resultid="11231" />
                    <RANKING order="4" place="4" resultid="10420" />
                    <RANKING order="5" place="5" resultid="12892" />
                    <RANKING order="6" place="-1" resultid="9681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15382" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12784" />
                    <RANKING order="2" place="2" resultid="11708" />
                    <RANKING order="3" place="3" resultid="10588" />
                    <RANKING order="4" place="-1" resultid="11966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15383" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11702" />
                    <RANKING order="2" place="2" resultid="9703" />
                    <RANKING order="3" place="3" resultid="10864" />
                    <RANKING order="4" place="4" resultid="10509" />
                    <RANKING order="5" place="-1" resultid="11057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15384" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9565" />
                    <RANKING order="2" place="2" resultid="9333" />
                    <RANKING order="3" place="3" resultid="10413" />
                    <RANKING order="4" place="4" resultid="11974" />
                    <RANKING order="5" place="5" resultid="12461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15385" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10651" />
                    <RANKING order="2" place="2" resultid="12014" />
                    <RANKING order="3" place="-1" resultid="11300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15386" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15387" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15388" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15389" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15390" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14316" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14317" daytime="18:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14318" daytime="18:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14319" daytime="18:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14320" daytime="18:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14321" daytime="18:35" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8582" daytime="20:28" gender="M" number="33" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15421" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9630" />
                    <RANKING order="2" place="2" resultid="9118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15422" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12769" />
                    <RANKING order="2" place="2" resultid="10381" />
                    <RANKING order="3" place="3" resultid="9945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15423" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12368" />
                    <RANKING order="2" place="2" resultid="9377" />
                    <RANKING order="3" place="3" resultid="12362" />
                    <RANKING order="4" place="4" resultid="12760" />
                    <RANKING order="5" place="-1" resultid="9829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15424" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12860" />
                    <RANKING order="2" place="2" resultid="10389" />
                    <RANKING order="3" place="3" resultid="10724" />
                    <RANKING order="4" place="4" resultid="10020" />
                    <RANKING order="5" place="-1" resultid="12006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15425" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12838" />
                    <RANKING order="2" place="2" resultid="12906" />
                    <RANKING order="3" place="3" resultid="9165" />
                    <RANKING order="4" place="4" resultid="9623" />
                    <RANKING order="5" place="5" resultid="10998" />
                    <RANKING order="6" place="-1" resultid="9645" />
                    <RANKING order="7" place="-1" resultid="11867" />
                    <RANKING order="8" place="-1" resultid="11938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15426" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9638" />
                    <RANKING order="2" place="2" resultid="8946" />
                    <RANKING order="3" place="3" resultid="11014" />
                    <RANKING order="4" place="4" resultid="9055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15427" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12428" />
                    <RANKING order="2" place="2" resultid="12400" />
                    <RANKING order="3" place="3" resultid="8849" />
                    <RANKING order="4" place="4" resultid="9469" />
                    <RANKING order="5" place="-1" resultid="8908" />
                    <RANKING order="6" place="-1" resultid="11913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15428" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9083" />
                    <RANKING order="2" place="2" resultid="9598" />
                    <RANKING order="3" place="3" resultid="11769" />
                    <RANKING order="4" place="4" resultid="12866" />
                    <RANKING order="5" place="5" resultid="9741" />
                    <RANKING order="6" place="-1" resultid="10092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15429" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9666" />
                    <RANKING order="2" place="2" resultid="10638" />
                    <RANKING order="3" place="3" resultid="11268" />
                    <RANKING order="4" place="4" resultid="9407" />
                    <RANKING order="5" place="5" resultid="9856" />
                    <RANKING order="6" place="-1" resultid="9889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15430" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11751" />
                    <RANKING order="2" place="2" resultid="11377" />
                    <RANKING order="3" place="3" resultid="10520" />
                    <RANKING order="4" place="4" resultid="10453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15431" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11824" />
                    <RANKING order="2" place="2" resultid="9712" />
                    <RANKING order="3" place="3" resultid="10255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15432" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8831" />
                    <RANKING order="2" place="-1" resultid="8886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15433" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15434" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15435" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14343" daytime="20:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14344" daytime="20:39" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14345" daytime="20:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14346" daytime="20:59" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14347" daytime="21:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14348" daytime="21:14" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2018-11-18" daytime="09:00" name="III Blok" number="4" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="8694" daytime="10:55" gender="M" number="39" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15511" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8977" />
                    <RANKING order="2" place="2" resultid="10327" />
                    <RANKING order="3" place="3" resultid="8989" />
                    <RANKING order="4" place="4" resultid="8927" />
                    <RANKING order="5" place="5" resultid="9120" />
                    <RANKING order="6" place="6" resultid="10604" />
                    <RANKING order="7" place="7" resultid="10611" />
                    <RANKING order="8" place="-1" resultid="9024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15512" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8992" />
                    <RANKING order="2" place="2" resultid="9149" />
                    <RANKING order="3" place="3" resultid="9031" />
                    <RANKING order="4" place="4" resultid="10783" />
                    <RANKING order="5" place="5" resultid="9108" />
                    <RANKING order="6" place="6" resultid="12746" />
                    <RANKING order="7" place="-1" resultid="9457" />
                    <RANKING order="8" place="-1" resultid="10801" />
                    <RANKING order="9" place="-1" resultid="10806" />
                    <RANKING order="10" place="-1" resultid="11403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15513" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9422" />
                    <RANKING order="2" place="2" resultid="10284" />
                    <RANKING order="3" place="3" resultid="11357" />
                    <RANKING order="4" place="4" resultid="10731" />
                    <RANKING order="5" place="5" resultid="10293" />
                    <RANKING order="6" place="6" resultid="10676" />
                    <RANKING order="7" place="7" resultid="12762" />
                    <RANKING order="8" place="8" resultid="9278" />
                    <RANKING order="9" place="9" resultid="12094" />
                    <RANKING order="10" place="-1" resultid="10300" />
                    <RANKING order="11" place="-1" resultid="12370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15514" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11947" />
                    <RANKING order="2" place="2" resultid="10045" />
                    <RANKING order="3" place="3" resultid="9909" />
                    <RANKING order="4" place="4" resultid="9985" />
                    <RANKING order="5" place="5" resultid="10371" />
                    <RANKING order="6" place="6" resultid="12861" />
                    <RANKING order="7" place="7" resultid="10067" />
                    <RANKING order="8" place="8" resultid="12080" />
                    <RANKING order="9" place="9" resultid="11881" />
                    <RANKING order="10" place="10" resultid="10022" />
                    <RANKING order="11" place="11" resultid="12421" />
                    <RANKING order="12" place="12" resultid="10079" />
                    <RANKING order="13" place="13" resultid="10056" />
                    <RANKING order="14" place="-1" resultid="11241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15515" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9284" />
                    <RANKING order="2" place="2" resultid="10247" />
                    <RANKING order="3" place="3" resultid="12847" />
                    <RANKING order="4" place="4" resultid="9625" />
                    <RANKING order="5" place="5" resultid="11874" />
                    <RANKING order="6" place="6" resultid="10001" />
                    <RANKING order="7" place="7" resultid="12108" />
                    <RANKING order="8" place="8" resultid="10569" />
                    <RANKING order="9" place="9" resultid="9326" />
                    <RANKING order="10" place="-1" resultid="9616" />
                    <RANKING order="11" place="-1" resultid="10664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15516" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11015" />
                    <RANKING order="2" place="2" resultid="11127" />
                    <RANKING order="3" place="3" resultid="11370" />
                    <RANKING order="4" place="4" resultid="12881" />
                    <RANKING order="5" place="5" resultid="11888" />
                    <RANKING order="6" place="-1" resultid="10583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15517" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10644" />
                    <RANKING order="2" place="2" resultid="11779" />
                    <RANKING order="3" place="3" resultid="9757" />
                    <RANKING order="4" place="4" resultid="12402" />
                    <RANKING order="5" place="5" resultid="8851" />
                    <RANKING order="6" place="6" resultid="8910" />
                    <RANKING order="7" place="7" resultid="9397" />
                    <RANKING order="8" place="8" resultid="11275" />
                    <RANKING order="9" place="-1" resultid="9432" />
                    <RANKING order="10" place="-1" resultid="9471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15518" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11200" />
                    <RANKING order="2" place="2" resultid="9041" />
                    <RANKING order="3" place="3" resultid="11082" />
                    <RANKING order="4" place="4" resultid="11770" />
                    <RANKING order="5" place="5" resultid="9883" />
                    <RANKING order="6" place="6" resultid="9743" />
                    <RANKING order="7" place="-1" resultid="12415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15519" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9668" />
                    <RANKING order="2" place="2" resultid="9130" />
                    <RANKING order="3" place="3" resultid="10350" />
                    <RANKING order="4" place="4" resultid="11269" />
                    <RANKING order="5" place="5" resultid="11757" />
                    <RANKING order="6" place="6" resultid="9696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15520" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11752" />
                    <RANKING order="2" place="2" resultid="11378" />
                    <RANKING order="3" place="3" resultid="13227" />
                    <RANKING order="4" place="4" resultid="9575" />
                    <RANKING order="5" place="5" resultid="11744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15521" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9837" />
                    <RANKING order="2" place="2" resultid="10625" />
                    <RANKING order="3" place="3" resultid="10446" />
                    <RANKING order="4" place="4" resultid="8825" />
                    <RANKING order="5" place="5" resultid="10504" />
                    <RANKING order="6" place="-1" resultid="11739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15522" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8859" />
                    <RANKING order="2" place="2" resultid="9505" />
                    <RANKING order="3" place="3" resultid="10534" />
                    <RANKING order="4" place="4" resultid="11817" />
                    <RANKING order="5" place="5" resultid="9749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15523" agemax="84" agemin="80" name="80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11385" />
                    <RANKING order="2" place="2" resultid="10433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15524" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9311" />
                    <RANKING order="2" place="2" resultid="9101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15525" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14379" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14380" daytime="10:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14381" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14382" daytime="11:01" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14383" daytime="11:03" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14384" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14385" daytime="11:07" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14386" daytime="11:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14387" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14388" daytime="11:11" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14389" daytime="11:13" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8662" daytime="10:07" gender="M" number="37" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15481" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9631" />
                    <RANKING order="2" place="2" resultid="10320" />
                    <RANKING order="3" place="3" resultid="9364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15482" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12771" />
                    <RANKING order="2" place="2" resultid="9496" />
                    <RANKING order="3" place="3" resultid="11325" />
                    <RANKING order="4" place="4" resultid="12745" />
                    <RANKING order="5" place="-1" resultid="9946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15483" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12363" />
                    <RANKING order="2" place="2" resultid="10720" />
                    <RANKING order="3" place="3" resultid="9277" />
                    <RANKING order="4" place="4" resultid="10376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15484" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10665" />
                    <RANKING order="2" place="2" resultid="9879" />
                    <RANKING order="3" place="3" resultid="9984" />
                    <RANKING order="4" place="4" resultid="11254" />
                    <RANKING order="5" place="5" resultid="10390" />
                    <RANKING order="6" place="6" resultid="10370" />
                    <RANKING order="7" place="7" resultid="10561" />
                    <RANKING order="8" place="8" resultid="10021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15485" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9615" />
                    <RANKING order="2" place="2" resultid="11939" />
                    <RANKING order="3" place="3" resultid="12907" />
                    <RANKING order="4" place="4" resultid="9167" />
                    <RANKING order="5" place="5" resultid="10999" />
                    <RANKING order="6" place="6" resultid="12876" />
                    <RANKING order="7" place="-1" resultid="9624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15486" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10478" />
                    <RANKING order="2" place="2" resultid="8919" />
                    <RANKING order="3" place="3" resultid="9053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15487" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13226" />
                    <RANKING order="2" place="2" resultid="11289" />
                    <RANKING order="3" place="3" resultid="11930" />
                    <RANKING order="4" place="4" resultid="11214" />
                    <RANKING order="5" place="5" resultid="9470" />
                    <RANKING order="6" place="-1" resultid="11788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15488" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9599" />
                    <RANKING order="2" place="2" resultid="9529" />
                    <RANKING order="3" place="3" resultid="9092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15489" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9890" />
                    <RANKING order="2" place="2" resultid="10639" />
                    <RANKING order="3" place="3" resultid="9409" />
                    <RANKING order="4" place="4" resultid="9858" />
                    <RANKING order="5" place="5" resultid="9695" />
                    <RANKING order="6" place="6" resultid="9842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15490" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11262" />
                    <RANKING order="2" place="2" resultid="8842" />
                    <RANKING order="3" place="3" resultid="10630" />
                    <RANKING order="4" place="4" resultid="9355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15491" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9836" />
                    <RANKING order="2" place="2" resultid="9541" />
                    <RANKING order="3" place="3" resultid="9735" />
                    <RANKING order="4" place="4" resultid="8824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15492" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8833" />
                    <RANKING order="2" place="2" resultid="10439" />
                    <RANKING order="3" place="3" resultid="11816" />
                    <RANKING order="4" place="4" resultid="8815" />
                    <RANKING order="5" place="-1" resultid="8887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15493" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15494" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15495" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14366" daytime="10:07" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14367" daytime="10:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14368" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14369" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14370" daytime="10:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14371" daytime="10:32" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8710" daytime="11:17" gender="X" number="40" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15621" agemax="99" agemin="80" name="80-99" calculate="TOTAL" />
                <AGEGROUP agegroupid="15622" agemax="119" agemin="100" name="100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12929" />
                    <RANKING order="2" place="2" resultid="11176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15623" agemax="159" agemin="120" name="120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10311" />
                    <RANKING order="2" place="2" resultid="12930" />
                    <RANKING order="3" place="3" resultid="10089" />
                    <RANKING order="4" place="4" resultid="10463" />
                    <RANKING order="5" place="5" resultid="12113" />
                    <RANKING order="6" place="-1" resultid="9225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15624" agemax="199" agemin="160" name="160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9937" />
                    <RANKING order="2" place="2" resultid="11030" />
                    <RANKING order="3" place="3" resultid="11906" />
                    <RANKING order="4" place="-1" resultid="12041" />
                    <RANKING order="5" place="-1" resultid="12454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15625" agemax="239" agemin="200" name="200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9113" />
                    <RANKING order="2" place="2" resultid="9774" />
                    <RANKING order="3" place="3" resultid="12931" />
                    <RANKING order="4" place="4" resultid="11790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15626" agemax="279" agemin="240" name="240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10659" />
                    <RANKING order="2" place="2" resultid="9776" />
                    <RANKING order="3" place="3" resultid="11415" />
                    <RANKING order="4" place="4" resultid="10894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15627" agemax="-1" agemin="280" name="280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9559" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14390" daytime="11:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14391" daytime="11:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14392" daytime="11:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8726" daytime="11:31" gender="F" number="41" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15526" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9389" />
                    <RANKING order="2" place="2" resultid="9895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15527" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9344" />
                    <RANKING order="2" place="2" resultid="12778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15528" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8956" />
                    <RANKING order="2" place="2" resultid="10279" />
                    <RANKING order="3" place="3" resultid="12445" />
                    <RANKING order="4" place="4" resultid="12901" />
                    <RANKING order="5" place="5" resultid="12073" />
                    <RANKING order="6" place="6" resultid="11052" />
                    <RANKING order="7" place="-1" resultid="12411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15529" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9463" />
                    <RANKING order="2" place="2" resultid="9812" />
                    <RANKING order="3" place="3" resultid="12436" />
                    <RANKING order="4" place="4" resultid="9079" />
                    <RANKING order="5" place="5" resultid="10692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15530" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11039" />
                    <RANKING order="2" place="2" resultid="8961" />
                    <RANKING order="3" place="3" resultid="10707" />
                    <RANKING order="4" place="4" resultid="11841" />
                    <RANKING order="5" place="5" resultid="8964" />
                    <RANKING order="6" place="6" resultid="10031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15531" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9548" />
                    <RANKING order="2" place="2" resultid="12376" />
                    <RANKING order="3" place="3" resultid="11233" />
                    <RANKING order="4" place="-1" resultid="10422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15532" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12787" />
                    <RANKING order="2" place="2" resultid="10589" />
                    <RANKING order="3" place="3" resultid="11968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15533" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15637" />
                    <RANKING order="2" place="2" resultid="9705" />
                    <RANKING order="3" place="3" resultid="12051" />
                    <RANKING order="4" place="4" resultid="11860" />
                    <RANKING order="5" place="5" resultid="10511" />
                    <RANKING order="6" place="6" resultid="9731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15534" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9567" />
                    <RANKING order="2" place="2" resultid="10415" />
                    <RANKING order="3" place="3" resultid="11067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15535" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10653" />
                    <RANKING order="2" place="2" resultid="11301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15536" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15537" agemax="79" agemin="75" name="75-79" />
                <AGEGROUP agegroupid="15538" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15539" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15540" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14393" daytime="11:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14394" daytime="11:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14395" daytime="11:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14396" daytime="11:59" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8646" daytime="09:43" gender="F" number="36" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15466" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8998" />
                    <RANKING order="2" place="2" resultid="9894" />
                    <RANKING order="3" place="3" resultid="9388" />
                    <RANKING order="4" place="4" resultid="12752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15467" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="9198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15468" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12444" />
                    <RANKING order="2" place="2" resultid="10270" />
                    <RANKING order="3" place="-1" resultid="9213" />
                    <RANKING order="4" place="-1" resultid="10687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15469" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12831" />
                    <RANKING order="2" place="2" resultid="9078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15470" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9265" />
                    <RANKING order="2" place="2" resultid="11852" />
                    <RANKING order="3" place="3" resultid="12803" />
                    <RANKING order="4" place="4" resultid="12471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15471" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9915" />
                    <RANKING order="2" place="2" resultid="12375" />
                    <RANKING order="3" place="3" resultid="10421" />
                    <RANKING order="4" place="4" resultid="12893" />
                    <RANKING order="5" place="-1" resultid="9688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15472" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12786" />
                    <RANKING order="2" place="2" resultid="11967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15473" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12050" />
                    <RANKING order="2" place="2" resultid="11859" />
                    <RANKING order="3" place="3" resultid="10510" />
                    <RANKING order="4" place="4" resultid="10865" />
                    <RANKING order="5" place="5" resultid="11988" />
                    <RANKING order="6" place="6" resultid="9730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15474" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9566" />
                    <RANKING order="2" place="2" resultid="9766" />
                    <RANKING order="3" place="3" resultid="10414" />
                    <RANKING order="4" place="4" resultid="9335" />
                    <RANKING order="5" place="5" resultid="11066" />
                    <RANKING order="6" place="-1" resultid="11975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15475" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10652" />
                    <RANKING order="2" place="2" resultid="8771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15476" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15477" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15478" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15479" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15480" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14362" daytime="09:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14363" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14364" daytime="09:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14365" daytime="10:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8742" daytime="12:16" gender="M" number="42" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15541" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15635" />
                    <RANKING order="2" place="2" resultid="9632" />
                    <RANKING order="3" place="3" resultid="9365" />
                    <RANKING order="4" place="4" resultid="15633" />
                    <RANKING order="5" place="-1" resultid="8978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15542" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10383" />
                    <RANKING order="2" place="2" resultid="9652" />
                    <RANKING order="3" place="3" resultid="12855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15543" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9317" />
                    <RANKING order="2" place="2" resultid="11329" />
                    <RANKING order="3" place="3" resultid="15629" />
                    <RANKING order="4" place="4" resultid="11358" />
                    <RANKING order="5" place="5" resultid="12095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15544" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11948" />
                    <RANKING order="2" place="2" resultid="11255" />
                    <RANKING order="3" place="3" resultid="12028" />
                    <RANKING order="4" place="4" resultid="10562" />
                    <RANKING order="5" place="5" resultid="12810" />
                    <RANKING order="6" place="-1" resultid="11882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15545" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12840" />
                    <RANKING order="2" place="2" resultid="12908" />
                    <RANKING order="3" place="3" resultid="8934" />
                    <RANKING order="4" place="4" resultid="11940" />
                    <RANKING order="5" place="5" resultid="11343" />
                    <RANKING order="6" place="6" resultid="10570" />
                    <RANKING order="7" place="7" resultid="11000" />
                    <RANKING order="8" place="8" resultid="12877" />
                    <RANKING order="9" place="9" resultid="12452" />
                    <RANKING order="10" place="10" resultid="9259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15546" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10584" />
                    <RANKING order="2" place="2" resultid="9640" />
                    <RANKING order="3" place="3" resultid="10700" />
                    <RANKING order="4" place="4" resultid="15636" />
                    <RANKING order="5" place="5" resultid="8948" />
                    <RANKING order="6" place="6" resultid="8902" />
                    <RANKING order="7" place="7" resultid="11371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15547" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8940" />
                    <RANKING order="2" place="2" resultid="11070" />
                    <RANKING order="3" place="3" resultid="12430" />
                    <RANKING order="4" place="4" resultid="11808" />
                    <RANKING order="5" place="5" resultid="11931" />
                    <RANKING order="6" place="6" resultid="11780" />
                    <RANKING order="7" place="7" resultid="12913" />
                    <RANKING order="8" place="8" resultid="11276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15548" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15631" />
                    <RANKING order="2" place="2" resultid="9600" />
                    <RANKING order="3" place="3" resultid="11771" />
                    <RANKING order="4" place="4" resultid="12868" />
                    <RANKING order="5" place="5" resultid="9402" />
                    <RANKING order="6" place="6" resultid="9093" />
                    <RANKING order="7" place="7" resultid="11763" />
                    <RANKING order="8" place="8" resultid="11296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15549" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8781" />
                    <RANKING order="2" place="2" resultid="12393" />
                    <RANKING order="3" place="3" resultid="10882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15550" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10358" />
                    <RANKING order="2" place="2" resultid="10631" />
                    <RANKING order="3" place="3" resultid="9356" />
                    <RANKING order="4" place="4" resultid="10455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15551" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9714" />
                    <RANKING order="2" place="2" resultid="11826" />
                    <RANKING order="3" place="3" resultid="8796" />
                    <RANKING order="4" place="4" resultid="12792" />
                    <RANKING order="5" place="5" resultid="8878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15552" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11162" />
                    <RANKING order="2" place="2" resultid="15591" />
                    <RANKING order="3" place="3" resultid="8816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15553" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15554" agemax="89" agemin="85" name="85 - 89">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15555" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14398" daytime="12:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14399" daytime="12:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14400" daytime="12:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14401" daytime="12:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14402" daytime="12:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14403" daytime="13:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14404" daytime="13:06" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8630" daytime="09:17" gender="M" number="35" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15451" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10796" />
                    <RANKING order="2" place="2" resultid="10326" />
                    <RANKING order="3" place="3" resultid="10945" />
                    <RANKING order="4" place="4" resultid="10776" />
                    <RANKING order="5" place="5" resultid="10319" />
                    <RANKING order="6" place="6" resultid="12886" />
                    <RANKING order="7" place="7" resultid="10345" />
                    <RANKING order="8" place="-1" resultid="9119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15452" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9477" />
                    <RANKING order="2" place="2" resultid="12770" />
                    <RANKING order="3" place="3" resultid="10951" />
                    <RANKING order="4" place="4" resultid="9651" />
                    <RANKING order="5" place="5" resultid="10382" />
                    <RANKING order="6" place="6" resultid="12854" />
                    <RANKING order="7" place="7" resultid="12022" />
                    <RANKING order="8" place="-1" resultid="9456" />
                    <RANKING order="9" place="-1" resultid="11194" />
                    <RANKING order="10" place="-1" resultid="11402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15453" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9929" />
                    <RANKING order="2" place="2" resultid="12369" />
                    <RANKING order="3" place="3" resultid="10292" />
                    <RANKING order="4" place="4" resultid="10967" />
                    <RANKING order="5" place="5" resultid="9378" />
                    <RANKING order="6" place="6" resultid="12761" />
                    <RANKING order="7" place="7" resultid="10935" />
                    <RANKING order="8" place="-1" resultid="9485" />
                    <RANKING order="9" place="-1" resultid="9958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15454" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10308" />
                    <RANKING order="2" place="2" resultid="10537" />
                    <RANKING order="3" place="3" resultid="9977" />
                    <RANKING order="4" place="4" resultid="12079" />
                    <RANKING order="5" place="5" resultid="11120" />
                    <RANKING order="6" place="6" resultid="12027" />
                    <RANKING order="7" place="7" resultid="10363" />
                    <RANKING order="8" place="8" resultid="10428" />
                    <RANKING order="9" place="-1" resultid="9878" />
                    <RANKING order="10" place="-1" resultid="9908" />
                    <RANKING order="11" place="-1" resultid="10725" />
                    <RANKING order="12" place="-1" resultid="12007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15455" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12839" />
                    <RANKING order="2" place="2" resultid="8933" />
                    <RANKING order="3" place="3" resultid="11953" />
                    <RANKING order="4" place="4" resultid="9166" />
                    <RANKING order="5" place="5" resultid="9993" />
                    <RANKING order="6" place="6" resultid="12107" />
                    <RANKING order="7" place="7" resultid="12451" />
                    <RANKING order="8" place="8" resultid="9325" />
                    <RANKING order="9" place="-1" resultid="9159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15456" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9639" />
                    <RANKING order="2" place="2" resultid="10576" />
                    <RANKING order="3" place="3" resultid="11391" />
                    <RANKING order="4" place="4" resultid="8947" />
                    <RANKING order="5" place="5" resultid="11020" />
                    <RANKING order="6" place="6" resultid="9349" />
                    <RANKING order="7" place="-1" resultid="8901" />
                    <RANKING order="8" place="-1" resultid="11109" />
                    <RANKING order="9" place="-1" resultid="11335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15457" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11069" />
                    <RANKING order="2" place="2" resultid="11288" />
                    <RANKING order="3" place="3" resultid="12401" />
                    <RANKING order="4" place="4" resultid="8850" />
                    <RANKING order="5" place="5" resultid="8909" />
                    <RANKING order="6" place="-1" resultid="12429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15458" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9040" />
                    <RANKING order="2" place="2" resultid="11959" />
                    <RANKING order="3" place="3" resultid="12867" />
                    <RANKING order="4" place="4" resultid="9742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15459" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12821" />
                    <RANKING order="2" place="2" resultid="11206" />
                    <RANKING order="3" place="3" resultid="9667" />
                    <RANKING order="4" place="4" resultid="9129" />
                    <RANKING order="5" place="5" resultid="9415" />
                    <RANKING order="6" place="6" resultid="9857" />
                    <RANKING order="7" place="-1" resultid="9408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15460" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10357" />
                    <RANKING order="2" place="2" resultid="8841" />
                    <RANKING order="3" place="3" resultid="10454" />
                    <RANKING order="4" place="-1" resultid="10521" />
                    <RANKING order="5" place="-1" resultid="11733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15461" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9924" />
                    <RANKING order="2" place="2" resultid="9713" />
                    <RANKING order="3" place="3" resultid="10256" />
                    <RANKING order="4" place="4" resultid="11825" />
                    <RANKING order="5" place="5" resultid="8877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15462" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8858" />
                    <RANKING order="2" place="2" resultid="11161" />
                    <RANKING order="3" place="3" resultid="8832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15463" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15464" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15465" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14353" daytime="09:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14354" daytime="09:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14355" daytime="09:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14356" daytime="09:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14357" daytime="09:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14358" daytime="09:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14359" daytime="09:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14360" daytime="09:36" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14361" daytime="09:38" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8678" daytime="10:39" gender="F" number="38" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15496" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11923" />
                    <RANKING order="2" place="2" resultid="8983" />
                    <RANKING order="3" place="3" resultid="9301" />
                    <RANKING order="4" place="4" resultid="9112" />
                    <RANKING order="5" place="5" resultid="12753" />
                    <RANKING order="6" place="6" resultid="10617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15497" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9012" />
                    <RANKING order="2" place="2" resultid="12797" />
                    <RANKING order="3" place="3" resultid="9343" />
                    <RANKING order="4" place="4" resultid="10962" />
                    <RANKING order="5" place="5" resultid="9491" />
                    <RANKING order="6" place="6" resultid="10745" />
                    <RANKING order="7" place="7" resultid="11352" />
                    <RANKING order="8" place="8" resultid="10670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15498" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10263" />
                    <RANKING order="2" place="2" resultid="10406" />
                    <RANKING order="3" place="3" resultid="10278" />
                    <RANKING order="4" place="4" resultid="11834" />
                    <RANKING order="5" place="5" resultid="10770" />
                    <RANKING order="6" place="6" resultid="12100" />
                    <RANKING order="7" place="-1" resultid="9205" />
                    <RANKING order="8" place="-1" resultid="9214" />
                    <RANKING order="9" place="-1" resultid="13300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15499" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11247" />
                    <RANKING order="2" place="2" resultid="9063" />
                    <RANKING order="3" place="-1" resultid="12383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15500" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9582" />
                    <RANKING order="2" place="2" resultid="11348" />
                    <RANKING order="3" place="3" resultid="13212" />
                    <RANKING order="4" place="4" resultid="8960" />
                    <RANKING order="5" place="5" resultid="11009" />
                    <RANKING order="6" place="6" resultid="9266" />
                    <RANKING order="7" place="7" resultid="10986" />
                    <RANKING order="8" place="8" resultid="12034" />
                    <RANKING order="9" place="9" resultid="11993" />
                    <RANKING order="10" place="-1" resultid="9864" />
                    <RANKING order="11" place="-1" resultid="11840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15501" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9547" />
                    <RANKING order="2" place="2" resultid="11232" />
                    <RANKING order="3" place="3" resultid="11715" />
                    <RANKING order="4" place="4" resultid="9591" />
                    <RANKING order="5" place="5" resultid="11846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15502" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9676" />
                    <RANKING order="2" place="2" resultid="10658" />
                    <RANKING order="3" place="3" resultid="9609" />
                    <RANKING order="4" place="4" resultid="11709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15503" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9872" />
                    <RANKING order="2" place="2" resultid="9043" />
                    <RANKING order="3" place="3" resultid="13295" />
                    <RANKING order="4" place="4" resultid="10866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15504" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11999" />
                    <RANKING order="2" place="2" resultid="11414" />
                    <RANKING order="3" place="3" resultid="10875" />
                    <RANKING order="4" place="4" resultid="11976" />
                    <RANKING order="5" place="5" resultid="12462" />
                    <RANKING order="6" place="-1" resultid="11697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15505" agemax="69" agemin="65" name="65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12015" />
                    <RANKING order="2" place="2" resultid="10526" />
                    <RANKING order="3" place="3" resultid="9516" />
                    <RANKING order="4" place="4" resultid="8772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15506" agemax="74" agemin="70" name="70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9553" />
                    <RANKING order="2" place="2" resultid="9722" />
                    <RANKING order="3" place="3" resultid="8808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15507" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15508" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15509" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15510" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14372" daytime="10:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14373" daytime="10:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14374" daytime="10:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14375" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14376" daytime="10:47" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14377" daytime="10:49" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14378" daytime="10:50" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8613" daytime="09:00" gender="F" number="34" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15436" agemax="24" agemin="20" name="20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11922" />
                    <RANKING order="2" place="2" resultid="12086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15437" agemax="29" agemin="25" name="25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15438" agemax="34" agemin="30" name="30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12900" />
                    <RANKING order="2" place="2" resultid="10405" />
                    <RANKING order="3" place="3" resultid="8955" />
                    <RANKING order="4" place="4" resultid="12072" />
                    <RANKING order="5" place="5" resultid="12410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15439" agemax="39" agemin="35" name="35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10074" />
                    <RANKING order="2" place="2" resultid="12830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15440" agemax="44" agemin="40" name="40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10469" />
                    <RANKING order="2" place="2" resultid="11008" />
                    <RANKING order="3" place="3" resultid="10985" />
                    <RANKING order="4" place="4" resultid="10706" />
                    <RANKING order="5" place="5" resultid="12470" />
                    <RANKING order="6" place="6" resultid="9772" />
                    <RANKING order="7" place="-1" resultid="11038" />
                    <RANKING order="8" place="-1" resultid="11803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15441" agemax="49" agemin="45" name="45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9900" />
                    <RANKING order="2" place="2" resultid="9682" />
                    <RANKING order="3" place="3" resultid="9687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15442" agemax="54" agemin="50" name="50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10657" />
                    <RANKING order="2" place="2" resultid="9608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15443" agemax="59" agemin="55" name="55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9871" />
                    <RANKING order="2" place="2" resultid="9047" />
                    <RANKING order="3" place="3" resultid="9704" />
                    <RANKING order="4" place="4" resultid="11987" />
                    <RANKING order="5" place="-1" resultid="11059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15444" agemax="64" agemin="60" name="60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9765" />
                    <RANKING order="2" place="2" resultid="10874" />
                    <RANKING order="3" place="3" resultid="9334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15445" agemax="69" agemin="65" name="65-69" />
                <AGEGROUP agegroupid="15446" agemax="74" agemin="70" name="70-74" />
                <AGEGROUP agegroupid="15447" agemax="79" agemin="75" name="75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15448" agemax="84" agemin="80" name="80-84" />
                <AGEGROUP agegroupid="15449" agemax="89" agemin="85" name="85 - 89" />
                <AGEGROUP agegroupid="15450" agemax="94" agemin="90" name="90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14349" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14350" daytime="09:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14351" daytime="09:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14352" daytime="09:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="RUS" clubid="9953" name="105th Element Dubna">
          <ATHLETES>
            <ATHLETE birthdate="1986-05-25" firstname="Dmitry" gender="M" lastname="Korobov " nation="POL" athleteid="9954">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9955" heatid="14157" lane="2" entrytime="00:00:26.50" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="9956" heatid="14234" lane="1" entrytime="00:00:59.00" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="9957" heatid="14300" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9958" heatid="14360" lane="9" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="9813" name="5STYL Warszawa">
          <CONTACT name="Korzeniowski" />
          <ATHLETES>
            <ATHLETE birthdate="1977-06-16" firstname="Adrian" gender="M" lastname="Kulisz" nation="POL" athleteid="9814">
              <RESULTS>
                <RESULT eventid="1075" points="421" reactiontime="+99" swimtime="00:00:31.70" resultid="9815" heatid="14149" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="8277" points="412" reactiontime="+94" swimtime="00:01:09.95" resultid="9816" heatid="14227" lane="4" entrytime="00:01:14.00" />
                <RESULT eventid="8406" points="391" reactiontime="+85" swimtime="00:01:29.73" resultid="9817" heatid="14279" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-09" firstname="Paweł" gender="M" lastname="Korzeniowski" nation="POL" athleteid="9823">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1075" points="986" reactiontime="+75" swimtime="00:00:22.23" resultid="9824" heatid="14161" lane="4" entrytime="00:00:22.99" />
                <RESULT eventid="1105" points="944" reactiontime="+78" swimtime="00:02:00.39" resultid="9825" heatid="14174" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.45" />
                    <SPLIT distance="100" swimtime="00:00:57.18" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8277" points="992" reactiontime="+77" swimtime="00:00:49.17" resultid="9826" heatid="14237" lane="5" entrytime="00:00:49.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="1032" reactiontime="+76" swimtime="00:00:54.41" resultid="9827" heatid="14255" lane="4" entrytime="00:00:54.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8454" points="930" swimtime="00:00:23.43" resultid="9828" heatid="14302" lane="4" entrytime="00:00:23.99" />
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="9829" heatid="14348" lane="4" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-02" firstname="Tomasz" gender="M" lastname="Iwańczyk" nation="POL" athleteid="9818">
              <RESULTS>
                <RESULT eventid="1075" points="360" reactiontime="+105" swimtime="00:00:31.10" resultid="9819" heatid="14149" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="8213" points="287" reactiontime="+93" swimtime="00:00:40.14" resultid="9820" heatid="14202" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="8277" points="335" reactiontime="+91" swimtime="00:01:10.57" resultid="9821" heatid="14226" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="430" reactiontime="+88" swimtime="00:01:21.22" resultid="9822" heatid="14277" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8993" name="Akademia WSB w Dąbrowie Górniczej" shortname="AWSB w Dąbrowie Górniczej">
          <ATHLETES>
            <ATHLETE birthdate="1996-05-27" firstname="Monika" gender="F" lastname="Kisiel" nation="POL" athleteid="8994">
              <RESULTS>
                <RESULT eventid="1135" points="558" reactiontime="+85" swimtime="00:11:05.46" resultid="8995" heatid="14178" lane="1" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:01:53.76" />
                    <SPLIT distance="200" swimtime="00:02:34.15" />
                    <SPLIT distance="250" swimtime="00:03:15.02" />
                    <SPLIT distance="300" swimtime="00:03:56.58" />
                    <SPLIT distance="350" swimtime="00:04:38.66" />
                    <SPLIT distance="400" swimtime="00:05:21.23" />
                    <SPLIT distance="450" swimtime="00:06:04.12" />
                    <SPLIT distance="500" swimtime="00:06:47.01" />
                    <SPLIT distance="550" swimtime="00:07:30.53" />
                    <SPLIT distance="600" swimtime="00:08:13.89" />
                    <SPLIT distance="650" swimtime="00:08:56.81" />
                    <SPLIT distance="700" swimtime="00:09:39.99" />
                    <SPLIT distance="750" swimtime="00:10:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="689" reactiontime="+88" swimtime="00:00:33.15" resultid="8996" heatid="14197" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="8470" points="733" reactiontime="+87" swimtime="00:01:11.40" resultid="8997" heatid="14307" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="615" reactiontime="+84" swimtime="00:02:34.91" resultid="8998" heatid="14365" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LAT" clubid="8776" name="Alytus Litwa">
          <ATHLETES>
            <ATHLETE birthdate="1957-08-05" firstname="Sigitas" gender="M" lastname="Katkevicius" nation="LAT" athleteid="8777">
              <RESULTS>
                <RESULT eventid="1105" points="895" reactiontime="+76" swimtime="00:02:42.32" resultid="8778" heatid="14171" lane="8" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:02:02.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="839" reactiontime="+85" swimtime="00:02:55.91" resultid="8779" heatid="14214" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:10.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="829" reactiontime="+103" swimtime="00:02:25.26" resultid="8780" heatid="14327" lane="0" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="813" reactiontime="+88" swimtime="00:05:16.10" resultid="8781" heatid="14401" lane="3" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                    <SPLIT distance="150" swimtime="00:01:56.25" />
                    <SPLIT distance="200" swimtime="00:02:36.44" />
                    <SPLIT distance="250" swimtime="00:03:17.20" />
                    <SPLIT distance="300" swimtime="00:03:58.04" />
                    <SPLIT distance="350" swimtime="00:04:38.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12754" name="AQUASFERA Masters Olsztyn">
          <CONTACT name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="12902">
              <RESULTS>
                <RESULT eventid="8179" points="697" reactiontime="+85" swimtime="00:18:44.45" resultid="12903" heatid="14189" lane="1" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:46.60" />
                    <SPLIT distance="200" swimtime="00:02:23.84" />
                    <SPLIT distance="250" swimtime="00:03:01.40" />
                    <SPLIT distance="300" swimtime="00:03:38.81" />
                    <SPLIT distance="350" swimtime="00:04:16.46" />
                    <SPLIT distance="400" swimtime="00:04:54.42" />
                    <SPLIT distance="450" swimtime="00:05:32.78" />
                    <SPLIT distance="500" swimtime="00:06:10.75" />
                    <SPLIT distance="550" swimtime="00:06:49.00" />
                    <SPLIT distance="600" swimtime="00:07:26.84" />
                    <SPLIT distance="650" swimtime="00:08:05.22" />
                    <SPLIT distance="700" swimtime="00:08:43.30" />
                    <SPLIT distance="750" swimtime="00:09:21.43" />
                    <SPLIT distance="800" swimtime="00:09:59.49" />
                    <SPLIT distance="850" swimtime="00:10:37.65" />
                    <SPLIT distance="900" swimtime="00:11:16.03" />
                    <SPLIT distance="950" swimtime="00:11:54.21" />
                    <SPLIT distance="1000" swimtime="00:12:31.66" />
                    <SPLIT distance="1050" swimtime="00:13:09.37" />
                    <SPLIT distance="1100" swimtime="00:13:47.34" />
                    <SPLIT distance="1150" swimtime="00:14:24.52" />
                    <SPLIT distance="1200" swimtime="00:15:01.97" />
                    <SPLIT distance="1250" swimtime="00:15:40.28" />
                    <SPLIT distance="1300" swimtime="00:16:17.27" />
                    <SPLIT distance="1350" swimtime="00:16:54.65" />
                    <SPLIT distance="1400" swimtime="00:17:32.00" />
                    <SPLIT distance="1450" swimtime="00:18:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="660" reactiontime="+76" swimtime="00:00:59.78" resultid="12904" heatid="14232" lane="3" entrytime="00:01:01.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="607" reactiontime="+61" swimtime="00:02:13.49" resultid="12905" heatid="14323" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:01:02.02" />
                    <SPLIT distance="150" swimtime="00:01:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="556" reactiontime="+77" swimtime="00:05:29.60" resultid="12906" heatid="14347" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:02:01.42" />
                    <SPLIT distance="200" swimtime="00:02:44.24" />
                    <SPLIT distance="250" swimtime="00:03:32.51" />
                    <SPLIT distance="300" swimtime="00:04:20.15" />
                    <SPLIT distance="350" swimtime="00:04:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="585" reactiontime="+74" swimtime="00:02:36.00" resultid="12907" heatid="14366" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="599" reactiontime="+82" swimtime="00:04:45.40" resultid="12908" heatid="14399" lane="3" entrytime="00:04:49.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:45.05" />
                    <SPLIT distance="200" swimtime="00:02:22.04" />
                    <SPLIT distance="250" swimtime="00:02:58.63" />
                    <SPLIT distance="300" swimtime="00:03:35.94" />
                    <SPLIT distance="350" swimtime="00:04:11.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-15" firstname="Mieszko" gender="M" lastname="Palmi-Kukiełko" nation="POL" athleteid="12763">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1105" points="815" reactiontime="+77" swimtime="00:02:09.04" resultid="12764" heatid="14174" lane="5" entrytime="00:02:11.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                    <SPLIT distance="150" swimtime="00:01:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8179" points="837" reactiontime="+82" swimtime="00:17:07.56" resultid="12765" heatid="14189" lane="3" entrytime="00:17:59.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:37.33" />
                    <SPLIT distance="200" swimtime="00:02:11.94" />
                    <SPLIT distance="250" swimtime="00:02:46.87" />
                    <SPLIT distance="300" swimtime="00:03:21.49" />
                    <SPLIT distance="350" swimtime="00:03:56.45" />
                    <SPLIT distance="400" swimtime="00:04:31.49" />
                    <SPLIT distance="450" swimtime="00:05:06.61" />
                    <SPLIT distance="500" swimtime="00:05:41.76" />
                    <SPLIT distance="550" swimtime="00:06:16.54" />
                    <SPLIT distance="600" swimtime="00:06:51.19" />
                    <SPLIT distance="650" swimtime="00:07:25.62" />
                    <SPLIT distance="700" swimtime="00:08:00.13" />
                    <SPLIT distance="750" swimtime="00:08:34.44" />
                    <SPLIT distance="800" swimtime="00:09:08.96" />
                    <SPLIT distance="850" swimtime="00:09:43.08" />
                    <SPLIT distance="900" swimtime="00:10:17.59" />
                    <SPLIT distance="950" swimtime="00:10:52.07" />
                    <SPLIT distance="1000" swimtime="00:11:26.60" />
                    <SPLIT distance="1050" swimtime="00:12:00.75" />
                    <SPLIT distance="1100" swimtime="00:12:34.94" />
                    <SPLIT distance="1150" swimtime="00:13:09.40" />
                    <SPLIT distance="1200" swimtime="00:13:43.93" />
                    <SPLIT distance="1250" swimtime="00:14:18.26" />
                    <SPLIT distance="1300" swimtime="00:14:52.76" />
                    <SPLIT distance="1350" swimtime="00:15:26.66" />
                    <SPLIT distance="1400" swimtime="00:16:00.89" />
                    <SPLIT distance="1450" swimtime="00:16:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="829" reactiontime="+72" swimtime="00:00:58.76" resultid="12766" heatid="14255" lane="8" entrytime="00:00:59.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="882" reactiontime="+79" swimtime="00:02:11.64" resultid="12767" heatid="14262" lane="4" entrytime="00:02:12.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:02.08" />
                    <SPLIT distance="150" swimtime="00:01:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="775" reactiontime="+88" swimtime="00:00:59.90" resultid="12768" heatid="14315" lane="6" entrytime="00:00:59.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8582" points="903" reactiontime="+75" swimtime="00:04:38.89" resultid="12769" heatid="14348" lane="3" entrytime="00:04:50.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                    <SPLIT distance="200" swimtime="00:02:15.87" />
                    <SPLIT distance="250" swimtime="00:02:55.36" />
                    <SPLIT distance="300" swimtime="00:03:35.01" />
                    <SPLIT distance="350" swimtime="00:04:07.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="869" reactiontime="+76" swimtime="00:00:56.50" resultid="12770" heatid="14361" lane="6" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8662" points="748" reactiontime="+78" swimtime="00:02:07.99" resultid="12771" heatid="14371" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:03.30" />
                    <SPLIT distance="150" swimtime="00:01:35.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="12823">
              <RESULTS>
                <RESULT eventid="1058" points="562" reactiontime="+92" swimtime="00:00:32.28" resultid="12824" heatid="14139" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1090" points="499" reactiontime="+90" swimtime="00:03:03.11" resultid="12825" heatid="14164" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                    <SPLIT distance="150" swimtime="00:02:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="588" reactiontime="+94" swimtime="00:00:38.05" resultid="12826" heatid="14196" lane="2" entrytime="00:00:37.50" />
                <RESULT eventid="8261" points="530" reactiontime="+85" swimtime="00:01:11.38" resultid="12827" heatid="14221" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="613" reactiontime="+79" swimtime="00:00:34.60" resultid="12828" heatid="14288" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="8470" points="457" reactiontime="+79" swimtime="00:01:25.57" resultid="12829" heatid="14306" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="387" reactiontime="+77" swimtime="00:01:29.43" resultid="12830" heatid="14351" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="456" reactiontime="+97" swimtime="00:03:05.43" resultid="12831" heatid="14365" lane="9" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:30.79" />
                    <SPLIT distance="150" swimtime="00:02:19.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-10-03" firstname="Bartosz" gender="M" lastname="Wolak" nation="POL" athleteid="12882">
              <RESULTS>
                <RESULT eventid="1075" points="675" reactiontime="+73" swimtime="00:00:26.15" resultid="12883" heatid="14157" lane="6" entrytime="00:00:26.34" />
                <RESULT eventid="8277" points="636" reactiontime="+80" swimtime="00:00:58.89" resultid="12884" heatid="14235" lane="2" entrytime="00:00:57.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="648" reactiontime="+73" swimtime="00:00:28.61" resultid="12885" heatid="14298" lane="6" entrytime="00:00:29.44" />
                <RESULT eventid="8630" points="562" reactiontime="+72" swimtime="00:01:05.79" resultid="12886" heatid="14359" lane="8" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Zaleska" nation="POL" athleteid="12894">
              <RESULTS>
                <RESULT eventid="1165" points="592" reactiontime="+82" swimtime="00:21:55.33" resultid="12895" heatid="14187" lane="7" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:19.86" />
                    <SPLIT distance="150" swimtime="00:02:02.69" />
                    <SPLIT distance="200" swimtime="00:02:46.08" />
                    <SPLIT distance="250" swimtime="00:03:29.50" />
                    <SPLIT distance="300" swimtime="00:04:12.54" />
                    <SPLIT distance="350" swimtime="00:04:56.07" />
                    <SPLIT distance="400" swimtime="00:05:39.53" />
                    <SPLIT distance="450" swimtime="00:06:23.20" />
                    <SPLIT distance="500" swimtime="00:07:07.12" />
                    <SPLIT distance="550" swimtime="00:07:50.97" />
                    <SPLIT distance="600" swimtime="00:08:34.81" />
                    <SPLIT distance="650" swimtime="00:09:18.72" />
                    <SPLIT distance="700" swimtime="00:10:03.16" />
                    <SPLIT distance="750" swimtime="00:10:47.63" />
                    <SPLIT distance="800" swimtime="00:11:31.83" />
                    <SPLIT distance="850" swimtime="00:12:16.43" />
                    <SPLIT distance="900" swimtime="00:13:01.03" />
                    <SPLIT distance="950" swimtime="00:13:45.91" />
                    <SPLIT distance="1000" swimtime="00:14:30.50" />
                    <SPLIT distance="1050" swimtime="00:15:15.26" />
                    <SPLIT distance="1100" swimtime="00:16:00.19" />
                    <SPLIT distance="1150" swimtime="00:16:44.26" />
                    <SPLIT distance="1200" swimtime="00:17:28.68" />
                    <SPLIT distance="1250" swimtime="00:18:13.14" />
                    <SPLIT distance="1300" swimtime="00:18:58.84" />
                    <SPLIT distance="1350" swimtime="00:19:43.74" />
                    <SPLIT distance="1400" swimtime="00:20:28.35" />
                    <SPLIT distance="1450" swimtime="00:21:12.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="553" reactiontime="+86" swimtime="00:00:36.97" resultid="12896" heatid="14195" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="8325" points="601" reactiontime="+82" swimtime="00:02:49.43" resultid="12897" heatid="14257" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="591" reactiontime="+87" swimtime="00:00:33.58" resultid="12898" heatid="14288" lane="6" entrytime="00:00:34.99" />
                <RESULT eventid="8502" points="545" reactiontime="+98" swimtime="00:02:34.11" resultid="12899" heatid="14320" lane="6" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="628" reactiontime="+86" swimtime="00:01:14.48" resultid="12900" heatid="14352" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="585" reactiontime="+78" swimtime="00:05:26.99" resultid="12901" heatid="14394" lane="3" entrytime="00:05:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:01.48" />
                    <SPLIT distance="200" swimtime="00:02:43.56" />
                    <SPLIT distance="250" swimtime="00:03:25.27" />
                    <SPLIT distance="300" swimtime="00:04:07.28" />
                    <SPLIT distance="350" swimtime="00:04:48.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="12755">
              <RESULTS>
                <RESULT eventid="1105" points="380" reactiontime="+90" swimtime="00:02:43.06" resultid="12756" heatid="14170" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="512" reactiontime="+72" swimtime="00:02:55.60" resultid="12757" heatid="14216" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:07.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="445" reactiontime="+82" swimtime="00:02:42.37" resultid="12758" heatid="14260" lane="4" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="463" reactiontime="+74" swimtime="00:01:19.26" resultid="12759" heatid="14281" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="441" reactiontime="+88" swimtime="00:05:50.58" resultid="12760" heatid="14343" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:52.66" />
                    <SPLIT distance="200" swimtime="00:03:41.16" />
                    <SPLIT distance="250" swimtime="00:04:30.43" />
                    <SPLIT distance="300" swimtime="00:05:10.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="384" reactiontime="+78" swimtime="00:01:12.38" resultid="12761" heatid="14358" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="423" reactiontime="+71" swimtime="00:00:37.03" resultid="12762" heatid="14386" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-18" firstname="Jacek" gender="M" lastname="Łuczak" nation="POL" athleteid="12843">
              <RESULTS>
                <RESULT eventid="1075" points="610" reactiontime="+76" swimtime="00:00:28.01" resultid="12844" heatid="14151" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="8406" points="565" reactiontime="+78" swimtime="00:01:19.37" resultid="12845" heatid="14278" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="497" reactiontime="+91" swimtime="00:00:31.71" resultid="12846" heatid="14295" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="8694" points="603" reactiontime="+69" swimtime="00:00:34.89" resultid="12847" heatid="14385" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-18" firstname="Danuta" gender="F" lastname="Wegen" nation="POL" athleteid="12887">
              <RESULTS>
                <RESULT eventid="1058" points="172" reactiontime="+127" swimtime="00:00:49.05" resultid="12888" heatid="14134" lane="3" />
                <RESULT eventid="8196" points="180" reactiontime="+99" swimtime="00:00:54.55" resultid="12889" heatid="14193" lane="9" />
                <RESULT eventid="8261" points="155" reactiontime="+101" swimtime="00:01:50.96" resultid="12890" heatid="14218" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="205" reactiontime="+105" swimtime="00:01:58.57" resultid="12891" heatid="14303" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="141" reactiontime="+113" swimtime="00:04:10.33" resultid="12892" heatid="14316" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.24" />
                    <SPLIT distance="100" swimtime="00:01:59.94" />
                    <SPLIT distance="150" swimtime="00:03:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="216" reactiontime="+93" swimtime="00:04:15.99" resultid="12893" heatid="14362" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.42" />
                    <SPLIT distance="100" swimtime="00:02:05.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="12798">
              <RESULTS>
                <RESULT eventid="1058" points="474" reactiontime="+91" swimtime="00:00:34.86" resultid="12799" heatid="14137" lane="2" entrytime="00:00:36.79" />
                <RESULT eventid="8196" points="515" reactiontime="+83" swimtime="00:00:38.09" resultid="12800" heatid="14195" lane="3" entrytime="00:00:40.19" />
                <RESULT eventid="8293" points="471" reactiontime="+79" swimtime="00:01:27.55" resultid="12801" heatid="14240" lane="7" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="512" reactiontime="+73" swimtime="00:01:24.91" resultid="12802" heatid="14305" lane="6" entrytime="00:01:35.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="425" reactiontime="+78" swimtime="00:03:18.66" resultid="12803" heatid="14362" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="12779">
              <RESULTS>
                <RESULT eventid="1090" points="533" swimtime="00:03:11.49" resultid="12780" heatid="14163" lane="5" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="150" swimtime="00:02:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="658" reactiontime="+97" swimtime="00:22:06.16" resultid="12781" heatid="14187" lane="2" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:07.55" />
                    <SPLIT distance="200" swimtime="00:02:51.24" />
                    <SPLIT distance="250" swimtime="00:03:35.00" />
                    <SPLIT distance="300" swimtime="00:04:18.69" />
                    <SPLIT distance="350" swimtime="00:05:02.22" />
                    <SPLIT distance="400" swimtime="00:05:45.89" />
                    <SPLIT distance="450" swimtime="00:06:29.52" />
                    <SPLIT distance="500" swimtime="00:07:14.19" />
                    <SPLIT distance="550" swimtime="00:07:58.58" />
                    <SPLIT distance="600" swimtime="00:08:42.72" />
                    <SPLIT distance="650" swimtime="00:09:27.37" />
                    <SPLIT distance="700" swimtime="00:10:11.72" />
                    <SPLIT distance="750" swimtime="00:10:56.31" />
                    <SPLIT distance="800" swimtime="00:11:40.60" />
                    <SPLIT distance="850" swimtime="00:12:25.20" />
                    <SPLIT distance="900" swimtime="00:13:09.91" />
                    <SPLIT distance="950" swimtime="00:13:55.10" />
                    <SPLIT distance="1000" swimtime="00:14:40.12" />
                    <SPLIT distance="1050" swimtime="00:15:24.94" />
                    <SPLIT distance="1100" swimtime="00:16:09.97" />
                    <SPLIT distance="1150" swimtime="00:16:54.79" />
                    <SPLIT distance="1200" swimtime="00:17:39.75" />
                    <SPLIT distance="1250" swimtime="00:18:24.47" />
                    <SPLIT distance="1300" swimtime="00:19:08.82" />
                    <SPLIT distance="1350" swimtime="00:19:53.11" />
                    <SPLIT distance="1400" swimtime="00:20:37.35" />
                    <SPLIT distance="1450" swimtime="00:21:22.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="552" swimtime="00:03:36.32" resultid="12782" heatid="14209" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                    <SPLIT distance="100" swimtime="00:01:45.27" />
                    <SPLIT distance="150" swimtime="00:02:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="561" reactiontime="+80" swimtime="00:01:15.12" resultid="12783" heatid="14221" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="591" reactiontime="+100" swimtime="00:02:40.66" resultid="12784" heatid="14317" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="489" reactiontime="+101" swimtime="00:07:01.61" resultid="12785" heatid="14341" lane="6" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                    <SPLIT distance="100" swimtime="00:01:48.26" />
                    <SPLIT distance="150" swimtime="00:03:38.73" />
                    <SPLIT distance="200" swimtime="00:04:35.40" />
                    <SPLIT distance="250" swimtime="00:05:33.26" />
                    <SPLIT distance="300" swimtime="00:06:17.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="440" reactiontime="+97" swimtime="00:03:26.96" resultid="12786" heatid="14363" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                    <SPLIT distance="100" swimtime="00:01:40.51" />
                    <SPLIT distance="150" swimtime="00:02:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="585" reactiontime="+91" swimtime="00:05:42.39" resultid="12787" heatid="14393" lane="0" entrytime="00:05:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:22.25" />
                    <SPLIT distance="150" swimtime="00:02:06.06" />
                    <SPLIT distance="200" swimtime="00:02:50.29" />
                    <SPLIT distance="250" swimtime="00:03:34.23" />
                    <SPLIT distance="300" swimtime="00:04:18.10" />
                    <SPLIT distance="350" swimtime="00:05:01.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="12869">
              <RESULTS>
                <RESULT eventid="1075" points="366" reactiontime="+83" swimtime="00:00:33.21" resultid="12870" heatid="14147" lane="2" entrytime="00:00:33.92" />
                <RESULT eventid="1150" points="417" reactiontime="+104" swimtime="00:11:24.39" resultid="12871" heatid="14185" lane="4" entrytime="00:12:17.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                    <SPLIT distance="200" swimtime="00:02:43.63" />
                    <SPLIT distance="250" swimtime="00:03:26.97" />
                    <SPLIT distance="300" swimtime="00:04:10.33" />
                    <SPLIT distance="350" swimtime="00:04:54.32" />
                    <SPLIT distance="400" swimtime="00:05:38.22" />
                    <SPLIT distance="450" swimtime="00:06:21.88" />
                    <SPLIT distance="500" swimtime="00:07:05.12" />
                    <SPLIT distance="550" swimtime="00:07:48.82" />
                    <SPLIT distance="600" swimtime="00:08:32.59" />
                    <SPLIT distance="650" swimtime="00:09:16.11" />
                    <SPLIT distance="700" swimtime="00:10:00.16" />
                    <SPLIT distance="750" swimtime="00:10:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="282" reactiontime="+82" swimtime="00:00:41.36" resultid="12872" heatid="14201" lane="1" entrytime="00:00:44.03" />
                <RESULT eventid="8277" points="352" reactiontime="+82" swimtime="00:01:13.68" resultid="12873" heatid="14227" lane="8" entrytime="00:01:15.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="288" reactiontime="+82" swimtime="00:00:38.05" resultid="12874" heatid="14292" lane="6" entrytime="00:00:41.06" />
                <RESULT eventid="8518" points="380" reactiontime="+104" swimtime="00:02:35.95" resultid="12875" heatid="14326" lane="0" entrytime="00:02:54.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:55.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="316" reactiontime="+75" swimtime="00:03:11.48" resultid="12876" heatid="14368" lane="8" entrytime="00:03:34.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="391" reactiontime="+90" swimtime="00:05:28.96" resultid="12877" heatid="14402" lane="3" entrytime="00:06:03.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:01:59.20" />
                    <SPLIT distance="200" swimtime="00:02:40.72" />
                    <SPLIT distance="250" swimtime="00:03:23.51" />
                    <SPLIT distance="300" swimtime="00:04:06.16" />
                    <SPLIT distance="350" swimtime="00:04:47.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-01" firstname="Adam" gender="M" lastname="Szmit" nation="POL" athleteid="12909">
              <RESULTS>
                <RESULT eventid="8277" points="446" reactiontime="+106" swimtime="00:01:13.86" resultid="12911" heatid="14228" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="455" reactiontime="+112" swimtime="00:02:41.85" resultid="12912" heatid="14327" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:16.95" />
                    <SPLIT distance="150" swimtime="00:02:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="456" reactiontime="+106" swimtime="00:05:38.40" resultid="12913" heatid="14401" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="200" swimtime="00:02:46.23" />
                    <SPLIT distance="350" swimtime="00:04:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="418" reactiontime="+104" swimtime="00:22:40.66" resultid="13205" heatid="14190" lane="8" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:05:50.51" />
                    <SPLIT distance="200" swimtime="00:11:54.74" />
                    <SPLIT distance="250" swimtime="00:14:14.33" />
                    <SPLIT distance="450" swimtime="00:15:46.40" />
                    <SPLIT distance="500" swimtime="00:18:06.49" />
                    <SPLIT distance="550" swimtime="00:18:52.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-18" firstname="Bogdan" gender="M" lastname="Milewski" nation="POL" athleteid="12878">
              <RESULTS>
                <RESULT eventid="8309" points="385" reactiontime="+92" swimtime="00:01:22.57" resultid="12879" heatid="14248" lane="1" entrytime="00:01:20.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="424" reactiontime="+86" swimtime="00:01:27.91" resultid="12880" heatid="14279" lane="5" entrytime="00:01:28.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="473" reactiontime="+80" swimtime="00:00:38.97" resultid="12881" heatid="14384" lane="8" entrytime="00:00:38.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="12804">
              <RESULTS>
                <RESULT eventid="1075" points="513" reactiontime="+82" swimtime="00:00:28.72" resultid="12805" heatid="14152" lane="7" entrytime="00:00:29.00" />
                <RESULT comment="przekroczony limit czasu" eventid="8179" reactiontime="+140" status="DSQ" swimtime="00:22:47.55" resultid="12806" heatid="14191" lane="5" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:22.98" />
                    <SPLIT distance="150" swimtime="00:02:07.01" />
                    <SPLIT distance="200" swimtime="00:02:50.94" />
                    <SPLIT distance="250" swimtime="00:03:36.84" />
                    <SPLIT distance="300" swimtime="00:04:22.21" />
                    <SPLIT distance="350" swimtime="00:05:07.76" />
                    <SPLIT distance="400" swimtime="00:05:53.54" />
                    <SPLIT distance="450" swimtime="00:07:25.92" />
                    <SPLIT distance="500" swimtime="00:08:13.06" />
                    <SPLIT distance="550" swimtime="00:08:59.76" />
                    <SPLIT distance="600" swimtime="00:09:45.69" />
                    <SPLIT distance="650" swimtime="00:10:31.68" />
                    <SPLIT distance="700" swimtime="00:11:18.08" />
                    <SPLIT distance="750" swimtime="00:12:03.31" />
                    <SPLIT distance="800" swimtime="00:12:49.83" />
                    <SPLIT distance="850" swimtime="00:13:36.26" />
                    <SPLIT distance="900" swimtime="00:14:22.62" />
                    <SPLIT distance="950" swimtime="00:15:09.58" />
                    <SPLIT distance="1000" swimtime="00:15:56.35" />
                    <SPLIT distance="1050" swimtime="00:16:43.06" />
                    <SPLIT distance="1100" swimtime="00:17:29.63" />
                    <SPLIT distance="1150" swimtime="00:18:16.83" />
                    <SPLIT distance="1200" swimtime="00:19:02.93" />
                    <SPLIT distance="1250" swimtime="00:19:48.50" />
                    <SPLIT distance="1300" swimtime="00:20:33.92" />
                    <SPLIT distance="1350" swimtime="00:22:03.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="528" reactiontime="+98" swimtime="00:01:03.62" resultid="12807" heatid="14231" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" reactiontime="+121" status="DNS" swimtime="00:00:00.00" resultid="12808" heatid="14292" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="8518" points="409" reactiontime="+123" swimtime="00:02:30.10" resultid="12809" heatid="14329" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="389" reactiontime="+100" swimtime="00:05:31.96" resultid="12810" heatid="14401" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="150" swimtime="00:01:56.93" />
                    <SPLIT distance="200" swimtime="00:02:40.28" />
                    <SPLIT distance="250" swimtime="00:03:24.22" />
                    <SPLIT distance="300" swimtime="00:04:08.03" />
                    <SPLIT distance="350" swimtime="00:04:51.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="12841">
              <RESULTS>
                <RESULT eventid="1150" points="433" reactiontime="+89" swimtime="00:11:26.66" resultid="12842" heatid="14184" lane="9" entrytime="00:12:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:04.10" />
                    <SPLIT distance="200" swimtime="00:02:47.80" />
                    <SPLIT distance="250" swimtime="00:03:31.31" />
                    <SPLIT distance="300" swimtime="00:04:14.84" />
                    <SPLIT distance="350" swimtime="00:04:58.62" />
                    <SPLIT distance="400" swimtime="00:05:42.56" />
                    <SPLIT distance="450" swimtime="00:06:26.48" />
                    <SPLIT distance="500" swimtime="00:07:10.75" />
                    <SPLIT distance="550" swimtime="00:07:55.09" />
                    <SPLIT distance="600" swimtime="00:08:38.06" />
                    <SPLIT distance="650" swimtime="00:09:21.05" />
                    <SPLIT distance="700" swimtime="00:10:03.54" />
                    <SPLIT distance="750" swimtime="00:10:46.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="12832">
              <RESULTS>
                <RESULT eventid="1105" points="724" reactiontime="+87" swimtime="00:02:22.39" resultid="12833" heatid="14173" lane="4" entrytime="00:02:23.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="757" reactiontime="+94" swimtime="00:09:21.38" resultid="12834" heatid="14182" lane="3" entrytime="00:09:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:06.45" />
                    <SPLIT distance="150" swimtime="00:01:41.48" />
                    <SPLIT distance="200" swimtime="00:02:16.95" />
                    <SPLIT distance="250" swimtime="00:02:52.37" />
                    <SPLIT distance="300" swimtime="00:03:27.78" />
                    <SPLIT distance="350" swimtime="00:04:03.30" />
                    <SPLIT distance="400" swimtime="00:04:38.69" />
                    <SPLIT distance="450" swimtime="00:05:14.26" />
                    <SPLIT distance="500" swimtime="00:05:49.88" />
                    <SPLIT distance="550" swimtime="00:06:25.71" />
                    <SPLIT distance="600" swimtime="00:07:01.20" />
                    <SPLIT distance="650" swimtime="00:07:36.61" />
                    <SPLIT distance="700" swimtime="00:08:11.81" />
                    <SPLIT distance="750" swimtime="00:08:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="816" reactiontime="+74" swimtime="00:00:55.71" resultid="12835" heatid="14236" lane="8" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="780" reactiontime="+75" swimtime="00:01:04.98" resultid="12836" heatid="14252" lane="5" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="743" reactiontime="+85" swimtime="00:02:04.75" resultid="12837" heatid="14333" lane="1" entrytime="00:02:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="150" swimtime="00:01:34.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="633" reactiontime="+92" swimtime="00:05:15.63" resultid="12838" heatid="14348" lane="1" entrytime="00:05:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                    <SPLIT distance="150" swimtime="00:01:53.87" />
                    <SPLIT distance="200" swimtime="00:02:35.22" />
                    <SPLIT distance="250" swimtime="00:03:19.76" />
                    <SPLIT distance="300" swimtime="00:04:04.72" />
                    <SPLIT distance="350" swimtime="00:04:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="773" reactiontime="+72" swimtime="00:01:01.68" resultid="12839" heatid="14359" lane="6" entrytime="00:01:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="730" reactiontime="+79" swimtime="00:04:27.17" resultid="12840" heatid="14398" lane="8" entrytime="00:04:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:38.09" />
                    <SPLIT distance="200" swimtime="00:02:12.11" />
                    <SPLIT distance="250" swimtime="00:02:46.16" />
                    <SPLIT distance="300" swimtime="00:03:20.42" />
                    <SPLIT distance="350" swimtime="00:03:54.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-19" firstname="Anna" gender="F" lastname="Głowacka" nation="POL" athleteid="12811">
              <RESULTS>
                <RESULT eventid="1058" points="278" reactiontime="+99" swimtime="00:00:40.78" resultid="12812" heatid="14136" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="8196" points="357" reactiontime="+74" swimtime="00:00:44.92" resultid="12813" heatid="14194" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-08" firstname="Justyna" gender="F" lastname="Łagowska" nation="POL" athleteid="12914">
              <RESULTS>
                <RESULT eventid="1058" points="282" reactiontime="+104" swimtime="00:00:40.60" resultid="12915" heatid="14134" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-06-18" firstname="Monika" gender="F" lastname="Pielowska" nation="POL" athleteid="12793">
              <RESULTS>
                <RESULT eventid="1058" points="809" reactiontime="+73" swimtime="00:00:27.63" resultid="12794" heatid="14141" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="12795" heatid="14223" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="8502" points="895" reactiontime="+76" swimtime="00:02:09.72" resultid="12796" heatid="14321" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.63" />
                    <SPLIT distance="150" swimtime="00:01:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="773" reactiontime="+66" swimtime="00:00:34.42" resultid="12797" heatid="14378" lane="5" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Zdzisław" gender="M" lastname="Choroszewski" nation="POL" athleteid="12788">
              <RESULTS>
                <RESULT eventid="1075" points="349" reactiontime="+102" swimtime="00:00:41.16" resultid="12789" heatid="14144" lane="3" entrytime="00:00:42.10" />
                <RESULT eventid="1150" points="329" reactiontime="+105" swimtime="00:16:36.19" resultid="12790" heatid="14186" lane="2" entrytime="00:16:53.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                    <SPLIT distance="100" swimtime="00:01:51.92" />
                    <SPLIT distance="150" swimtime="00:02:52.49" />
                    <SPLIT distance="200" swimtime="00:03:54.68" />
                    <SPLIT distance="250" swimtime="00:04:58.95" />
                    <SPLIT distance="300" swimtime="00:06:01.43" />
                    <SPLIT distance="350" swimtime="00:07:06.64" />
                    <SPLIT distance="400" swimtime="00:08:10.97" />
                    <SPLIT distance="450" swimtime="00:09:13.12" />
                    <SPLIT distance="500" swimtime="00:10:17.46" />
                    <SPLIT distance="550" swimtime="00:11:23.50" />
                    <SPLIT distance="600" swimtime="00:12:27.86" />
                    <SPLIT distance="650" swimtime="00:13:32.29" />
                    <SPLIT distance="700" swimtime="00:14:35.27" />
                    <SPLIT distance="750" swimtime="00:15:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="288" reactiontime="+83" swimtime="00:03:48.01" resultid="12791" heatid="14323" lane="4" entrytime="00:03:56.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                    <SPLIT distance="100" swimtime="00:01:44.42" />
                    <SPLIT distance="150" swimtime="00:02:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="343" reactiontime="+98" swimtime="00:07:58.15" resultid="12792" heatid="14403" lane="9" entrytime="00:08:34.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.10" />
                    <SPLIT distance="100" swimtime="00:01:49.50" />
                    <SPLIT distance="150" swimtime="00:02:50.12" />
                    <SPLIT distance="200" swimtime="00:03:52.21" />
                    <SPLIT distance="250" swimtime="00:04:54.91" />
                    <SPLIT distance="300" swimtime="00:05:58.05" />
                    <SPLIT distance="350" swimtime="00:06:59.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-28" firstname="Maciej" gender="M" lastname="Zembrzuski" nation="POL" athleteid="12848">
              <RESULTS>
                <RESULT eventid="1105" points="554" reactiontime="+94" swimtime="00:02:26.79" resultid="12849" heatid="14172" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="575" reactiontime="+96" swimtime="00:10:18.83" resultid="12850" heatid="14182" lane="1" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                    <SPLIT distance="200" swimtime="00:02:25.86" />
                    <SPLIT distance="250" swimtime="00:03:03.65" />
                    <SPLIT distance="300" swimtime="00:03:41.70" />
                    <SPLIT distance="350" swimtime="00:04:20.40" />
                    <SPLIT distance="400" swimtime="00:04:59.35" />
                    <SPLIT distance="450" swimtime="00:05:38.21" />
                    <SPLIT distance="500" swimtime="00:06:17.76" />
                    <SPLIT distance="550" swimtime="00:06:57.59" />
                    <SPLIT distance="600" swimtime="00:07:37.64" />
                    <SPLIT distance="650" swimtime="00:08:18.40" />
                    <SPLIT distance="700" swimtime="00:08:59.20" />
                    <SPLIT distance="750" swimtime="00:09:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="686" reactiontime="+87" swimtime="00:00:55.06" resultid="12851" heatid="14237" lane="0" entrytime="00:00:54.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="783" reactiontime="+49" swimtime="00:00:25.71" resultid="12852" heatid="14302" lane="0" entrytime="00:00:25.87" />
                <RESULT eventid="8518" points="723" reactiontime="+86" swimtime="00:02:05.37" resultid="12853" heatid="14332" lane="4" entrytime="00:02:05.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:01.15" />
                    <SPLIT distance="150" swimtime="00:01:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="690" reactiontime="+81" swimtime="00:01:01.02" resultid="12854" heatid="14361" lane="1" entrytime="00:00:58.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="643" reactiontime="+81" swimtime="00:04:43.10" resultid="12855" heatid="14399" lane="2" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:07.97" />
                    <SPLIT distance="150" swimtime="00:01:43.61" />
                    <SPLIT distance="200" swimtime="00:02:19.60" />
                    <SPLIT distance="250" swimtime="00:02:55.47" />
                    <SPLIT distance="300" swimtime="00:03:32.04" />
                    <SPLIT distance="350" swimtime="00:04:08.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-15" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="12856">
              <RESULTS>
                <RESULT eventid="1075" points="666" reactiontime="+73" swimtime="00:00:26.33" resultid="12857" heatid="14153" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="8245" points="710" reactiontime="+84" swimtime="00:02:37.59" resultid="12858" heatid="14217" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:56.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="712" reactiontime="+73" swimtime="00:01:11.69" resultid="12859" heatid="14282" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="567" reactiontime="+75" swimtime="00:05:29.69" resultid="12860" heatid="14346" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:02:44.13" />
                    <SPLIT distance="250" swimtime="00:03:27.09" />
                    <SPLIT distance="300" swimtime="00:04:11.33" />
                    <SPLIT distance="350" swimtime="00:04:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="655" reactiontime="+79" swimtime="00:00:33.24" resultid="12861" heatid="14387" lane="9" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-01" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="12862">
              <RESULTS>
                <RESULT eventid="1150" points="563" reactiontime="+113" swimtime="00:11:52.77" resultid="12863" heatid="14185" lane="2" entrytime="00:12:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                    <SPLIT distance="200" swimtime="00:02:49.64" />
                    <SPLIT distance="250" swimtime="00:03:34.25" />
                    <SPLIT distance="300" swimtime="00:04:19.18" />
                    <SPLIT distance="350" swimtime="00:05:04.45" />
                    <SPLIT distance="400" swimtime="00:05:49.70" />
                    <SPLIT distance="450" swimtime="00:06:35.03" />
                    <SPLIT distance="500" swimtime="00:07:20.82" />
                    <SPLIT distance="550" swimtime="00:08:06.38" />
                    <SPLIT distance="600" swimtime="00:08:52.01" />
                    <SPLIT distance="650" swimtime="00:09:37.24" />
                    <SPLIT distance="700" swimtime="00:10:23.00" />
                    <SPLIT distance="750" swimtime="00:11:08.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="579" reactiontime="+95" swimtime="00:03:14.33" resultid="12864" heatid="14214" lane="7" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="505" reactiontime="+104" swimtime="00:01:22.58" resultid="12865" heatid="14247" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="530" reactiontime="+103" swimtime="00:06:38.69" resultid="12866" heatid="14345" lane="7" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:39.41" />
                    <SPLIT distance="150" swimtime="00:02:33.59" />
                    <SPLIT distance="200" swimtime="00:03:28.07" />
                    <SPLIT distance="250" swimtime="00:04:20.55" />
                    <SPLIT distance="300" swimtime="00:05:13.74" />
                    <SPLIT distance="350" swimtime="00:05:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="353" reactiontime="+92" swimtime="00:01:31.62" resultid="12867" heatid="14355" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="535" reactiontime="+89" swimtime="00:05:49.15" resultid="12868" heatid="14402" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                    <SPLIT distance="200" swimtime="00:02:48.67" />
                    <SPLIT distance="250" swimtime="00:03:34.10" />
                    <SPLIT distance="300" swimtime="00:04:19.99" />
                    <SPLIT distance="350" swimtime="00:05:05.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-15" firstname="Patryk" gender="M" lastname="Poniatowski" nation="POL" athleteid="12916">
              <RESULTS>
                <RESULT comment="M5 - Pływak nie przeniósł ramion do przodu nad lustrem wody." eventid="8454" reactiontime="+69" status="DSQ" swimtime="00:00:24.18" resultid="12917" heatid="14300" lane="8" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="12814">
              <RESULTS>
                <RESULT eventid="1075" points="814" reactiontime="+92" swimtime="00:00:28.74" resultid="12815" heatid="14152" lane="5" entrytime="00:00:28.90" />
                <RESULT eventid="1105" points="1012" reactiontime="+87" swimtime="00:02:35.79" resultid="12816" heatid="14171" lane="6" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:59.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="876" reactiontime="+100" swimtime="00:00:33.22" resultid="12817" heatid="14204" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="8341" points="861" reactiontime="+94" swimtime="00:02:47.89" resultid="12818" heatid="14261" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="794" reactiontime="+87" swimtime="00:00:31.48" resultid="12819" heatid="14295" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="8518" points="924" reactiontime="+96" swimtime="00:02:20.10" resultid="12820" heatid="14329" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="873" reactiontime="+87" swimtime="00:01:10.51" resultid="12821" heatid="14358" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Oriana" gender="F" lastname="Lewandowska" nation="POL" athleteid="12772">
              <RESULTS>
                <RESULT eventid="1135" points="805" reactiontime="+93" swimtime="00:09:58.21" resultid="12773" heatid="14178" lane="4" entrytime="00:09:58.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                    <SPLIT distance="200" swimtime="00:02:30.23" />
                    <SPLIT distance="250" swimtime="00:03:08.53" />
                    <SPLIT distance="300" swimtime="00:03:46.40" />
                    <SPLIT distance="350" swimtime="00:04:24.30" />
                    <SPLIT distance="400" swimtime="00:05:02.02" />
                    <SPLIT distance="450" swimtime="00:05:38.72" />
                    <SPLIT distance="500" swimtime="00:06:15.47" />
                    <SPLIT distance="550" swimtime="00:06:53.10" />
                    <SPLIT distance="600" swimtime="00:07:30.75" />
                    <SPLIT distance="650" swimtime="00:08:08.57" />
                    <SPLIT distance="700" swimtime="00:08:46.24" />
                    <SPLIT distance="750" swimtime="00:09:23.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="891" reactiontime="+84" swimtime="00:02:23.24" resultid="12774" heatid="14257" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="719" reactiontime="+68" swimtime="00:00:31.32" resultid="12775" heatid="14289" lane="9" entrytime="00:00:33.50" />
                <RESULT eventid="8502" points="687" reactiontime="+101" swimtime="00:02:21.69" resultid="12776" heatid="14321" lane="2" entrytime="00:02:19.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="737" reactiontime="+81" swimtime="00:01:08.11" resultid="12777" heatid="14352" lane="4" entrytime="00:01:09.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="749" reactiontime="+85" swimtime="00:04:54.84" resultid="12778" heatid="14393" lane="5" entrytime="00:04:48.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:50.31" />
                    <SPLIT distance="200" swimtime="00:02:28.23" />
                    <SPLIT distance="250" swimtime="00:03:05.47" />
                    <SPLIT distance="300" swimtime="00:03:42.71" />
                    <SPLIT distance="350" swimtime="00:04:19.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-28" firstname="Dawid" gender="M" lastname="Zieja" nation="POL" athleteid="12918">
              <RESULTS>
                <RESULT eventid="1075" points="782" reactiontime="+75" swimtime="00:00:24.79" resultid="12919" heatid="14160" lane="9" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="HARPAGANY" number="4">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+79" swimtime="00:01:50.66" resultid="12920" heatid="14268" lane="2" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:26.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12763" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="12856" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="12848" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="12918" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="BESTIE" number="5">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+93" swimtime="00:02:08.74" resultid="12924" heatid="14266" lane="4" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:37.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12814" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="12843" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="12832" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="12862" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="ORŁY" number="7">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="8550" reactiontime="+73" swimtime="00:01:36.09" resultid="12926" heatid="14339" lane="6" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.58" />
                    <SPLIT distance="100" swimtime="00:00:48.45" />
                    <SPLIT distance="150" swimtime="00:01:12.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12916" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="12848" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="12918" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="12763" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="SOKOŁY" number="8">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+80" swimtime="00:01:46.77" resultid="12927" heatid="14338" lane="5" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="100" swimtime="00:00:53.42" />
                    <SPLIT distance="150" swimtime="00:01:21.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12902" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="12856" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="12843" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="12832" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="HEROSY" number="9">
              <RESULTS>
                <RESULT eventid="8550" swimtime="00:02:01.59" resultid="12928" heatid="14337" lane="3" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:01.04" />
                    <SPLIT distance="150" swimtime="00:01:32.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12814" number="1" />
                    <RELAYPOSITION athleteid="12878" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="12862" number="3" reactiontime="+198" />
                    <RELAYPOSITION athleteid="12804" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="SENIORITY" number="3">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+95" swimtime="00:02:14.00" resultid="12922" heatid="14264" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12894" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="12793" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="12772" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="12823" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="BABY NIEPRUSKIE" number="6">
              <RESULTS>
                <RESULT eventid="8534" reactiontime="+71" swimtime="00:02:02.70" resultid="12925" heatid="14335" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                    <SPLIT distance="150" swimtime="00:01:30.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12793" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="12772" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="12823" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="12894" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="SMERFY" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+77" swimtime="00:01:57.87" resultid="12921" heatid="14177" lane="9" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                    <SPLIT distance="100" swimtime="00:00:50.82" />
                    <SPLIT distance="150" swimtime="00:01:23.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12918" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="12832" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="12823" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="12779" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="GUMISIE" number="3">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+86" swimtime="00:01:47.69" resultid="12923" heatid="14177" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="100" swimtime="00:00:50.60" />
                    <SPLIT distance="150" swimtime="00:01:17.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12848" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="12763" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="12793" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="12772" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="MALAGA" number="10">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="8710" reactiontime="+67" swimtime="00:01:56.67" resultid="12929" heatid="14392" lane="4" entrytime="00:01:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.97" />
                    <SPLIT distance="100" swimtime="00:01:01.13" />
                    <SPLIT distance="150" swimtime="00:01:32.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12763" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="12793" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="12772" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="12918" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="TIKI TAKI" number="11">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+68" swimtime="00:02:05.72" resultid="12930" heatid="14392" lane="7" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="100" swimtime="00:01:00.19" />
                    <SPLIT distance="150" swimtime="00:01:33.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12916" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="12856" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="12894" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="12823" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="KASZTANKI" number="12">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+84" swimtime="00:02:21.93" resultid="12931" heatid="14391" lane="8" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:47.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12798" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="12878" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="12814" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="12779" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="POM" clubid="10240" name="AquaStars Gdynia">
          <CONTACT email="mariuszgolon5@wp.pl" name="Mariusz Golon" phone="609649755" />
          <ATHLETES>
            <ATHLETE birthdate="1978-11-20" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="10241">
              <RESULTS>
                <RESULT eventid="1075" points="691" reactiontime="+89" swimtime="00:00:26.87" resultid="10242" heatid="14150" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="8213" points="605" reactiontime="+86" swimtime="00:00:32.10" resultid="10243" heatid="14202" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="8309" points="684" reactiontime="+83" swimtime="00:01:07.87" resultid="10244" heatid="14250" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="617" reactiontime="+91" swimtime="00:01:17.08" resultid="10245" heatid="14276" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="672" reactiontime="+88" swimtime="00:00:28.68" resultid="10246" heatid="14297" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="8694" points="693" reactiontime="+82" swimtime="00:00:33.32" resultid="10247" heatid="14383" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="9094" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóraa" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" license="100611700315" athleteid="9095">
              <RESULTS>
                <RESULT eventid="8179" reactiontime="+89" swimtime="00:45:22.06" resultid="9096" heatid="14191" lane="7" entrytime="00:44:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.13" />
                    <SPLIT distance="100" swimtime="00:02:51.47" />
                    <SPLIT distance="150" swimtime="00:04:21.01" />
                    <SPLIT distance="200" swimtime="00:05:49.18" />
                    <SPLIT distance="250" swimtime="00:07:17.44" />
                    <SPLIT distance="300" swimtime="00:08:46.26" />
                    <SPLIT distance="350" swimtime="00:10:18.25" />
                    <SPLIT distance="400" swimtime="00:11:49.98" />
                    <SPLIT distance="450" swimtime="00:13:23.41" />
                    <SPLIT distance="500" swimtime="00:14:56.87" />
                    <SPLIT distance="550" swimtime="00:16:31.40" />
                    <SPLIT distance="600" swimtime="00:18:05.77" />
                    <SPLIT distance="650" swimtime="00:19:37.89" />
                    <SPLIT distance="700" swimtime="00:21:12.53" />
                    <SPLIT distance="750" swimtime="00:22:50.53" />
                    <SPLIT distance="800" swimtime="00:24:25.84" />
                    <SPLIT distance="850" swimtime="00:26:01.97" />
                    <SPLIT distance="900" swimtime="00:27:39.69" />
                    <SPLIT distance="950" swimtime="00:29:18.82" />
                    <SPLIT distance="1000" swimtime="00:30:54.63" />
                    <SPLIT distance="1050" swimtime="00:32:30.75" />
                    <SPLIT distance="1100" swimtime="00:34:09.19" />
                    <SPLIT distance="1150" swimtime="00:35:46.61" />
                    <SPLIT distance="1200" swimtime="00:37:25.09" />
                    <SPLIT distance="1250" swimtime="00:39:01.49" />
                    <SPLIT distance="1300" swimtime="00:40:36.56" />
                    <SPLIT distance="1350" swimtime="00:42:11.65" />
                    <SPLIT distance="1400" swimtime="00:43:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="328" swimtime="00:06:09.53" resultid="9097" heatid="14212" lane="0" entrytime="00:05:23.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.80" />
                    <SPLIT distance="100" swimtime="00:03:07.26" />
                    <SPLIT distance="150" swimtime="00:04:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="198" reactiontime="+100" swimtime="00:02:29.36" resultid="9098" heatid="14224" lane="3" entrytime="00:02:30.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="214" reactiontime="+110" swimtime="00:02:53.15" resultid="9099" heatid="14275" lane="4" entrytime="00:02:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="204" reactiontime="+149" swimtime="00:05:30.69" resultid="9100" heatid="14323" lane="7" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.83" />
                    <SPLIT distance="100" swimtime="00:02:45.87" />
                    <SPLIT distance="150" swimtime="00:04:11.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="226" reactiontime="+111" swimtime="00:01:17.97" resultid="9101" heatid="14380" lane="0" entrytime="00:01:08.57" />
                <RESULT eventid="8742" points="291" reactiontime="+149" swimtime="00:11:15.79" resultid="9102" heatid="14404" lane="6" entrytime="00:10:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.56" />
                    <SPLIT distance="100" swimtime="00:02:43.36" />
                    <SPLIT distance="150" swimtime="00:04:12.77" />
                    <SPLIT distance="200" swimtime="00:05:37.54" />
                    <SPLIT distance="250" swimtime="00:07:05.62" />
                    <SPLIT distance="300" swimtime="00:08:32.35" />
                    <SPLIT distance="350" swimtime="00:09:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="213" reactiontime="+95" swimtime="00:01:04.96" resultid="9302" heatid="14143" lane="1" entrytime="00:01:00.21" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9103" name="AZS KU UW">
          <CONTACT city="Warszawa" email="mbaranowski@fuw.edu.pl" internet="http://www.azs.uw.edu.pl/" name="Baranowski Marek" state="MAZ" street="ul. Dobra 56/66, p. 162" zip="00-312" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" athleteid="9104">
              <RESULTS>
                <RESULT eventid="1075" points="712" reactiontime="+73" swimtime="00:00:25.57" resultid="9105" heatid="14158" lane="5" entrytime="00:00:25.80" entrycourse="SCM" />
                <RESULT eventid="8277" points="706" reactiontime="+72" swimtime="00:00:54.54" resultid="9106" heatid="14236" lane="3" entrytime="00:00:55.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="764" reactiontime="+72" swimtime="00:02:03.08" resultid="9107" heatid="14333" lane="6" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="100" swimtime="00:00:57.43" />
                    <SPLIT distance="150" swimtime="00:01:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="666" reactiontime="+73" swimtime="00:00:32.36" resultid="9108" heatid="14388" lane="9" entrytime="00:00:33.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-08-27" firstname="Edyta" gender="F" lastname="Ilcewicz" nation="POL" athleteid="9109">
              <RESULTS>
                <RESULT eventid="8293" points="706" reactiontime="+69" swimtime="00:01:10.94" resultid="9110" heatid="14243" lane="8" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="705" reactiontime="+81" swimtime="00:01:19.47" resultid="9111" heatid="14274" lane="1" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="697" reactiontime="+73" swimtime="00:00:37.03" resultid="9112" heatid="14378" lane="0" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS PWSZ R" nation="POL" region="SLA" clubid="9660" name="AZS PWSZ Racibórz">
          <CONTACT city="Raciborz" email="adip45@poczta.onet.pl" name="PIECHULA" state="ŚLA" street="SŁOWACKIEGO" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-11-04" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="9661">
              <RESULTS>
                <RESULT eventid="1105" points="644" reactiontime="+106" swimtime="00:03:01.10" resultid="9662" heatid="14169" lane="3" entrytime="00:03:09.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:17.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="577" reactiontime="+110" swimtime="00:03:19.24" resultid="9663" heatid="14214" lane="1" entrytime="00:03:21.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:35.51" />
                    <SPLIT distance="150" swimtime="00:02:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="514" reactiontime="+93" swimtime="00:03:19.37" resultid="9664" heatid="14260" lane="9" entrytime="00:03:20.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:34.88" />
                    <SPLIT distance="150" swimtime="00:02:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="584" reactiontime="+100" swimtime="00:01:28.35" resultid="9665" heatid="14278" lane="4" entrytime="00:01:30.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="612" reactiontime="+100" swimtime="00:06:39.86" resultid="9666" heatid="14345" lane="6" entrytime="00:06:45.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:35.97" />
                    <SPLIT distance="150" swimtime="00:02:28.95" />
                    <SPLIT distance="200" swimtime="00:03:20.48" />
                    <SPLIT distance="250" swimtime="00:04:16.47" />
                    <SPLIT distance="300" swimtime="00:05:12.36" />
                    <SPLIT distance="350" swimtime="00:05:58.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="447" reactiontime="+91" swimtime="00:01:28.14" resultid="9667" heatid="14356" lane="1" entrytime="00:01:24.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="576" reactiontime="+85" swimtime="00:00:39.33" resultid="9668" heatid="14383" lane="7" entrytime="00:00:40.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10695" name="CityZen Poznań">
          <CONTACT city="Daszewice" email="gmo@o2.pl" name="MONCZAK, Grzegorz" phone="608639696" zip="61-160" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-05" firstname="Kinga" gender="F" lastname="Jaruga" nation="POL" athleteid="10701">
              <RESULTS>
                <RESULT eventid="1165" points="535" reactiontime="+110" swimtime="00:22:59.91" resultid="10702" heatid="14187" lane="1" entrytime="00:23:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:09.67" />
                    <SPLIT distance="200" swimtime="00:02:55.15" />
                    <SPLIT distance="250" swimtime="00:03:40.82" />
                    <SPLIT distance="300" swimtime="00:04:26.68" />
                    <SPLIT distance="350" swimtime="00:05:12.49" />
                    <SPLIT distance="400" swimtime="00:05:58.66" />
                    <SPLIT distance="450" swimtime="00:06:44.99" />
                    <SPLIT distance="500" swimtime="00:07:31.52" />
                    <SPLIT distance="550" swimtime="00:08:17.84" />
                    <SPLIT distance="600" swimtime="00:09:04.39" />
                    <SPLIT distance="650" swimtime="00:09:50.86" />
                    <SPLIT distance="700" swimtime="00:10:37.56" />
                    <SPLIT distance="750" swimtime="00:11:24.24" />
                    <SPLIT distance="800" swimtime="00:12:10.83" />
                    <SPLIT distance="850" swimtime="00:12:57.56" />
                    <SPLIT distance="900" swimtime="00:13:44.18" />
                    <SPLIT distance="950" swimtime="00:14:30.77" />
                    <SPLIT distance="1000" swimtime="00:15:17.70" />
                    <SPLIT distance="1050" swimtime="00:16:04.05" />
                    <SPLIT distance="1100" swimtime="00:16:50.65" />
                    <SPLIT distance="1150" swimtime="00:17:37.10" />
                    <SPLIT distance="1200" swimtime="00:18:23.76" />
                    <SPLIT distance="1250" swimtime="00:19:09.95" />
                    <SPLIT distance="1300" swimtime="00:19:56.89" />
                    <SPLIT distance="1350" swimtime="00:20:43.54" />
                    <SPLIT distance="1400" swimtime="00:21:29.73" />
                    <SPLIT distance="1450" swimtime="00:22:15.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="315" reactiontime="+100" swimtime="00:03:36.92" resultid="10703" heatid="14257" lane="1" entrytime="00:03:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="100" swimtime="00:01:42.02" />
                    <SPLIT distance="150" swimtime="00:02:39.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" status="DNS" swimtime="00:00:00.00" resultid="10704" heatid="14305" lane="4" entrytime="00:01:29.99" entrycourse="SCM" />
                <RESULT eventid="8502" points="446" reactiontime="+95" swimtime="00:02:49.17" resultid="10705" heatid="14320" lane="9" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:21.23" />
                    <SPLIT distance="150" swimtime="00:02:06.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="353" reactiontime="+71" swimtime="00:01:33.47" resultid="10706" heatid="14351" lane="7" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="502" reactiontime="+92" swimtime="00:05:48.37" resultid="10707" heatid="14395" lane="6" entrytime="00:06:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                    <SPLIT distance="200" swimtime="00:02:51.66" />
                    <SPLIT distance="250" swimtime="00:03:36.46" />
                    <SPLIT distance="300" swimtime="00:04:21.81" />
                    <SPLIT distance="350" swimtime="00:05:05.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="10696">
              <RESULTS>
                <RESULT eventid="8179" points="721" reactiontime="+93" swimtime="00:18:22.04" resultid="10697" heatid="14189" lane="2" entrytime="00:18:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:44.90" />
                    <SPLIT distance="200" swimtime="00:02:21.50" />
                    <SPLIT distance="250" swimtime="00:02:58.31" />
                    <SPLIT distance="300" swimtime="00:03:34.68" />
                    <SPLIT distance="350" swimtime="00:04:11.23" />
                    <SPLIT distance="400" swimtime="00:04:48.16" />
                    <SPLIT distance="450" swimtime="00:05:24.79" />
                    <SPLIT distance="500" swimtime="00:06:01.65" />
                    <SPLIT distance="550" swimtime="00:06:38.47" />
                    <SPLIT distance="600" swimtime="00:07:15.39" />
                    <SPLIT distance="650" swimtime="00:07:52.35" />
                    <SPLIT distance="700" swimtime="00:08:29.46" />
                    <SPLIT distance="750" swimtime="00:09:06.41" />
                    <SPLIT distance="800" swimtime="00:09:43.46" />
                    <SPLIT distance="850" swimtime="00:10:20.73" />
                    <SPLIT distance="900" swimtime="00:10:57.56" />
                    <SPLIT distance="950" swimtime="00:11:34.78" />
                    <SPLIT distance="1000" swimtime="00:12:12.08" />
                    <SPLIT distance="1050" swimtime="00:12:49.33" />
                    <SPLIT distance="1100" swimtime="00:13:26.58" />
                    <SPLIT distance="1150" swimtime="00:14:03.82" />
                    <SPLIT distance="1200" swimtime="00:14:41.33" />
                    <SPLIT distance="1250" swimtime="00:15:18.38" />
                    <SPLIT distance="1300" swimtime="00:15:55.51" />
                    <SPLIT distance="1350" swimtime="00:16:32.63" />
                    <SPLIT distance="1400" swimtime="00:17:09.53" />
                    <SPLIT distance="1450" swimtime="00:17:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="680" reactiontime="+80" swimtime="00:01:00.16" resultid="10698" heatid="14234" lane="8" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="689" reactiontime="+78" swimtime="00:02:09.89" resultid="10699" heatid="14331" lane="5" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="150" swimtime="00:01:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="688" reactiontime="+81" swimtime="00:04:38.51" resultid="10700" heatid="14398" lane="0" entrytime="00:04:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:41.59" />
                    <SPLIT distance="200" swimtime="00:02:17.42" />
                    <SPLIT distance="250" swimtime="00:02:52.98" />
                    <SPLIT distance="300" swimtime="00:03:28.70" />
                    <SPLIT distance="350" swimtime="00:04:03.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GBR" clubid="8928" name="Concept Swimming Club">
          <CONTACT city="London" email="info@conceptswimming.com" name="Bartlomiej Kulaga" phone="+447783308258" street="35 Croftongate Way" zip="SE4 2DL" />
          <ATHLETES>
            <ATHLETE birthdate="1978-03-09" firstname="Aleksandra" gender="F" lastname="Morkisz" nation="GBR" athleteid="8957">
              <RESULTS>
                <RESULT eventid="8229" points="640" reactiontime="+95" swimtime="00:03:12.68" resultid="8958" heatid="14210" lane="4" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:32.58" />
                    <SPLIT distance="150" swimtime="00:02:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="595" reactiontime="+84" swimtime="00:01:29.95" resultid="8959" heatid="14273" lane="8" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="552" reactiontime="+88" swimtime="00:00:41.85" resultid="8960" heatid="14376" lane="1" entrytime="00:00:40.30" />
                <RESULT eventid="8726" points="537" reactiontime="+99" swimtime="00:05:40.62" resultid="8961" heatid="14393" lane="8" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:02:01.52" />
                    <SPLIT distance="200" swimtime="00:02:45.43" />
                    <SPLIT distance="250" swimtime="00:03:29.66" />
                    <SPLIT distance="300" swimtime="00:04:13.94" />
                    <SPLIT distance="350" swimtime="00:04:58.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-07-05" firstname="Peter" gender="M" lastname="Dixon" nation="GBR" athleteid="8935">
              <RESULTS>
                <RESULT eventid="1150" points="957" reactiontime="+88" swimtime="00:09:05.46" resultid="8936" heatid="14182" lane="6" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                    <SPLIT distance="150" swimtime="00:01:35.98" />
                    <SPLIT distance="200" swimtime="00:02:10.22" />
                    <SPLIT distance="250" swimtime="00:02:44.77" />
                    <SPLIT distance="300" swimtime="00:03:19.38" />
                    <SPLIT distance="350" swimtime="00:03:54.32" />
                    <SPLIT distance="400" swimtime="00:04:29.23" />
                    <SPLIT distance="450" swimtime="00:05:04.18" />
                    <SPLIT distance="500" swimtime="00:05:38.86" />
                    <SPLIT distance="550" swimtime="00:06:13.77" />
                    <SPLIT distance="600" swimtime="00:06:48.52" />
                    <SPLIT distance="650" swimtime="00:07:23.04" />
                    <SPLIT distance="700" swimtime="00:07:57.68" />
                    <SPLIT distance="750" swimtime="00:08:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="1000" reactiontime="+90" swimtime="00:00:56.44" resultid="8937" heatid="14235" lane="4" entrytime="00:00:57.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="833" reactiontime="+81" swimtime="00:02:27.63" resultid="8938" heatid="14262" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="983" reactiontime="+98" swimtime="00:02:05.27" resultid="8939" heatid="14333" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:01:01.00" />
                    <SPLIT distance="150" swimtime="00:01:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="965" reactiontime="+79" swimtime="00:04:23.53" resultid="8940" heatid="14398" lane="7" entrytime="00:04:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="150" swimtime="00:01:36.43" />
                    <SPLIT distance="200" swimtime="00:02:09.86" />
                    <SPLIT distance="250" swimtime="00:02:43.13" />
                    <SPLIT distance="300" swimtime="00:03:17.14" />
                    <SPLIT distance="350" swimtime="00:03:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="931" reactiontime="+88" swimtime="00:00:26.02" resultid="10726" heatid="14157" lane="4" entrytime="00:00:26.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-10" firstname="Christopher" gender="M" lastname="Morgan" nation="GBR" athleteid="8941">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="8942" heatid="14172" lane="3" entrytime="00:02:32.00" />
                <RESULT eventid="1150" points="686" reactiontime="+89" swimtime="00:09:49.38" resultid="8943" heatid="14182" lane="7" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:08.07" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                    <SPLIT distance="200" swimtime="00:02:21.38" />
                    <SPLIT distance="250" swimtime="00:02:58.43" />
                    <SPLIT distance="300" swimtime="00:03:35.03" />
                    <SPLIT distance="350" swimtime="00:04:12.17" />
                    <SPLIT distance="400" swimtime="00:04:49.69" />
                    <SPLIT distance="450" swimtime="00:05:26.87" />
                    <SPLIT distance="500" swimtime="00:06:04.12" />
                    <SPLIT distance="550" swimtime="00:06:42.07" />
                    <SPLIT distance="600" swimtime="00:07:19.94" />
                    <SPLIT distance="650" swimtime="00:07:57.78" />
                    <SPLIT distance="700" swimtime="00:08:35.70" />
                    <SPLIT distance="750" swimtime="00:09:13.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="680" reactiontime="+91" swimtime="00:02:47.89" resultid="8944" heatid="14217" lane="0" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="652" reactiontime="+78" swimtime="00:02:31.78" resultid="8945" heatid="14261" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="743" reactiontime="+69" swimtime="00:05:19.09" resultid="8946" heatid="14348" lane="8" entrytime="00:05:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:54.79" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="250" swimtime="00:03:21.83" />
                    <SPLIT distance="300" swimtime="00:04:06.38" />
                    <SPLIT distance="350" swimtime="00:04:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="641" reactiontime="+77" swimtime="00:01:08.17" resultid="8947" heatid="14359" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="507" reactiontime="+84" swimtime="00:05:08.33" resultid="8948" heatid="14398" lane="9" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:49.41" />
                    <SPLIT distance="200" swimtime="00:02:29.28" />
                    <SPLIT distance="250" swimtime="00:03:08.83" />
                    <SPLIT distance="300" swimtime="00:03:48.99" />
                    <SPLIT distance="350" swimtime="00:04:29.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-21" firstname="Lee" gender="F" lastname="Griffin" nation="GBR" athleteid="8962">
              <RESULTS>
                <RESULT comment="przekroczony limit czasu" eventid="1165" reactiontime="+111" status="DSQ" swimtime="00:29:13.24" resultid="8963" heatid="14188" lane="3" entrytime="00:26:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                    <SPLIT distance="100" swimtime="00:01:47.91" />
                    <SPLIT distance="150" swimtime="00:02:45.69" />
                    <SPLIT distance="200" swimtime="00:03:43.39" />
                    <SPLIT distance="250" swimtime="00:04:41.87" />
                    <SPLIT distance="300" swimtime="00:05:40.28" />
                    <SPLIT distance="350" swimtime="00:06:38.36" />
                    <SPLIT distance="400" swimtime="00:07:36.74" />
                    <SPLIT distance="450" swimtime="00:08:35.24" />
                    <SPLIT distance="500" swimtime="00:09:33.39" />
                    <SPLIT distance="550" swimtime="00:10:32.38" />
                    <SPLIT distance="600" swimtime="00:11:30.50" />
                    <SPLIT distance="650" swimtime="00:12:29.42" />
                    <SPLIT distance="700" swimtime="00:13:28.34" />
                    <SPLIT distance="750" swimtime="00:14:27.51" />
                    <SPLIT distance="800" swimtime="00:15:26.47" />
                    <SPLIT distance="850" swimtime="00:16:25.22" />
                    <SPLIT distance="900" swimtime="00:17:24.50" />
                    <SPLIT distance="950" swimtime="00:18:23.86" />
                    <SPLIT distance="1000" swimtime="00:19:22.95" />
                    <SPLIT distance="1050" swimtime="00:20:22.30" />
                    <SPLIT distance="1100" swimtime="00:21:22.54" />
                    <SPLIT distance="1150" swimtime="00:22:21.31" />
                    <SPLIT distance="1200" swimtime="00:23:21.14" />
                    <SPLIT distance="1250" swimtime="00:24:20.84" />
                    <SPLIT distance="1300" swimtime="00:25:20.26" />
                    <SPLIT distance="1350" swimtime="00:26:19.37" />
                    <SPLIT distance="1400" swimtime="00:27:18.09" />
                    <SPLIT distance="1450" swimtime="00:28:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="345" reactiontime="+111" swimtime="00:06:34.54" resultid="8964" heatid="14395" lane="9" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:44.47" />
                    <SPLIT distance="150" swimtime="00:02:42.57" />
                    <SPLIT distance="200" swimtime="00:03:41.10" />
                    <SPLIT distance="250" swimtime="00:04:39.14" />
                    <SPLIT distance="300" swimtime="00:05:36.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-08" firstname="Bartlomiej" gender="M" lastname="Kulaga" nation="GBR" athleteid="8929">
              <RESULTS>
                <RESULT eventid="8179" points="664" reactiontime="+94" swimtime="00:19:02.37" resultid="8930" heatid="14189" lane="0" entrytime="00:19:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:42.26" />
                    <SPLIT distance="200" swimtime="00:02:18.73" />
                    <SPLIT distance="250" swimtime="00:02:55.67" />
                    <SPLIT distance="300" swimtime="00:03:33.26" />
                    <SPLIT distance="350" swimtime="00:04:10.62" />
                    <SPLIT distance="400" swimtime="00:04:48.31" />
                    <SPLIT distance="450" swimtime="00:05:26.13" />
                    <SPLIT distance="500" swimtime="00:06:03.57" />
                    <SPLIT distance="550" swimtime="00:06:41.41" />
                    <SPLIT distance="600" swimtime="00:07:19.91" />
                    <SPLIT distance="650" swimtime="00:07:58.43" />
                    <SPLIT distance="700" swimtime="00:08:36.92" />
                    <SPLIT distance="750" swimtime="00:09:15.60" />
                    <SPLIT distance="800" swimtime="00:09:53.95" />
                    <SPLIT distance="850" swimtime="00:10:32.47" />
                    <SPLIT distance="900" swimtime="00:11:11.95" />
                    <SPLIT distance="950" swimtime="00:11:51.13" />
                    <SPLIT distance="1000" swimtime="00:12:30.27" />
                    <SPLIT distance="1050" swimtime="00:13:09.32" />
                    <SPLIT distance="1100" swimtime="00:13:47.71" />
                    <SPLIT distance="1150" swimtime="00:14:26.16" />
                    <SPLIT distance="1200" swimtime="00:15:05.39" />
                    <SPLIT distance="1250" swimtime="00:15:45.18" />
                    <SPLIT distance="1300" swimtime="00:16:25.44" />
                    <SPLIT distance="1350" swimtime="00:17:04.73" />
                    <SPLIT distance="1400" swimtime="00:17:44.06" />
                    <SPLIT distance="1450" swimtime="00:18:23.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="544" reactiontime="+97" swimtime="00:02:34.33" resultid="8931" heatid="14261" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="628" reactiontime="+87" swimtime="00:02:11.94" resultid="8932" heatid="14332" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:04.91" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="673" reactiontime="+84" swimtime="00:01:04.58" resultid="8933" heatid="14359" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="598" reactiontime="+85" swimtime="00:04:45.66" resultid="8934" heatid="14398" lane="5" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:44.04" />
                    <SPLIT distance="200" swimtime="00:02:20.70" />
                    <SPLIT distance="250" swimtime="00:02:57.10" />
                    <SPLIT distance="300" swimtime="00:03:33.93" />
                    <SPLIT distance="350" swimtime="00:04:10.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-15" firstname="Jessica" gender="F" lastname="Thorpe" nation="GBR" athleteid="8949">
              <RESULTS>
                <RESULT eventid="1090" points="638" reactiontime="+93" swimtime="00:02:46.10" resultid="8950" heatid="14165" lane="2" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:02:05.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="809" reactiontime="+74" swimtime="00:10:12.07" resultid="8951" heatid="14178" lane="5" entrytime="00:10:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.50" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                    <SPLIT distance="200" swimtime="00:02:27.42" />
                    <SPLIT distance="250" swimtime="00:03:06.06" />
                    <SPLIT distance="300" swimtime="00:03:44.63" />
                    <SPLIT distance="350" swimtime="00:04:23.25" />
                    <SPLIT distance="400" swimtime="00:05:02.27" />
                    <SPLIT distance="450" swimtime="00:05:40.76" />
                    <SPLIT distance="500" swimtime="00:06:19.51" />
                    <SPLIT distance="550" swimtime="00:06:58.56" />
                    <SPLIT distance="600" swimtime="00:07:37.42" />
                    <SPLIT distance="650" swimtime="00:08:16.32" />
                    <SPLIT distance="700" swimtime="00:08:55.13" />
                    <SPLIT distance="750" swimtime="00:09:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="563" reactiontime="+73" swimtime="00:03:04.99" resultid="8952" heatid="14211" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:01:26.48" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="540" reactiontime="+91" swimtime="00:01:19.60" resultid="8953" heatid="14243" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="8954" heatid="14342" lane="6" entrytime="00:05:35.00" />
                <RESULT eventid="8613" points="562" reactiontime="+78" swimtime="00:01:17.27" resultid="8955" heatid="14352" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="742" reactiontime="+79" swimtime="00:05:02.05" resultid="8956" heatid="14393" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                    <SPLIT distance="200" swimtime="00:02:28.68" />
                    <SPLIT distance="250" swimtime="00:03:07.39" />
                    <SPLIT distance="300" swimtime="00:03:45.88" />
                    <SPLIT distance="350" swimtime="00:04:24.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="10313" name="CSIR MOS Dąbrowa Górnicza">
          <CONTACT email="mariuszwaliczek@interia.pl" name="Waliczek" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1997-06-01" firstname="Dawid" gender="M" lastname="Nowodworski" nation="POL" license="102711700137" athleteid="10321">
              <RESULTS>
                <RESULT eventid="1075" points="938" reactiontime="+76" swimtime="00:00:23.43" resultid="10322" heatid="14161" lane="3" entrytime="00:00:23.00" />
                <RESULT eventid="8213" points="912" reactiontime="+92" swimtime="00:00:26.71" resultid="10323" heatid="14207" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="8309" points="951" reactiontime="+73" swimtime="00:00:57.17" resultid="10324" heatid="14255" lane="5" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="1011" reactiontime="+43" swimtime="00:00:24.67" resultid="10325" heatid="14302" lane="2" entrytime="00:00:25.00" />
                <RESULT eventid="8630" points="871" reactiontime="+78" swimtime="00:00:56.86" resultid="10326" heatid="14361" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="901" reactiontime="+70" swimtime="00:00:29.25" resultid="10327" heatid="14389" lane="2" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-22" firstname="Anna" gender="F" lastname="Teresko" nation="POL" license="102711100021" athleteid="10334">
              <RESULTS>
                <RESULT eventid="8196" points="766" reactiontime="+76" swimtime="00:00:31.99" resultid="10335" heatid="14197" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="8325" points="804" reactiontime="+80" swimtime="00:02:25.63" resultid="10336" heatid="14257" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="834" reactiontime="+87" swimtime="00:01:08.40" resultid="10337" heatid="14307" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="861" reactiontime="+88" swimtime="00:02:09.42" resultid="10338" heatid="14321" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="10339" heatid="14342" lane="5" entrytime="00:05:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="10314">
              <RESULTS>
                <RESULT eventid="8213" points="627" reactiontime="+73" swimtime="00:00:30.27" resultid="10315" heatid="14207" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="10316" heatid="14262" lane="0" entrytime="00:02:30.00" />
                <RESULT eventid="8454" points="788" reactiontime="+71" swimtime="00:00:26.80" resultid="10317" heatid="14301" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="8486" points="607" reactiontime="+87" swimtime="00:01:05.14" resultid="10318" heatid="14315" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="611" reactiontime="+76" swimtime="00:01:03.99" resultid="10319" heatid="14361" lane="0" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="583" reactiontime="+76" swimtime="00:02:29.76" resultid="10320" heatid="14371" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-21" firstname="Patryk" gender="M" lastname="Droś" nation="POL" license="102711200122" athleteid="10328">
              <RESULTS>
                <RESULT eventid="8245" points="758" reactiontime="+71" swimtime="00:02:30.31" resultid="10329" heatid="14217" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="10330" heatid="14237" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="8341" points="540" reactiontime="+72" swimtime="00:02:33.24" resultid="10331" heatid="14262" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="840" reactiontime="+71" swimtime="00:01:05.42" resultid="10332" heatid="14284" lane="6" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="787" reactiontime="+77" swimtime="00:01:59.17" resultid="10333" heatid="14333" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="100" swimtime="00:00:58.17" />
                    <SPLIT distance="150" swimtime="00:01:28.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10464" name="Delfin Masters Łódz">
          <CONTACT email="cewa@poczta.fm" name="Ewa Kadłubiec" phone="604627966" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-12" firstname="Maja" gender="F" lastname="Klusek" nation="POL" athleteid="10465">
              <RESULTS>
                <RESULT eventid="1090" points="513" reactiontime="+101" swimtime="00:03:03.30" resultid="10466" heatid="14164" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                    <SPLIT distance="150" swimtime="00:02:18.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="463" reactiontime="+99" swimtime="00:03:10.82" resultid="10467" heatid="14257" lane="9" entrytime="00:03:15.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                    <SPLIT distance="150" swimtime="00:02:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="558" reactiontime="+108" swimtime="00:00:36.28" resultid="10468" heatid="14288" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="8613" points="473" reactiontime="+107" swimtime="00:01:24.81" resultid="10469" heatid="14352" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12739" name="Dąbrowska Szkoła Pływania">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="12740">
              <RESULTS>
                <RESULT eventid="8213" points="324" reactiontime="+73" swimtime="00:00:36.45" resultid="12741" heatid="14200" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="8245" points="479" reactiontime="+72" swimtime="00:02:56.84" resultid="12742" heatid="14213" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:02:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="521" reactiontime="+78" swimtime="00:01:17.04" resultid="12743" heatid="14276" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="379" reactiontime="+73" swimtime="00:01:16.05" resultid="12744" heatid="14310" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="279" reactiontime="+69" swimtime="00:02:57.72" resultid="12745" heatid="14367" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="100" swimtime="00:01:28.81" />
                    <SPLIT distance="150" swimtime="00:02:15.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="492" reactiontime="+72" swimtime="00:00:35.78" resultid="12746" heatid="14380" lane="6" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-03-24" firstname="Kinga" gender="F" lastname="Pluta" nation="POL" athleteid="12747">
              <RESULTS>
                <RESULT eventid="8196" points="404" reactiontime="+83" swimtime="00:00:39.60" resultid="12748" heatid="14194" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="8229" points="509" reactiontime="+70" swimtime="00:03:10.14" resultid="12749" heatid="14209" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="150" swimtime="00:02:18.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="570" reactiontime="+81" swimtime="00:01:25.26" resultid="12750" heatid="14271" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="480" reactiontime="+83" swimtime="00:01:22.22" resultid="12751" heatid="14304" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="426" reactiontime="+82" swimtime="00:02:55.05" resultid="12752" heatid="14363" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                    <SPLIT distance="150" swimtime="00:02:10.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="580" reactiontime="+72" swimtime="00:00:39.37" resultid="12753" heatid="14374" lane="9" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="10563" name="Euro-Lviv MSC">
          <CONTACT email="mk.dmitry@gmail.com" name="Melnyk Dmytro" phone="+380965422460" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="10564">
              <RESULTS>
                <RESULT eventid="1075" points="798" reactiontime="+65" swimtime="00:00:25.61" resultid="10565" heatid="14158" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1150" points="533" reactiontime="+83" swimtime="00:10:30.72" resultid="10566" heatid="14183" lane="4" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:51.05" />
                    <SPLIT distance="200" swimtime="00:02:30.93" />
                    <SPLIT distance="250" swimtime="00:03:10.84" />
                    <SPLIT distance="300" swimtime="00:03:51.28" />
                    <SPLIT distance="350" swimtime="00:04:31.87" />
                    <SPLIT distance="400" swimtime="00:05:12.33" />
                    <SPLIT distance="450" swimtime="00:05:53.12" />
                    <SPLIT distance="500" swimtime="00:06:33.84" />
                    <SPLIT distance="550" swimtime="00:07:54.64" />
                    <SPLIT distance="600" swimtime="00:08:35.26" />
                    <SPLIT distance="650" swimtime="00:09:15.82" />
                    <SPLIT distance="700" swimtime="00:09:56.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="755" reactiontime="+74" swimtime="00:00:57.18" resultid="10567" heatid="14234" lane="4" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="732" reactiontime="+70" swimtime="00:01:12.80" resultid="10568" heatid="14283" lane="8" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="271" reactiontime="+64" swimtime="00:00:45.57" resultid="10569" heatid="14388" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="8742" points="506" reactiontime="+96" swimtime="00:05:01.89" resultid="10570" heatid="14400" lane="5" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                    <SPLIT distance="200" swimtime="00:02:29.30" />
                    <SPLIT distance="250" swimtime="00:03:08.09" />
                    <SPLIT distance="300" swimtime="00:03:46.80" />
                    <SPLIT distance="350" swimtime="00:04:25.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-02-27" firstname="Olena" gender="F" lastname="Pereyaslova" nation="UKR" athleteid="10585">
              <RESULTS>
                <RESULT eventid="1058" points="572" reactiontime="+100" swimtime="00:00:34.33" resultid="10586" heatid="14138" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="8261" points="511" reactiontime="+99" swimtime="00:01:17.48" resultid="10587" heatid="14220" lane="5" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="463" reactiontime="+82" swimtime="00:02:54.34" resultid="10588" heatid="14319" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="435" reactiontime="+86" swimtime="00:06:17.72" resultid="10589" heatid="14395" lane="8" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:28.73" />
                    <SPLIT distance="150" swimtime="00:02:18.19" />
                    <SPLIT distance="200" swimtime="00:03:08.00" />
                    <SPLIT distance="250" swimtime="00:03:56.77" />
                    <SPLIT distance="300" swimtime="00:04:45.39" />
                    <SPLIT distance="350" swimtime="00:05:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="10571">
              <RESULTS>
                <RESULT eventid="1075" points="751" reactiontime="+93" swimtime="00:00:26.26" resultid="10572" heatid="14158" lane="3" entrytime="00:00:25.95" />
                <RESULT eventid="8277" points="747" reactiontime="+87" swimtime="00:00:58.30" resultid="10573" heatid="14235" lane="1" entrytime="00:00:57.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="709" reactiontime="+80" swimtime="00:02:27.60" resultid="10574" heatid="14262" lane="8" entrytime="00:02:28.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="904" reactiontime="+71" swimtime="00:00:27.34" resultid="10575" heatid="14301" lane="9" entrytime="00:00:27.40" />
                <RESULT eventid="8630" points="778" reactiontime="+82" swimtime="00:01:03.93" resultid="10576" heatid="14359" lane="2" entrytime="00:01:04.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-18" firstname="Vladyslav" gender="M" lastname="Horovoy" nation="UKR" athleteid="10577">
              <RESULTS>
                <RESULT eventid="1105" points="964" reactiontime="+89" swimtime="00:02:16.94" resultid="10578" heatid="14174" lane="0" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:45.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="774" reactiontime="+75" swimtime="00:00:30.35" resultid="10579" heatid="14205" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="8309" points="904" reactiontime="+80" swimtime="00:01:02.11" resultid="10580" heatid="14254" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="900" reactiontime="+79" swimtime="00:01:08.40" resultid="10581" heatid="14283" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="834" reactiontime="+73" swimtime="00:02:01.84" resultid="10582" heatid="14333" lane="7" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:00:58.49" />
                    <SPLIT distance="150" swimtime="00:01:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K1 - Pływak wykonał kopnięcie delfinowe po pierwszym kopnięciu do stylu klasycznego (pierwszy ruch po starcie lub nawrocie)." eventid="8694" reactiontime="+69" status="DSQ" swimtime="00:00:30.99" resultid="10583" heatid="14388" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="8742" points="783" reactiontime="+73" swimtime="00:04:26.71" resultid="10584" heatid="14398" lane="2" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:05.68" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                    <SPLIT distance="200" swimtime="00:02:15.38" />
                    <SPLIT distance="250" swimtime="00:02:49.90" />
                    <SPLIT distance="300" swimtime="00:03:24.03" />
                    <SPLIT distance="350" swimtime="00:03:56.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10498" name="Gdynia Masters">
          <CONTACT name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="10527">
              <RESULTS>
                <RESULT eventid="1075" points="367" reactiontime="+115" swimtime="00:00:43.69" resultid="10528" heatid="14144" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1105" points="341" reactiontime="+121" swimtime="00:04:31.79" resultid="10529" heatid="14168" lane="0" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.87" />
                    <SPLIT distance="100" swimtime="00:03:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="381" reactiontime="+96" swimtime="00:00:52.25" resultid="10530" heatid="14200" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="8309" points="363" reactiontime="+120" swimtime="00:01:56.99" resultid="10531" heatid="14246" lane="1" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="376" reactiontime="+107" swimtime="00:02:00.13" resultid="10532" heatid="14277" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="267" reactiontime="+111" swimtime="00:02:09.43" resultid="10533" heatid="14310" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="483" reactiontime="+124" swimtime="00:00:49.95" resultid="10534" heatid="14381" lane="9" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="10517">
              <RESULTS>
                <RESULT eventid="8179" points="380" reactiontime="+123" swimtime="00:30:22.31" resultid="10518" heatid="14191" lane="0" entrytime="00:29:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:02:51.58" />
                    <SPLIT distance="150" swimtime="00:03:53.15" />
                    <SPLIT distance="200" swimtime="00:04:53.77" />
                    <SPLIT distance="250" swimtime="00:06:56.33" />
                    <SPLIT distance="300" swimtime="00:08:57.72" />
                    <SPLIT distance="350" swimtime="00:09:58.12" />
                    <SPLIT distance="400" swimtime="00:10:58.96" />
                    <SPLIT distance="450" swimtime="00:12:01.22" />
                    <SPLIT distance="500" swimtime="00:13:03.13" />
                    <SPLIT distance="550" swimtime="00:14:05.58" />
                    <SPLIT distance="600" swimtime="00:15:06.77" />
                    <SPLIT distance="650" swimtime="00:16:06.65" />
                    <SPLIT distance="700" swimtime="00:17:09.29" />
                    <SPLIT distance="750" swimtime="00:18:10.78" />
                    <SPLIT distance="800" swimtime="00:19:13.77" />
                    <SPLIT distance="850" swimtime="00:20:15.07" />
                    <SPLIT distance="900" swimtime="00:21:16.87" />
                    <SPLIT distance="950" swimtime="00:22:18.37" />
                    <SPLIT distance="1000" swimtime="00:23:20.59" />
                    <SPLIT distance="1050" swimtime="00:24:20.94" />
                    <SPLIT distance="1100" swimtime="00:26:26.01" />
                    <SPLIT distance="1150" swimtime="00:27:28.14" />
                    <SPLIT distance="1200" swimtime="00:28:27.38" />
                    <SPLIT distance="1250" swimtime="00:29:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="162" reactiontime="+104" swimtime="00:05:06.98" resultid="10519" heatid="14259" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.00" />
                    <SPLIT distance="100" swimtime="00:02:14.70" />
                    <SPLIT distance="150" swimtime="00:03:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="353" reactiontime="+111" swimtime="00:08:40.64" resultid="10520" heatid="14344" lane="6" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.63" />
                    <SPLIT distance="100" swimtime="00:02:27.32" />
                    <SPLIT distance="150" swimtime="00:03:35.64" />
                    <SPLIT distance="200" swimtime="00:04:40.93" />
                    <SPLIT distance="250" swimtime="00:05:44.21" />
                    <SPLIT distance="300" swimtime="00:06:47.65" />
                    <SPLIT distance="350" swimtime="00:07:48.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="10521" heatid="14354" lane="8" entrytime="00:02:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Grażyna" gender="F" lastname="Heisler" nation="POL" athleteid="10522">
              <RESULTS>
                <RESULT eventid="1058" points="432" reactiontime="+101" swimtime="00:00:42.63" resultid="10523" heatid="14135" lane="4" entrytime="00:00:47.00" />
                <RESULT eventid="8293" points="362" reactiontime="+106" swimtime="00:01:54.84" resultid="10524" heatid="14239" lane="8" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="370" reactiontime="+84" swimtime="00:02:01.88" resultid="10525" heatid="14304" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="360" reactiontime="+101" swimtime="00:00:57.95" resultid="10526" heatid="14373" lane="8" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="10499">
              <RESULTS>
                <RESULT eventid="1075" points="413" reactiontime="+101" swimtime="00:00:38.92" resultid="10500" heatid="14145" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="8213" points="164" reactiontime="+99" swimtime="00:01:03.27" resultid="10501" heatid="14200" lane="9" entrytime="00:00:58.00" />
                <RESULT eventid="8309" points="241" reactiontime="+109" swimtime="00:02:05.88" resultid="10502" heatid="14245" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="331" reactiontime="+98" swimtime="00:00:46.74" resultid="10503" heatid="14292" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="8694" points="163" reactiontime="+91" swimtime="00:01:04.92" resultid="10504" heatid="14380" lane="3" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Józef" gender="M" lastname="Stopiński" nation="POL" athleteid="10535">
              <RESULTS>
                <RESULT eventid="8454" points="793" reactiontime="+77" swimtime="00:00:26.88" resultid="10536" heatid="14300" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="8630" points="811" reactiontime="+66" swimtime="00:00:59.19" resultid="10537" heatid="14360" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="10505">
              <RESULTS>
                <RESULT eventid="8196" points="463" reactiontime="+94" swimtime="00:00:46.64" resultid="10506" heatid="14194" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="8261" points="389" reactiontime="+108" swimtime="00:01:27.80" resultid="10507" heatid="14219" lane="3" entrytime="00:01:28.00" />
                <RESULT eventid="8470" points="382" reactiontime="+82" swimtime="00:01:47.62" resultid="10508" heatid="14305" lane="3" entrytime="00:01:32.00" />
                <RESULT eventid="8502" points="317" reactiontime="+114" swimtime="00:03:22.91" resultid="10509" heatid="14318" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:35.80" />
                    <SPLIT distance="150" swimtime="00:02:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="420" reactiontime="+94" swimtime="00:03:39.58" resultid="10510" heatid="14364" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="334" reactiontime="+109" swimtime="00:07:04.79" resultid="10511" heatid="14395" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:35.55" />
                    <SPLIT distance="150" swimtime="00:02:30.18" />
                    <SPLIT distance="200" swimtime="00:03:25.35" />
                    <SPLIT distance="250" swimtime="00:04:20.69" />
                    <SPLIT distance="300" swimtime="00:05:16.32" />
                    <SPLIT distance="350" swimtime="00:06:12.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="10512">
              <RESULTS>
                <RESULT eventid="8245" points="715" reactiontime="+93" swimtime="00:03:23.69" resultid="10513" heatid="14214" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:35.20" />
                    <SPLIT distance="150" swimtime="00:02:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10514" heatid="14247" lane="9" entrytime="00:01:36.00" />
                <RESULT eventid="8406" points="700" reactiontime="+100" swimtime="00:01:29.43" resultid="10515" heatid="14278" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="10516" heatid="14292" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="8694" points="685" reactiontime="+93" swimtime="00:00:39.57" resultid="13227" heatid="14382" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+119" swimtime="00:02:46.94" resultid="10538" heatid="14336" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:11.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10527" number="1" reactiontime="+119" />
                    <RELAYPOSITION athleteid="10499" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10517" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="10512" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8373" reactiontime="+93" swimtime="00:03:02.36" resultid="10539" heatid="14265" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:34.86" />
                    <SPLIT distance="150" swimtime="00:02:20.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10527" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="10512" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="10499" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="10517" number="4" reactiontime="+80" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+85" swimtime="00:02:53.22" resultid="11415" heatid="14390" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                    <SPLIT distance="150" swimtime="00:02:11.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10505" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="10512" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="10499" number="3" reactiontime="+11" />
                    <RELAYPOSITION athleteid="10522" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10829" name="IKS Konstancin">
          <CONTACT email="RAFAL@JUCHNO.COM" name="JUCHNO" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="10830">
              <RESULTS>
                <RESULT eventid="1075" points="687" reactiontime="+74" swimtime="00:00:27.05" resultid="10831" heatid="14153" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1105" points="593" reactiontime="+80" swimtime="00:02:41.01" resultid="10832" heatid="14170" lane="3" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="701" reactiontime="+85" swimtime="00:00:59.57" resultid="10833" heatid="14233" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="562" reactiontime="+81" swimtime="00:01:12.77" resultid="10834" heatid="14249" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="622" reactiontime="+81" swimtime="00:00:30.97" resultid="10835" heatid="14296" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="8518" points="636" reactiontime="+66" swimtime="00:02:13.38" resultid="10836" heatid="14331" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:04.03" />
                    <SPLIT distance="150" swimtime="00:01:39.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-03" firstname="Rafal" gender="M" lastname="Juchno" nation="POL" license="103714700087" athleteid="11111">
              <RESULTS>
                <RESULT eventid="1075" points="583" reactiontime="+93" swimtime="00:00:28.43" resultid="11112" heatid="14150" lane="5" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="456" reactiontime="+86" swimtime="00:01:07.65" resultid="11113" heatid="14229" lane="8" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="422" reactiontime="+90" swimtime="00:01:27.42" resultid="11114" heatid="14279" lane="8" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="353" reactiontime="+95" swimtime="00:00:35.54" resultid="11115" heatid="14293" lane="4" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-02-23" firstname="Maciej" gender="M" lastname="Piłatowicz" nation="POL" athleteid="11103">
              <RESULTS>
                <RESULT eventid="8179" status="DNS" swimtime="00:00:00.00" resultid="11104" heatid="14192" lane="5" entrytime="00:23:00.00" entrycourse="SCM" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="11105" heatid="14229" lane="7" entrytime="00:01:08.00" entrycourse="SCM" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="11106" heatid="14248" lane="7" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="11107" heatid="14294" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="11108" heatid="14328" lane="1" entrytime="00:02:30.00" entrycourse="SCM" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="11109" heatid="14356" lane="7" entrytime="00:01:20.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="PDL" clubid="11116" name="ISWIM Białystok">
          <CONTACT city="Białystok" email="biuro@iswim.bialystok.pl" internet="www.iswim.bialystok.pl" name="Sebastian Humbla" phone="782997050" state="PDL" street="Wierzbowa 3" zip="15-743" />
          <ATHLETES>
            <ATHLETE birthdate="1979-02-13" firstname="Świderski" gender="M" lastname="Dawid" nation="POL" athleteid="11117">
              <RESULTS>
                <RESULT eventid="1075" points="596" reactiontime="+93" swimtime="00:00:27.32" resultid="11118" heatid="14155" lane="6" entrytime="00:00:27.20" entrycourse="SCM" />
                <RESULT eventid="8454" points="634" reactiontime="+88" swimtime="00:00:28.96" resultid="11119" heatid="14299" lane="4" entrytime="00:00:28.30" entrycourse="SCM" />
                <RESULT eventid="8630" points="581" reactiontime="+89" swimtime="00:01:06.14" resultid="11120" heatid="14360" lane="0" entrytime="00:01:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Agnieszka" gender="F" lastname="Stefanowska" nation="POL" athleteid="11143">
              <RESULTS>
                <RESULT eventid="1135" points="328" reactiontime="+90" swimtime="00:13:53.38" resultid="11144" heatid="14179" lane="3" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:17.99" />
                    <SPLIT distance="200" swimtime="00:03:08.74" />
                    <SPLIT distance="250" swimtime="00:04:00.50" />
                    <SPLIT distance="300" swimtime="00:04:53.72" />
                    <SPLIT distance="350" swimtime="00:05:47.07" />
                    <SPLIT distance="400" swimtime="00:06:42.01" />
                    <SPLIT distance="450" swimtime="00:07:36.89" />
                    <SPLIT distance="500" swimtime="00:08:31.43" />
                    <SPLIT distance="550" swimtime="00:09:25.27" />
                    <SPLIT distance="600" swimtime="00:10:19.85" />
                    <SPLIT distance="650" swimtime="00:11:15.30" />
                    <SPLIT distance="700" swimtime="00:12:09.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="261" reactiontime="+91" swimtime="00:03:51.00" resultid="11145" heatid="14256" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="357" reactiontime="+175" swimtime="00:03:02.17" resultid="11146" heatid="14319" lane="1" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:26.05" />
                    <SPLIT distance="150" swimtime="00:02:15.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-24" firstname="Sebastian" gender="M" lastname="Humbla" nation="POL" athleteid="11135">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1075" reactiontime="+71" status="DSQ" swimtime="00:00:26.76" resultid="11136" heatid="14157" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="8277" points="577" reactiontime="+105" swimtime="00:01:01.76" resultid="11137" heatid="14234" lane="3" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8454" reactiontime="+84" status="DSQ" swimtime="00:00:29.51" resultid="11138" heatid="14299" lane="2" entrytime="00:00:28.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-08-27" firstname="Józek" gender="M" lastname="Sawicki" nation="POL" athleteid="11139">
              <RESULTS>
                <RESULT eventid="1150" points="514" reactiontime="+89" swimtime="00:10:42.10" resultid="11140" heatid="14182" lane="2" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="200" swimtime="00:02:30.30" />
                    <SPLIT distance="250" swimtime="00:03:11.57" />
                    <SPLIT distance="300" swimtime="00:03:53.62" />
                    <SPLIT distance="350" swimtime="00:04:35.87" />
                    <SPLIT distance="400" swimtime="00:05:16.76" />
                    <SPLIT distance="450" swimtime="00:05:58.74" />
                    <SPLIT distance="500" swimtime="00:06:41.08" />
                    <SPLIT distance="550" swimtime="00:08:03.87" />
                    <SPLIT distance="600" swimtime="00:08:45.16" />
                    <SPLIT distance="650" swimtime="00:09:26.32" />
                    <SPLIT distance="700" swimtime="00:10:05.21" />
                    <SPLIT distance="750" swimtime="00:10:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="452" reactiontime="+76" swimtime="00:01:03.30" resultid="11141" heatid="14235" lane="7" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="11142" heatid="14332" lane="3" entrytime="00:02:06.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-12" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="11124">
              <RESULTS>
                <RESULT eventid="8213" points="614" reactiontime="+77" swimtime="00:00:32.78" resultid="11125" heatid="14204" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="11126" heatid="14281" lane="0" entrytime="00:01:22.00" />
                <RESULT eventid="8694" points="749" reactiontime="+84" swimtime="00:00:33.43" resultid="11127" heatid="14387" lane="7" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-09-21" firstname="Bartek" gender="M" lastname="Markowski" nation="POL" athleteid="11147">
              <RESULTS>
                <RESULT eventid="1150" points="269" reactiontime="+106" swimtime="00:13:11.76" resultid="11148" heatid="14184" lane="3" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:12.06" />
                    <SPLIT distance="200" swimtime="00:03:01.92" />
                    <SPLIT distance="250" swimtime="00:03:53.37" />
                    <SPLIT distance="300" swimtime="00:04:44.70" />
                    <SPLIT distance="350" swimtime="00:05:35.89" />
                    <SPLIT distance="400" swimtime="00:06:27.31" />
                    <SPLIT distance="450" swimtime="00:07:19.05" />
                    <SPLIT distance="500" swimtime="00:08:11.08" />
                    <SPLIT distance="550" swimtime="00:09:03.19" />
                    <SPLIT distance="600" swimtime="00:09:54.90" />
                    <SPLIT distance="650" swimtime="00:10:46.39" />
                    <SPLIT distance="700" swimtime="00:11:37.66" />
                    <SPLIT distance="750" swimtime="00:12:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="335" reactiontime="+91" swimtime="00:01:14.94" resultid="11149" heatid="14228" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="278" reactiontime="+96" swimtime="00:02:53.03" resultid="11150" heatid="14327" lane="8" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:05.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-20" firstname="Ewa" gender="F" lastname="Markowska" nation="POL" athleteid="11128">
              <RESULTS>
                <RESULT comment="przekroczony limit czasu" eventid="1165" reactiontime="+112" status="DSQ" swimtime="00:27:46.78" resultid="11129" heatid="14188" lane="6" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:02:30.38" />
                    <SPLIT distance="200" swimtime="00:03:24.30" />
                    <SPLIT distance="250" swimtime="00:04:19.29" />
                    <SPLIT distance="300" swimtime="00:05:15.70" />
                    <SPLIT distance="350" swimtime="00:06:11.42" />
                    <SPLIT distance="400" swimtime="00:07:07.89" />
                    <SPLIT distance="450" swimtime="00:08:03.99" />
                    <SPLIT distance="500" swimtime="00:09:00.44" />
                    <SPLIT distance="550" swimtime="00:09:56.72" />
                    <SPLIT distance="600" swimtime="00:10:51.06" />
                    <SPLIT distance="650" swimtime="00:11:46.63" />
                    <SPLIT distance="700" swimtime="00:12:43.84" />
                    <SPLIT distance="750" swimtime="00:13:40.66" />
                    <SPLIT distance="800" swimtime="00:14:37.30" />
                    <SPLIT distance="850" swimtime="00:15:34.45" />
                    <SPLIT distance="900" swimtime="00:16:31.18" />
                    <SPLIT distance="950" swimtime="00:17:28.69" />
                    <SPLIT distance="1000" swimtime="00:18:25.65" />
                    <SPLIT distance="1050" swimtime="00:19:23.68" />
                    <SPLIT distance="1100" swimtime="00:20:21.81" />
                    <SPLIT distance="1150" swimtime="00:21:18.59" />
                    <SPLIT distance="1200" swimtime="00:22:16.37" />
                    <SPLIT distance="1250" swimtime="00:23:15.43" />
                    <SPLIT distance="1300" swimtime="00:24:12.43" />
                    <SPLIT distance="1350" swimtime="00:25:10.00" />
                    <SPLIT distance="1400" swimtime="00:26:04.73" />
                    <SPLIT distance="1450" swimtime="00:27:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="131" swimtime="00:04:51.29" resultid="11130" heatid="14256" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                    <SPLIT distance="100" swimtime="00:02:08.29" />
                    <SPLIT distance="150" swimtime="00:03:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="273" swimtime="00:08:06.05" resultid="11131" heatid="14341" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:02:04.23" />
                    <SPLIT distance="150" swimtime="00:03:12.04" />
                    <SPLIT distance="200" swimtime="00:04:15.80" />
                    <SPLIT distance="250" swimtime="00:05:17.76" />
                    <SPLIT distance="300" swimtime="00:06:19.58" />
                    <SPLIT distance="350" swimtime="00:07:14.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-10" firstname="Dawid" gender="M" lastname="Perkowski" nation="POL" athleteid="11132">
              <RESULTS>
                <RESULT eventid="8341" points="590" reactiontime="+74" swimtime="00:02:28.78" resultid="11133" heatid="14262" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="786" reactiontime="+60" swimtime="00:00:26.82" resultid="11134" heatid="14301" lane="7" entrytime="00:00:26.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-16" firstname="Karol" gender="M" lastname="Traciecki" nation="POL" athleteid="11121">
              <RESULTS>
                <RESULT eventid="1105" points="406" reactiontime="+99" swimtime="00:02:52.62" resultid="11122" heatid="14172" lane="5" entrytime="00:02:30.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="483" reactiontime="+108" swimtime="00:03:02.02" resultid="11123" heatid="14216" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:24.48" />
                    <SPLIT distance="150" swimtime="00:02:13.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+78" swimtime="00:02:06.12" resultid="11151" heatid="14268" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:39.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11124" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="11121" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="11117" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="11135" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+87" swimtime="00:01:51.13" resultid="11153" heatid="14339" lane="0" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                    <SPLIT distance="100" swimtime="00:00:56.66" />
                    <SPLIT distance="150" swimtime="00:01:23.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11139" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="11124" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="11117" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="11135" number="4" reactiontime="+82" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11044" name="Jedynka Elbląg Masters">
          <CONTACT city="Elbląg" email="tomwysocki@onet.eu" name="Wysocki" phone="696427414" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1984-12-19" firstname="Krzysztof" gender="M" lastname="Kluge" nation="POL" athleteid="11074">
              <RESULTS>
                <RESULT eventid="1075" points="499" reactiontime="+79" swimtime="00:00:27.89" resultid="11075" heatid="14154" lane="5" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="11068">
              <RESULTS>
                <RESULT eventid="8630" points="901" reactiontime="+73" swimtime="00:01:04.46" resultid="11069" heatid="14358" lane="5" entrytime="00:01:06.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="814" reactiontime="+71" swimtime="00:04:38.94" resultid="11070" heatid="14399" lane="7" entrytime="00:04:43.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                    <SPLIT distance="150" swimtime="00:01:40.69" />
                    <SPLIT distance="200" swimtime="00:02:16.41" />
                    <SPLIT distance="250" swimtime="00:02:52.69" />
                    <SPLIT distance="300" swimtime="00:03:28.81" />
                    <SPLIT distance="350" swimtime="00:04:04.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="11047">
              <RESULTS>
                <RESULT eventid="1058" points="231" reactiontime="+107" swimtime="00:00:42.57" resultid="11048" heatid="14136" lane="0" entrytime="00:00:45.14" />
                <RESULT comment="przekroczony limit czasu" eventid="1135" reactiontime="+99" status="DSQ" swimtime="00:14:26.26" resultid="11049" heatid="14179" lane="6" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:31.39" />
                    <SPLIT distance="200" swimtime="00:03:26.31" />
                    <SPLIT distance="250" swimtime="00:04:22.31" />
                    <SPLIT distance="300" swimtime="00:05:17.91" />
                    <SPLIT distance="350" swimtime="00:06:13.48" />
                    <SPLIT distance="400" swimtime="00:07:09.06" />
                    <SPLIT distance="450" swimtime="00:08:04.21" />
                    <SPLIT distance="500" swimtime="00:08:59.53" />
                    <SPLIT distance="550" swimtime="00:09:54.88" />
                    <SPLIT distance="600" swimtime="00:10:49.81" />
                    <SPLIT distance="650" swimtime="00:11:44.31" />
                    <SPLIT distance="700" swimtime="00:12:39.27" />
                    <SPLIT distance="750" swimtime="00:13:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="236" reactiontime="+101" swimtime="00:01:32.97" resultid="11050" heatid="14219" lane="7" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="243" reactiontime="+124" swimtime="00:03:21.72" resultid="11051" heatid="14318" lane="1" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:36.69" />
                    <SPLIT distance="150" swimtime="00:02:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="264" reactiontime="+110" swimtime="00:07:06.07" resultid="11052" heatid="14396" lane="5" entrytime="00:07:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="100" swimtime="00:01:39.59" />
                    <SPLIT distance="150" swimtime="00:02:33.81" />
                    <SPLIT distance="200" swimtime="00:03:29.21" />
                    <SPLIT distance="250" swimtime="00:04:24.72" />
                    <SPLIT distance="300" swimtime="00:05:20.23" />
                    <SPLIT distance="350" swimtime="00:06:14.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-18" firstname="Tomasz" gender="M" lastname="Gleb" nation="POL" athleteid="11071">
              <RESULTS>
                <RESULT eventid="1075" points="536" reactiontime="+102" swimtime="00:00:31.27" resultid="11072" heatid="14150" lane="0" entrytime="00:00:30.25" />
                <RESULT eventid="8179" points="452" reactiontime="+114" swimtime="00:22:05.82" resultid="11073" heatid="14190" lane="0" entrytime="00:22:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:20.89" />
                    <SPLIT distance="150" swimtime="00:02:04.03" />
                    <SPLIT distance="200" swimtime="00:02:47.64" />
                    <SPLIT distance="250" swimtime="00:03:31.70" />
                    <SPLIT distance="300" swimtime="00:04:16.14" />
                    <SPLIT distance="350" swimtime="00:05:00.32" />
                    <SPLIT distance="400" swimtime="00:05:44.87" />
                    <SPLIT distance="450" swimtime="00:06:28.92" />
                    <SPLIT distance="500" swimtime="00:07:13.39" />
                    <SPLIT distance="550" swimtime="00:07:57.69" />
                    <SPLIT distance="600" swimtime="00:08:42.30" />
                    <SPLIT distance="650" swimtime="00:09:26.95" />
                    <SPLIT distance="700" swimtime="00:10:12.31" />
                    <SPLIT distance="750" swimtime="00:10:57.36" />
                    <SPLIT distance="800" swimtime="00:11:42.14" />
                    <SPLIT distance="850" swimtime="00:12:27.27" />
                    <SPLIT distance="900" swimtime="00:13:12.21" />
                    <SPLIT distance="950" swimtime="00:13:57.53" />
                    <SPLIT distance="1000" swimtime="00:14:42.43" />
                    <SPLIT distance="1050" swimtime="00:15:26.76" />
                    <SPLIT distance="1100" swimtime="00:16:10.84" />
                    <SPLIT distance="1150" swimtime="00:16:54.67" />
                    <SPLIT distance="1200" swimtime="00:17:39.15" />
                    <SPLIT distance="1250" swimtime="00:18:24.63" />
                    <SPLIT distance="1300" swimtime="00:19:09.65" />
                    <SPLIT distance="1350" swimtime="00:19:55.08" />
                    <SPLIT distance="1400" swimtime="00:20:39.86" />
                    <SPLIT distance="1450" swimtime="00:21:24.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="11053">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="11054" heatid="14163" lane="9" entrytime="00:04:12.00" />
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="11055" heatid="14180" lane="5" entrytime="00:14:45.00" />
                <RESULT eventid="8325" status="DNS" swimtime="00:00:00.00" resultid="11056" heatid="14256" lane="7" entrytime="00:04:25.00" />
                <RESULT eventid="8502" status="DNS" swimtime="00:00:00.00" resultid="11057" heatid="14318" lane="9" entrytime="00:03:35.00" />
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="11058" heatid="14340" lane="6" entrytime="00:08:55.00" />
                <RESULT eventid="8613" status="DNS" swimtime="00:00:00.00" resultid="11059" heatid="14350" lane="8" entrytime="00:02:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner Mateusiak" nation="POL" athleteid="11061">
              <RESULTS>
                <RESULT eventid="1135" status="DNF" swimtime="00:00:00.00" resultid="11062" heatid="14181" lane="4" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.03" />
                    <SPLIT distance="100" swimtime="00:02:32.21" />
                    <SPLIT distance="150" swimtime="00:03:52.49" />
                    <SPLIT distance="200" swimtime="00:05:13.40" />
                    <SPLIT distance="250" swimtime="00:06:33.62" />
                    <SPLIT distance="300" swimtime="00:07:52.38" />
                    <SPLIT distance="350" swimtime="00:09:12.09" />
                    <SPLIT distance="400" swimtime="00:10:31.70" />
                    <SPLIT distance="450" swimtime="00:11:51.06" />
                    <SPLIT distance="500" swimtime="00:13:10.56" />
                    <SPLIT distance="550" swimtime="00:14:30.24" />
                    <SPLIT distance="600" swimtime="00:15:49.21" />
                    <SPLIT distance="650" swimtime="00:17:08.32" />
                    <SPLIT distance="700" swimtime="00:18:24.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="108" swimtime="00:06:33.55" resultid="11063" heatid="14208" lane="7" entrytime="00:05:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.28" />
                    <SPLIT distance="100" swimtime="00:03:19.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="83" swimtime="00:03:16.83" resultid="11064" heatid="14269" lane="5" />
                <RESULT eventid="8470" points="152" reactiontime="+112" swimtime="00:02:36.99" resultid="11065" heatid="14304" lane="1" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="167" reactiontime="+75" swimtime="00:05:31.56" resultid="11066" heatid="14362" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.86" />
                    <SPLIT distance="100" swimtime="00:02:44.54" />
                    <SPLIT distance="150" swimtime="00:04:11.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="169" swimtime="00:10:32.78" resultid="11067" heatid="14396" lane="9" entrytime="00:10:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.70" />
                    <SPLIT distance="100" swimtime="00:02:30.05" />
                    <SPLIT distance="150" swimtime="00:03:52.98" />
                    <SPLIT distance="200" swimtime="00:05:14.26" />
                    <SPLIT distance="250" swimtime="00:06:34.26" />
                    <SPLIT distance="300" swimtime="00:07:53.11" />
                    <SPLIT distance="350" swimtime="00:09:11.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-21" firstname="Tomasz" gender="M" lastname="Wysocki" nation="POL" athleteid="11045">
              <RESULTS>
                <RESULT eventid="1075" points="747" reactiontime="+79" swimtime="00:00:25.34" resultid="11046" heatid="14158" lane="4" entrytime="00:00:25.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBS" clubid="8999" name="K.P. Stilon Gorzów Wlkp.">
          <CONTACT city="Gorzów Wlkp." email="kpstilon@hotmail.com" internet="http://www.kpstilon.gorzow.eu" name="K.Świderski" phone="512 428 265" state="LUBUS" street="UL. Słowiańska 1/ 42" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="9000">
              <RESULTS>
                <RESULT eventid="8179" points="370" reactiontime="+119" swimtime="00:27:16.63" resultid="9001" heatid="14191" lane="1" entrytime="00:27:12.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:38.88" />
                    <SPLIT distance="150" swimtime="00:02:33.03" />
                    <SPLIT distance="200" swimtime="00:03:27.79" />
                    <SPLIT distance="250" swimtime="00:04:23.07" />
                    <SPLIT distance="300" swimtime="00:05:17.76" />
                    <SPLIT distance="350" swimtime="00:06:13.04" />
                    <SPLIT distance="400" swimtime="00:07:07.65" />
                    <SPLIT distance="450" swimtime="00:08:03.03" />
                    <SPLIT distance="500" swimtime="00:08:58.81" />
                    <SPLIT distance="550" swimtime="00:09:54.29" />
                    <SPLIT distance="600" swimtime="00:10:50.14" />
                    <SPLIT distance="650" swimtime="00:11:45.80" />
                    <SPLIT distance="700" swimtime="00:12:41.26" />
                    <SPLIT distance="750" swimtime="00:13:36.15" />
                    <SPLIT distance="800" swimtime="00:14:31.25" />
                    <SPLIT distance="850" swimtime="00:15:26.24" />
                    <SPLIT distance="900" swimtime="00:16:20.98" />
                    <SPLIT distance="950" swimtime="00:17:16.47" />
                    <SPLIT distance="1000" swimtime="00:18:11.67" />
                    <SPLIT distance="1050" swimtime="00:19:06.81" />
                    <SPLIT distance="1100" swimtime="00:20:01.70" />
                    <SPLIT distance="1150" swimtime="00:20:57.70" />
                    <SPLIT distance="1200" swimtime="00:21:53.69" />
                    <SPLIT distance="1250" swimtime="00:22:48.82" />
                    <SPLIT distance="1300" swimtime="00:23:43.34" />
                    <SPLIT distance="1350" swimtime="00:24:37.66" />
                    <SPLIT distance="1400" swimtime="00:25:32.31" />
                    <SPLIT distance="1450" swimtime="00:26:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="266" reactiontime="+116" swimtime="00:01:33.06" resultid="9002" heatid="14225" lane="5" entrytime="00:01:28.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="9003" heatid="14310" lane="9" entrytime="00:02:05.00" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="9004" heatid="14324" lane="5" entrytime="00:03:17.35" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="11076" name="Kauno Takas">
          <CONTACT city="Kaunas" email="kaunotakas@gmail.com" name="Romaldas Bickauskas" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas Antanas" gender="M" lastname="Juodeska" nation="LTU" athleteid="11077">
              <RESULTS>
                <RESULT eventid="1075" points="643" reactiontime="+73" swimtime="00:00:30.21" resultid="11078" heatid="14151" lane="9" entrytime="00:00:29.99" />
                <RESULT eventid="8213" points="623" reactiontime="+86" swimtime="00:00:34.35" resultid="11079" heatid="14204" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="8309" points="637" reactiontime="+78" swimtime="00:01:16.42" resultid="11080" heatid="14249" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="568" reactiontime="+83" swimtime="00:01:18.19" resultid="11081" heatid="14312" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="563" reactiontime="+74" swimtime="00:00:36.93" resultid="11082" heatid="14385" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="10090" name="Kharkiv, Ukraine">
          <ATHLETES>
            <ATHLETE birthdate="1963-11-11" firstname="Mykhaylo" gender="M" lastname="Zakharchevskiy" nation="UKR" athleteid="10091">
              <RESULTS>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="10092" heatid="14345" lane="1" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PŁYWAK" nation="POL" region="WAR" clubid="10598" name="KPiRS PŁYWAK Płock">
          <CONTACT city="Płock" email="pawel.powichrowski@wp.pl" name="Powichrowski Paweł" phone="603694397" state="MAZ" street="Wiatraki 11 B" zip="09-402" />
          <ATHLETES>
            <ATHLETE birthdate="1998-05-02" firstname="Jakub" gender="M" lastname="Cichocki" nation="POL" athleteid="10606">
              <RESULTS>
                <RESULT eventid="8245" points="485" reactiontime="+86" swimtime="00:02:54.43" resultid="10607" heatid="14217" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="546" reactiontime="+72" swimtime="00:01:08.78" resultid="10608" heatid="14254" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="478" reactiontime="+83" swimtime="00:01:18.95" resultid="10609" heatid="14283" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="573" reactiontime="+78" swimtime="00:00:29.81" resultid="10610" heatid="14297" lane="6" entrytime="00:00:30.30" />
                <RESULT eventid="8694" points="440" reactiontime="+81" swimtime="00:00:37.15" resultid="10611" heatid="14387" lane="5" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-02-06" firstname="Dominik" gender="M" lastname="Bruchajzer" nation="POL" athleteid="10599">
              <RESULTS>
                <RESULT eventid="8277" points="611" reactiontime="+75" swimtime="00:00:59.69" resultid="10600" heatid="14235" lane="5" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="521" reactiontime="+80" swimtime="00:01:09.85" resultid="10601" heatid="14253" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="566" reactiontime="+77" swimtime="00:00:29.93" resultid="10602" heatid="14296" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="10603" heatid="14331" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="8694" points="444" reactiontime="+74" swimtime="00:00:37.02" resultid="10604" heatid="14387" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="8742" points="435" reactiontime="+157" swimtime="00:05:23.75" resultid="15633" heatid="14404" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:51.94" />
                    <SPLIT distance="200" swimtime="00:02:33.29" />
                    <SPLIT distance="250" swimtime="00:03:15.82" />
                    <SPLIT distance="300" swimtime="00:03:59.28" />
                    <SPLIT distance="350" swimtime="00:04:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-02" firstname="Katarzyna" gender="F" lastname="Janiszkiewicz" nation="POL" athleteid="10612">
              <RESULTS>
                <RESULT eventid="8229" points="424" reactiontime="+84" swimtime="00:03:22.12" resultid="10613" heatid="14209" lane="6" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:35.10" />
                    <SPLIT distance="150" swimtime="00:02:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="500" reactiontime="+85" swimtime="00:01:19.59" resultid="10614" heatid="14240" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="457" reactiontime="+92" swimtime="00:01:31.79" resultid="10615" heatid="14271" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="540" reactiontime="+92" swimtime="00:00:34.29" resultid="10616" heatid="14287" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="8678" points="528" reactiontime="+87" swimtime="00:00:40.62" resultid="10617" heatid="14375" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="KR" clubid="9669" name="Kraków Masters" shortname="Korona Kraków Masters">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz-Musiał" nation="POL" athleteid="9724">
              <RESULTS>
                <RESULT eventid="1165" points="273" swimtime="00:31:33.38" resultid="9725" heatid="14188" lane="7" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                    <SPLIT distance="100" swimtime="00:01:49.22" />
                    <SPLIT distance="150" swimtime="00:02:51.02" />
                    <SPLIT distance="200" swimtime="00:03:53.01" />
                    <SPLIT distance="250" swimtime="00:04:56.19" />
                    <SPLIT distance="300" swimtime="00:06:00.46" />
                    <SPLIT distance="350" swimtime="00:07:03.30" />
                    <SPLIT distance="400" swimtime="00:08:06.52" />
                    <SPLIT distance="450" swimtime="00:09:09.49" />
                    <SPLIT distance="500" swimtime="00:10:12.14" />
                    <SPLIT distance="550" swimtime="00:11:16.24" />
                    <SPLIT distance="600" swimtime="00:12:20.39" />
                    <SPLIT distance="650" swimtime="00:13:23.04" />
                    <SPLIT distance="700" swimtime="00:14:27.89" />
                    <SPLIT distance="750" swimtime="00:15:30.64" />
                    <SPLIT distance="800" swimtime="00:16:34.14" />
                    <SPLIT distance="850" swimtime="00:17:37.75" />
                    <SPLIT distance="900" swimtime="00:18:41.17" />
                    <SPLIT distance="950" swimtime="00:19:47.43" />
                    <SPLIT distance="1000" swimtime="00:20:50.73" />
                    <SPLIT distance="1050" swimtime="00:21:55.37" />
                    <SPLIT distance="1100" swimtime="00:22:58.85" />
                    <SPLIT distance="1150" swimtime="00:24:02.54" />
                    <SPLIT distance="1200" swimtime="00:25:07.08" />
                    <SPLIT distance="1250" swimtime="00:26:11.65" />
                    <SPLIT distance="1300" swimtime="00:27:15.81" />
                    <SPLIT distance="1350" swimtime="00:28:21.14" />
                    <SPLIT distance="1400" swimtime="00:29:24.74" />
                    <SPLIT distance="1450" swimtime="00:30:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="197" reactiontime="+120" swimtime="00:05:18.15" resultid="9726" heatid="14208" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.33" />
                    <SPLIT distance="100" swimtime="00:02:32.29" />
                    <SPLIT distance="150" swimtime="00:03:53.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="190" reactiontime="+93" swimtime="00:05:07.97" resultid="9727" heatid="14256" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.57" />
                    <SPLIT distance="100" swimtime="00:02:25.47" />
                    <SPLIT distance="150" swimtime="00:03:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="187" reactiontime="+101" swimtime="00:02:26.34" resultid="9728" heatid="14269" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="239" reactiontime="+102" swimtime="00:09:55.47" resultid="9729" heatid="14340" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.84" />
                    <SPLIT distance="100" swimtime="00:02:20.38" />
                    <SPLIT distance="150" swimtime="00:03:39.71" />
                    <SPLIT distance="200" swimtime="00:04:56.81" />
                    <SPLIT distance="250" swimtime="00:06:22.66" />
                    <SPLIT distance="300" swimtime="00:07:48.32" />
                    <SPLIT distance="350" swimtime="00:08:52.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="176" reactiontime="+56" swimtime="00:04:53.05" resultid="9730" heatid="14362" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.61" />
                    <SPLIT distance="100" swimtime="00:02:21.14" />
                    <SPLIT distance="150" swimtime="00:03:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="193" reactiontime="+103" swimtime="00:08:29.67" resultid="9731" heatid="14396" lane="2" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.63" />
                    <SPLIT distance="100" swimtime="00:01:56.16" />
                    <SPLIT distance="150" swimtime="00:03:01.88" />
                    <SPLIT distance="200" swimtime="00:04:07.33" />
                    <SPLIT distance="250" swimtime="00:05:13.00" />
                    <SPLIT distance="300" swimtime="00:06:19.03" />
                    <SPLIT distance="350" swimtime="00:07:23.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-07-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="9750">
              <RESULTS>
                <RESULT eventid="1075" points="721" reactiontime="+71" swimtime="00:00:25.65" resultid="9751" heatid="14158" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="8277" points="670" reactiontime="+82" swimtime="00:00:58.77" resultid="9752" heatid="14224" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="569" reactiontime="+75" swimtime="00:01:08.52" resultid="9753" heatid="14253" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="454" reactiontime="+86" swimtime="00:01:13.41" resultid="9754" heatid="14308" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="9744">
              <RESULTS>
                <RESULT eventid="1075" points="322" reactiontime="+105" swimtime="00:00:45.62" resultid="9745" heatid="14144" lane="0" entrytime="00:00:45.50" />
                <RESULT eventid="8179" points="381" reactiontime="+115" swimtime="00:32:52.22" resultid="9746" heatid="14190" lane="9" entrytime="00:42:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.89" />
                    <SPLIT distance="100" swimtime="00:02:04.57" />
                    <SPLIT distance="150" swimtime="00:03:11.39" />
                    <SPLIT distance="200" swimtime="00:04:18.03" />
                    <SPLIT distance="250" swimtime="00:05:27.12" />
                    <SPLIT distance="300" swimtime="00:06:33.26" />
                    <SPLIT distance="350" swimtime="00:07:39.73" />
                    <SPLIT distance="400" swimtime="00:08:46.33" />
                    <SPLIT distance="450" swimtime="00:09:52.15" />
                    <SPLIT distance="500" swimtime="00:10:58.70" />
                    <SPLIT distance="550" swimtime="00:12:05.00" />
                    <SPLIT distance="600" swimtime="00:13:11.51" />
                    <SPLIT distance="650" swimtime="00:14:17.52" />
                    <SPLIT distance="700" swimtime="00:15:23.69" />
                    <SPLIT distance="750" swimtime="00:16:29.98" />
                    <SPLIT distance="800" swimtime="00:17:36.30" />
                    <SPLIT distance="850" swimtime="00:18:40.79" />
                    <SPLIT distance="900" swimtime="00:19:46.27" />
                    <SPLIT distance="950" swimtime="00:20:52.62" />
                    <SPLIT distance="1000" swimtime="00:21:58.49" />
                    <SPLIT distance="1050" swimtime="00:23:04.63" />
                    <SPLIT distance="1100" swimtime="00:24:11.19" />
                    <SPLIT distance="1150" swimtime="00:25:17.35" />
                    <SPLIT distance="1200" swimtime="00:26:23.53" />
                    <SPLIT distance="1250" swimtime="00:27:29.58" />
                    <SPLIT distance="1300" swimtime="00:28:35.56" />
                    <SPLIT distance="1350" swimtime="00:29:41.14" />
                    <SPLIT distance="1400" swimtime="00:30:46.97" />
                    <SPLIT distance="1450" swimtime="00:31:52.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="334" reactiontime="+116" swimtime="00:01:42.48" resultid="9747" heatid="14225" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="298" reactiontime="+124" swimtime="00:03:57.94" resultid="9748" heatid="14324" lane="8" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:52.13" />
                    <SPLIT distance="150" swimtime="00:02:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="181" reactiontime="+119" swimtime="00:01:09.24" resultid="9749" heatid="14380" lane="7" entrytime="00:01:02.00" />
                <RESULT eventid="8742" points="299" reactiontime="+169" swimtime="00:08:47.89" resultid="15591" heatid="14404" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.65" />
                    <SPLIT distance="100" swimtime="00:02:07.77" />
                    <SPLIT distance="150" swimtime="00:03:16.33" />
                    <SPLIT distance="200" swimtime="00:04:24.85" />
                    <SPLIT distance="250" swimtime="00:05:33.16" />
                    <SPLIT distance="300" swimtime="00:06:40.52" />
                    <SPLIT distance="350" swimtime="00:07:47.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="9767">
              <RESULTS>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="9768" heatid="14187" lane="4" entrytime="00:16:15.00" />
                <RESULT eventid="8293" points="244" reactiontime="+128" swimtime="00:01:49.03" resultid="9769" heatid="14239" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="184" reactiontime="+123" swimtime="00:00:52.43" resultid="9770" heatid="14285" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="8502" points="138" reactiontime="+146" swimtime="00:04:09.65" resultid="9771" heatid="14317" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.14" />
                    <SPLIT distance="100" swimtime="00:01:45.79" />
                    <SPLIT distance="150" swimtime="00:02:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="165" reactiontime="+106" swimtime="00:02:00.33" resultid="9772" heatid="14350" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-24" firstname="Grzegorz" gender="M" lastname="Mucha" nation="POL" athleteid="9755">
              <RESULTS>
                <RESULT eventid="8406" points="556" reactiontime="+93" swimtime="00:01:24.56" resultid="9756" heatid="14280" lane="7" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="590" reactiontime="+87" swimtime="00:00:36.67" resultid="9757" heatid="14386" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="9706">
              <RESULTS>
                <RESULT eventid="1105" points="467" reactiontime="+126" swimtime="00:03:48.97" resultid="9707" heatid="14168" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:48.89" />
                    <SPLIT distance="150" swimtime="00:02:55.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="487" reactiontime="+144" swimtime="00:14:33.94" resultid="9708" heatid="14186" lane="4" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.89" />
                    <SPLIT distance="100" swimtime="00:01:48.28" />
                    <SPLIT distance="150" swimtime="00:02:44.31" />
                    <SPLIT distance="200" swimtime="00:03:40.53" />
                    <SPLIT distance="250" swimtime="00:04:36.27" />
                    <SPLIT distance="300" swimtime="00:05:31.25" />
                    <SPLIT distance="350" swimtime="00:06:26.50" />
                    <SPLIT distance="400" swimtime="00:07:22.38" />
                    <SPLIT distance="450" swimtime="00:08:17.53" />
                    <SPLIT distance="500" swimtime="00:09:12.96" />
                    <SPLIT distance="550" swimtime="00:10:08.48" />
                    <SPLIT distance="600" swimtime="00:11:03.44" />
                    <SPLIT distance="650" swimtime="00:11:58.00" />
                    <SPLIT distance="700" swimtime="00:12:53.79" />
                    <SPLIT distance="750" swimtime="00:13:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="683" reactiontime="+127" swimtime="00:01:17.01" resultid="9709" heatid="14227" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" reactiontime="+155" status="DNF" swimtime="00:00:00.00" resultid="9710" heatid="14259" lane="0" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.54" />
                    <SPLIT distance="100" swimtime="00:02:05.28" />
                    <SPLIT distance="150" swimtime="00:03:22.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="570" reactiontime="+128" swimtime="00:03:01.56" resultid="9711" heatid="14325" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="150" swimtime="00:02:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="441" reactiontime="+158" swimtime="00:08:40.31" resultid="9712" heatid="14344" lane="3" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.43" />
                    <SPLIT distance="100" swimtime="00:02:08.80" />
                    <SPLIT distance="150" swimtime="00:03:20.81" />
                    <SPLIT distance="200" swimtime="00:05:43.48" />
                    <SPLIT distance="250" swimtime="00:06:54.72" />
                    <SPLIT distance="300" swimtime="00:07:50.07" />
                    <SPLIT distance="350" swimtime="00:08:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="371" reactiontime="+126" swimtime="00:01:52.47" resultid="9713" heatid="14355" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="537" reactiontime="+131" swimtime="00:06:51.69" resultid="9714" heatid="14403" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:40.26" />
                    <SPLIT distance="150" swimtime="00:02:33.53" />
                    <SPLIT distance="200" swimtime="00:03:25.90" />
                    <SPLIT distance="250" swimtime="00:04:19.18" />
                    <SPLIT distance="300" swimtime="00:05:13.25" />
                    <SPLIT distance="350" swimtime="00:06:06.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="9758">
              <RESULTS>
                <RESULT eventid="1058" points="617" reactiontime="+106" swimtime="00:00:36.41" resultid="9759" heatid="14137" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1135" points="599" reactiontime="+124" swimtime="00:14:16.15" resultid="9760" heatid="14180" lane="3" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:34.77" />
                    <SPLIT distance="150" swimtime="00:02:28.44" />
                    <SPLIT distance="200" swimtime="00:03:21.45" />
                    <SPLIT distance="250" swimtime="00:04:16.01" />
                    <SPLIT distance="300" swimtime="00:05:10.16" />
                    <SPLIT distance="350" swimtime="00:06:05.70" />
                    <SPLIT distance="400" swimtime="00:07:01.13" />
                    <SPLIT distance="450" swimtime="00:07:55.67" />
                    <SPLIT distance="500" swimtime="00:08:50.34" />
                    <SPLIT distance="550" swimtime="00:10:40.20" />
                    <SPLIT distance="600" swimtime="00:11:35.27" />
                    <SPLIT distance="650" swimtime="00:12:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="680" reactiontime="+93" swimtime="00:00:43.77" resultid="9761" heatid="14194" lane="3" entrytime="00:00:47.00" />
                <RESULT eventid="8325" points="650" reactiontime="+126" swimtime="00:03:54.54" resultid="9762" heatid="14256" lane="6" entrytime="00:04:04.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:49.65" />
                    <SPLIT distance="150" swimtime="00:02:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="504" reactiontime="+108" swimtime="00:00:41.99" resultid="9763" heatid="14286" lane="7" entrytime="00:00:46.19" />
                <RESULT eventid="8566" points="548" reactiontime="+113" swimtime="00:07:45.96" resultid="9764" heatid="14340" lane="5" entrytime="00:08:14.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                    <SPLIT distance="100" swimtime="00:01:53.88" />
                    <SPLIT distance="150" swimtime="00:02:53.82" />
                    <SPLIT distance="200" swimtime="00:03:53.74" />
                    <SPLIT distance="250" swimtime="00:04:58.40" />
                    <SPLIT distance="300" swimtime="00:06:01.88" />
                    <SPLIT distance="350" swimtime="00:06:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="459" reactiontime="+109" swimtime="00:01:45.57" resultid="9765" heatid="14350" lane="6" entrytime="00:01:46.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="524" swimtime="00:03:46.86" resultid="9766" heatid="14363" lane="6" entrytime="00:03:45.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                    <SPLIT distance="100" swimtime="00:01:49.90" />
                    <SPLIT distance="150" swimtime="00:02:51.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="9689">
              <RESULTS>
                <RESULT eventid="1075" points="143" reactiontime="+115" swimtime="00:00:51.31" resultid="9690" heatid="14143" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="8213" points="110" reactiontime="+96" swimtime="00:01:06.32" resultid="9691" heatid="14199" lane="6" entrytime="00:01:04.00" />
                <RESULT eventid="8277" points="138" reactiontime="+124" swimtime="00:01:55.79" resultid="9692" heatid="14225" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="122" reactiontime="+119" swimtime="00:02:28.82" resultid="9693" heatid="14276" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="128" reactiontime="+105" swimtime="00:04:30.33" resultid="9694" heatid="14323" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                    <SPLIT distance="100" swimtime="00:02:04.92" />
                    <SPLIT distance="150" swimtime="00:03:18.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="121" reactiontime="+109" swimtime="00:05:20.57" resultid="9695" heatid="14367" lane="9" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.65" />
                    <SPLIT distance="100" swimtime="00:02:34.33" />
                    <SPLIT distance="150" swimtime="00:03:57.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="125" reactiontime="+120" swimtime="00:01:05.42" resultid="9696" heatid="14380" lane="8" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="9732">
              <RESULTS>
                <RESULT eventid="8213" points="141" reactiontime="+147" swimtime="00:01:06.54" resultid="9733" heatid="14200" lane="0" entrytime="00:00:58.00" />
                <RESULT eventid="8486" points="191" reactiontime="+152" swimtime="00:02:10.37" resultid="9734" heatid="14309" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="256" reactiontime="+97" swimtime="00:04:46.24" resultid="9735" heatid="14367" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.43" />
                    <SPLIT distance="100" swimtime="00:02:16.96" />
                    <SPLIT distance="150" swimtime="00:03:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="9670">
              <RESULTS>
                <RESULT eventid="1058" points="845" reactiontime="+73" swimtime="00:00:30.14" resultid="9671" heatid="14141" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="8196" points="822" reactiontime="+66" swimtime="00:00:35.45" resultid="9672" heatid="14196" lane="4" entrytime="00:00:36.50" />
                <RESULT eventid="8293" points="836" reactiontime="+82" swimtime="00:01:16.03" resultid="9673" heatid="14242" lane="3" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="861" reactiontime="+80" swimtime="00:00:32.74" resultid="9674" heatid="14288" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="8470" points="710" reactiontime="+81" swimtime="00:01:20.93" resultid="9675" heatid="14307" lane="9" entrytime="00:01:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="937" reactiontime="+77" swimtime="00:00:37.28" resultid="9676" heatid="14378" lane="9" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="9677">
              <RESULTS>
                <RESULT eventid="1058" points="808" reactiontime="+72" swimtime="00:00:29.33" resultid="9678" heatid="14141" lane="7" entrytime="00:00:29.20" />
                <RESULT eventid="8261" points="672" reactiontime="+92" swimtime="00:01:08.07" resultid="9679" heatid="14223" lane="0" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="811" reactiontime="+79" swimtime="00:00:32.18" resultid="9680" heatid="14289" lane="8" entrytime="00:00:32.40" />
                <RESULT eventid="8502" status="DNS" swimtime="00:00:00.00" resultid="9681" heatid="14321" lane="9" entrytime="00:02:32.00" />
                <RESULT eventid="8613" points="634" reactiontime="+84" swimtime="00:01:16.88" resultid="9682" heatid="14352" lane="8" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-10-20" firstname="Janusz" gender="M" lastname="Toporski" nation="POL" athleteid="9736">
              <RESULTS>
                <RESULT eventid="1105" points="307" reactiontime="+101" swimtime="00:03:35.56" resultid="9737" heatid="14168" lane="2" entrytime="00:03:41.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                    <SPLIT distance="150" swimtime="00:02:48.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="451" reactiontime="+89" swimtime="00:03:31.25" resultid="9738" heatid="14213" lane="6" entrytime="00:03:30.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.31" />
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="150" swimtime="00:02:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="280" reactiontime="+99" swimtime="00:01:40.49" resultid="9739" heatid="14246" lane="3" entrytime="00:01:39.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="301" reactiontime="+91" swimtime="00:01:41.65" resultid="9740" heatid="14277" lane="5" entrytime="00:01:41.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="311" reactiontime="+94" swimtime="00:07:56.08" resultid="9741" heatid="14344" lane="4" entrytime="00:08:05.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.36" />
                    <SPLIT distance="100" swimtime="00:01:53.78" />
                    <SPLIT distance="150" swimtime="00:03:00.01" />
                    <SPLIT distance="200" swimtime="00:04:10.88" />
                    <SPLIT distance="250" swimtime="00:05:12.16" />
                    <SPLIT distance="300" swimtime="00:06:10.20" />
                    <SPLIT distance="350" swimtime="00:07:06.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="221" reactiontime="+100" swimtime="00:01:47.03" resultid="9742" heatid="14355" lane="0" entrytime="00:01:42.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="278" reactiontime="+94" swimtime="00:00:46.70" resultid="9743" heatid="14381" lane="1" entrytime="00:00:47.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="9697">
              <RESULTS>
                <RESULT eventid="1058" points="677" reactiontime="+91" swimtime="00:00:33.68" resultid="9698" heatid="14138" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1135" points="561" reactiontime="+105" swimtime="00:12:18.41" resultid="9699" heatid="14179" lane="4" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                    <SPLIT distance="200" swimtime="00:02:57.47" />
                    <SPLIT distance="250" swimtime="00:03:44.59" />
                    <SPLIT distance="300" swimtime="00:04:32.63" />
                    <SPLIT distance="350" swimtime="00:05:20.22" />
                    <SPLIT distance="400" swimtime="00:06:06.95" />
                    <SPLIT distance="450" swimtime="00:06:53.69" />
                    <SPLIT distance="500" swimtime="00:07:40.27" />
                    <SPLIT distance="550" swimtime="00:08:27.38" />
                    <SPLIT distance="600" swimtime="00:09:14.26" />
                    <SPLIT distance="650" swimtime="00:10:01.14" />
                    <SPLIT distance="700" swimtime="00:10:48.18" />
                    <SPLIT distance="750" swimtime="00:11:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="613" reactiontime="+102" swimtime="00:01:15.49" resultid="9700" heatid="14221" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="687" reactiontime="+108" swimtime="00:03:20.84" resultid="9701" heatid="14256" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:32.90" />
                    <SPLIT distance="150" swimtime="00:02:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="638" reactiontime="+99" swimtime="00:00:38.02" resultid="9702" heatid="14287" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="8502" points="570" reactiontime="+100" swimtime="00:02:46.87" resultid="9703" heatid="14320" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="722" reactiontime="+90" swimtime="00:01:27.68" resultid="9704" heatid="14351" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="605" reactiontime="+102" swimtime="00:05:48.70" resultid="9705" heatid="14394" lane="8" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:21.65" />
                    <SPLIT distance="150" swimtime="00:02:06.10" />
                    <SPLIT distance="200" swimtime="00:02:51.38" />
                    <SPLIT distance="250" swimtime="00:03:37.06" />
                    <SPLIT distance="300" swimtime="00:04:22.10" />
                    <SPLIT distance="350" swimtime="00:05:07.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="9683">
              <RESULTS>
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="9684" heatid="14220" lane="7" entrytime="00:01:19.00" />
                <RESULT eventid="8438" points="514" reactiontime="+93" swimtime="00:00:37.46" resultid="9685" heatid="14287" lane="5" entrytime="00:00:37.90" />
                <RESULT eventid="8566" points="400" reactiontime="+108" swimtime="00:07:18.63" resultid="9686" heatid="14341" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:43.93" />
                    <SPLIT distance="150" swimtime="00:02:44.51" />
                    <SPLIT distance="200" swimtime="00:03:43.63" />
                    <SPLIT distance="250" swimtime="00:04:46.41" />
                    <SPLIT distance="300" swimtime="00:05:47.11" />
                    <SPLIT distance="350" swimtime="00:06:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="350" reactiontime="+81" swimtime="00:01:33.70" resultid="9687" heatid="14350" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="9688" heatid="14364" lane="1" entrytime="00:03:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="9715">
              <RESULTS>
                <RESULT eventid="1058" points="113" reactiontime="+108" swimtime="00:01:08.84" resultid="9716" heatid="14135" lane="0" entrytime="00:01:02.00" />
                <RESULT eventid="1090" points="87" reactiontime="+123" swimtime="00:07:10.34" resultid="9717" heatid="14162" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:53.74" />
                    <SPLIT distance="100" swimtime="00:04:02.95" />
                    <SPLIT distance="150" swimtime="00:05:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="137" reactiontime="+125" swimtime="00:02:24.63" resultid="9718" heatid="14218" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="89" reactiontime="+113" swimtime="00:03:06.23" resultid="9719" heatid="14239" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="159" reactiontime="+120" swimtime="00:02:59.03" resultid="9720" heatid="14270" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="45" reactiontime="+155" swimtime="00:01:42.58" resultid="9721" heatid="14285" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="8678" points="206" reactiontime="+108" swimtime="00:01:13.10" resultid="9722" heatid="14373" lane="9" entrytime="00:01:08.00" />
                <RESULT eventid="8726" points="145" reactiontime="+124" swimtime="00:12:02.41" resultid="9723" heatid="14396" lane="0" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.46" />
                    <SPLIT distance="100" swimtime="00:02:42.65" />
                    <SPLIT distance="150" swimtime="00:04:13.45" />
                    <SPLIT distance="200" swimtime="00:05:42.14" />
                    <SPLIT distance="250" swimtime="00:07:18.08" />
                    <SPLIT distance="300" swimtime="00:08:53.25" />
                    <SPLIT distance="350" swimtime="00:10:25.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków" number="1">
              <RESULTS>
                <RESULT eventid="8550" swimtime="00:02:29.91" resultid="9779" heatid="14337" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9744" number="1" />
                    <RELAYPOSITION athleteid="9755" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="9736" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="9706" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8373" reactiontime="+106" swimtime="00:02:56.46" resultid="9780" heatid="14265" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                    <SPLIT distance="100" swimtime="00:01:26.33" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9706" number="1" reactiontime="+106" />
                    <RELAYPOSITION athleteid="9755" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="9736" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="9744" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków" number="1">
              <RESULTS>
                <RESULT eventid="8534" reactiontime="+82" swimtime="00:02:07.09" resultid="9777" heatid="14335" lane="6" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:04.56" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9670" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="9683" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="9697" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="9677" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8357" reactiontime="+86" swimtime="00:02:24.38" resultid="9778" heatid="14264" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                    <SPLIT distance="150" swimtime="00:01:55.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9697" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="9670" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="9683" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9677" number="4" reactiontime="+1" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+87" swimtime="00:01:56.26" resultid="9773" heatid="14177" lane="2" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:01.75" />
                    <SPLIT distance="150" swimtime="00:01:30.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9670" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="9755" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="9677" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="9750" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+60" swimtime="00:02:20.15" resultid="9774" heatid="14391" lane="2" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:46.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9670" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="9755" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="9677" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="9706" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+115" swimtime="00:02:23.56" resultid="9775" heatid="14175" lane="3" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9697" number="1" reactiontime="+115" />
                    <RELAYPOSITION athleteid="9758" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="9706" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="9736" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+83" swimtime="00:02:52.66" resultid="9776" heatid="14390" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:01:52.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9758" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="9736" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9683" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="9744" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="8790" name="KS Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANWOL@POCZTA.ONET.PL" name="WOLNIEWICZ JANUSZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="8791">
              <RESULTS>
                <RESULT eventid="1075" points="459" reactiontime="+94" swimtime="00:00:37.57" resultid="8792" heatid="14146" lane="0" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="8179" points="447" reactiontime="+113" swimtime="00:30:11.64" resultid="8793" heatid="14191" lane="9" entrytime="00:30:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:44.90" />
                    <SPLIT distance="150" swimtime="00:02:42.60" />
                    <SPLIT distance="200" swimtime="00:03:41.86" />
                    <SPLIT distance="250" swimtime="00:04:41.92" />
                    <SPLIT distance="300" swimtime="00:05:42.59" />
                    <SPLIT distance="350" swimtime="00:06:43.22" />
                    <SPLIT distance="400" swimtime="00:07:43.48" />
                    <SPLIT distance="450" swimtime="00:08:44.19" />
                    <SPLIT distance="500" swimtime="00:09:45.11" />
                    <SPLIT distance="550" swimtime="00:10:44.46" />
                    <SPLIT distance="600" swimtime="00:11:44.82" />
                    <SPLIT distance="650" swimtime="00:12:44.57" />
                    <SPLIT distance="700" swimtime="00:13:45.07" />
                    <SPLIT distance="750" swimtime="00:14:45.25" />
                    <SPLIT distance="800" swimtime="00:15:46.97" />
                    <SPLIT distance="850" swimtime="00:16:49.02" />
                    <SPLIT distance="900" swimtime="00:17:50.15" />
                    <SPLIT distance="950" swimtime="00:18:52.68" />
                    <SPLIT distance="1000" swimtime="00:19:54.65" />
                    <SPLIT distance="1050" swimtime="00:20:57.40" />
                    <SPLIT distance="1100" swimtime="00:21:59.10" />
                    <SPLIT distance="1150" swimtime="00:23:02.49" />
                    <SPLIT distance="1200" swimtime="00:24:05.38" />
                    <SPLIT distance="1250" swimtime="00:25:05.20" />
                    <SPLIT distance="1300" swimtime="00:26:07.13" />
                    <SPLIT distance="1350" swimtime="00:27:09.38" />
                    <SPLIT distance="1400" swimtime="00:28:12.31" />
                    <SPLIT distance="1450" swimtime="00:29:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="496" reactiontime="+96" swimtime="00:01:25.67" resultid="8794" heatid="14226" lane="1" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="404" reactiontime="+100" swimtime="00:03:23.58" resultid="8795" heatid="14324" lane="6" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:34.31" />
                    <SPLIT distance="150" swimtime="00:02:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="403" reactiontime="+97" swimtime="00:07:33.13" resultid="8796" heatid="14403" lane="7" entrytime="00:07:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.55" />
                    <SPLIT distance="100" swimtime="00:01:42.15" />
                    <SPLIT distance="150" swimtime="00:02:39.96" />
                    <SPLIT distance="200" swimtime="00:03:37.89" />
                    <SPLIT distance="250" swimtime="00:04:36.87" />
                    <SPLIT distance="300" swimtime="00:05:36.75" />
                    <SPLIT distance="350" swimtime="00:06:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKO" nation="POL" region="WAR" clubid="9416" name="KS MAKO Warszawa">
          <CONTACT email="ania.plywanie@gmail.com" name="Anna Dąbrowska" phone="601 480 280" />
          <ATHLETES>
            <ATHLETE birthdate="1976-05-14" firstname="Dominik" gender="M" lastname="Markowski" nation="POL" athleteid="9438">
              <RESULTS>
                <RESULT eventid="8213" points="244" reactiontime="+87" swimtime="00:00:43.39" resultid="9439" heatid="14201" lane="4" entrytime="00:00:41.53" />
                <RESULT eventid="8277" points="227" reactiontime="+70" swimtime="00:01:25.34" resultid="9440" heatid="14226" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="243" reactiontime="+84" swimtime="00:01:35.80" resultid="9441" heatid="14244" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="9442" heatid="14310" lane="5" entrytime="00:01:40.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="9417">
              <RESULTS>
                <RESULT eventid="1075" points="890" reactiontime="+67" swimtime="00:00:23.00" resultid="9418" heatid="14161" lane="9" entrytime="00:00:23.90" />
                <RESULT eventid="8309" points="888" reactiontime="+73" swimtime="00:00:57.22" resultid="9419" heatid="14255" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="998" reactiontime="+73" swimtime="00:01:01.37" resultid="9420" heatid="14284" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="771" swimtime="00:00:24.94" resultid="9421" heatid="14302" lane="1" entrytime="00:00:25.50" />
                <RESULT eventid="8694" points="977" reactiontime="+67" swimtime="00:00:28.02" resultid="9422" heatid="14389" lane="3" entrytime="00:00:28.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarek" gender="M" lastname="Bystry" nation="POL" athleteid="9443">
              <RESULTS>
                <RESULT eventid="1075" points="620" reactiontime="+70" swimtime="00:00:27.85" resultid="9444" heatid="14153" lane="6" entrytime="00:00:28.20" />
                <RESULT eventid="8277" points="611" reactiontime="+80" swimtime="00:01:01.34" resultid="9445" heatid="14232" lane="5" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="529" reactiontime="+75" swimtime="00:01:13.96" resultid="9446" heatid="14249" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="528" reactiontime="+84" swimtime="00:00:31.09" resultid="9447" heatid="14298" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="8518" points="494" reactiontime="+71" swimtime="00:02:22.93" resultid="9448" heatid="14329" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:45.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-06-07" firstname="Piotr" gender="M" lastname="Kieżun" nation="POL" athleteid="9423">
              <RESULTS>
                <RESULT eventid="1075" points="399" reactiontime="+80" swimtime="00:00:31.22" resultid="9424" heatid="14147" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="8277" points="355" reactiontime="+105" swimtime="00:01:12.58" resultid="9425" heatid="14229" lane="0" entrytime="00:01:08.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="279" reactiontime="+79" swimtime="00:02:50.57" resultid="9426" heatid="14326" lane="8" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:02:05.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="9427">
              <RESULTS>
                <RESULT eventid="1075" points="298" reactiontime="+83" swimtime="00:00:38.02" resultid="9428" heatid="14145" lane="2" entrytime="00:00:39.37" />
                <RESULT eventid="8309" points="249" reactiontime="+85" swimtime="00:01:43.42" resultid="9429" heatid="14246" lane="0" entrytime="00:01:50.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="343" reactiontime="+88" swimtime="00:01:39.34" resultid="9430" heatid="14277" lane="3" entrytime="00:01:43.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="213" reactiontime="+81" swimtime="00:03:28.55" resultid="9431" heatid="14322" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:38.87" />
                    <SPLIT distance="150" swimtime="00:02:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8694" reactiontime="+50" status="DSQ" swimtime="00:00:00.00" resultid="9432" heatid="14381" lane="3" entrytime="00:00:45.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="9433">
              <RESULTS>
                <RESULT eventid="8277" points="307" reactiontime="+89" swimtime="00:01:18.42" resultid="9434" heatid="14226" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="285" reactiontime="+93" swimtime="00:01:31.20" resultid="9435" heatid="14245" lane="6" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="316" reactiontime="+109" swimtime="00:01:36.89" resultid="9436" heatid="14276" lane="5" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="248" reactiontime="+106" swimtime="00:03:02.46" resultid="9437" heatid="14323" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:01:28.77" />
                    <SPLIT distance="150" swimtime="00:02:15.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+76" swimtime="00:02:30.75" resultid="9449" heatid="14266" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:24.02" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9438" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="9427" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9443" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="9433" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8550" reactiontime="+70" status="DSQ" swimtime="00:01:55.66" resultid="9450" heatid="14338" lane="8" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.14" />
                    <SPLIT distance="100" swimtime="00:00:50.53" />
                    <SPLIT distance="150" swimtime="00:01:20.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9417" number="1" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="9443" number="2" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="9423" number="3" reactiontime="+33" status="DSQ" />
                    <RELAYPOSITION athleteid="9438" number="4" reactiontime="-43" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="10258" name="KS Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztoff" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="10285">
              <RESULTS>
                <RESULT eventid="1075" points="697" reactiontime="+80" swimtime="00:00:24.95" resultid="10286" heatid="14159" lane="4" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="545" reactiontime="+82" swimtime="00:02:24.60" resultid="10287" heatid="14171" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="728" reactiontime="+78" swimtime="00:00:29.45" resultid="10288" heatid="14206" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="8309" points="657" reactiontime="+80" swimtime="00:01:03.25" resultid="10289" heatid="14253" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="10290" heatid="14299" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="8486" points="721" reactiontime="+79" swimtime="00:01:04.18" resultid="10291" heatid="14314" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="649" reactiontime="+78" swimtime="00:01:00.76" resultid="10292" heatid="14358" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="643" reactiontime="+76" swimtime="00:00:32.22" resultid="10293" heatid="14386" lane="0" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="10264">
              <RESULTS>
                <RESULT eventid="1058" points="508" reactiontime="+84" swimtime="00:00:32.75" resultid="10265" heatid="14139" lane="1" entrytime="00:00:32.90" entrycourse="SCM" />
                <RESULT eventid="8229" status="DNS" swimtime="00:00:00.00" resultid="10266" heatid="14208" lane="9" />
                <RESULT eventid="8261" points="451" swimtime="00:01:14.90" resultid="10267" heatid="14221" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="391" reactiontime="+111" swimtime="00:01:30.92" resultid="10268" heatid="14303" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="433" swimtime="00:02:46.38" resultid="10269" heatid="14320" lane="0" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="396" reactiontime="+99" swimtime="00:03:12.70" resultid="10270" heatid="14364" lane="6" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                    <SPLIT distance="100" swimtime="00:01:34.79" />
                    <SPLIT distance="150" swimtime="00:02:23.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" license="102001600127" athleteid="10259">
              <RESULTS>
                <RESULT eventid="1058" points="815" reactiontime="+78" swimtime="00:00:27.98" resultid="10260" heatid="14134" lane="4" />
                <RESULT eventid="8261" points="803" reactiontime="+82" swimtime="00:01:01.83" resultid="10261" heatid="14223" lane="1" entrytime="00:01:04.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="731" reactiontime="+74" swimtime="00:01:16.86" resultid="10262" heatid="14274" lane="7" entrytime="00:01:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="725" reactiontime="+72" swimtime="00:00:34.89" resultid="10263" heatid="14378" lane="8" entrytime="00:00:35.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" license="102001700126" athleteid="10301">
              <RESULTS>
                <RESULT eventid="1075" points="831" reactiontime="+74" swimtime="00:00:24.46" resultid="10302" heatid="14142" lane="5" />
                <RESULT eventid="1105" points="919" reactiontime="+80" swimtime="00:02:10.93" resultid="10303" heatid="14174" lane="3" entrytime="00:02:13.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="100" swimtime="00:01:00.51" />
                    <SPLIT distance="150" swimtime="00:01:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="830" reactiontime="+70" swimtime="00:00:27.74" resultid="10304" heatid="14198" lane="3" />
                <RESULT comment="K1 - Pływak wykonał kopnięcie delfinowe po pierwszym kopnięciu do stylu klasycznego (pierwszy ruch po starcie lub nawrocie)., Z3" eventid="8309" reactiontime="+71" status="DSQ" swimtime="00:00:59.08" resultid="10305" heatid="14255" lane="9" entrytime="00:01:01.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="799" reactiontime="+84" swimtime="00:00:26.81" resultid="10306" heatid="14291" lane="0" />
                <RESULT eventid="8486" points="871" reactiontime="+86" swimtime="00:00:59.09" resultid="10307" heatid="14315" lane="3" entrytime="00:00:59.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="854" reactiontime="+76" swimtime="00:00:58.16" resultid="10308" heatid="14353" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="859" reactiontime="+63" swimtime="00:02:07.84" resultid="10665" heatid="14371" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:01.50" />
                    <SPLIT distance="150" swimtime="00:01:34.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="10280">
              <RESULTS>
                <RESULT eventid="1075" points="641" reactiontime="+85" swimtime="00:00:25.66" resultid="10281" heatid="14159" lane="6" entrytime="00:00:25.20" entrycourse="SCM" />
                <RESULT eventid="8245" points="664" reactiontime="+90" swimtime="00:02:41.03" resultid="10282" heatid="14216" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:15.69" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="664" reactiontime="+84" swimtime="00:01:10.31" resultid="10283" heatid="14283" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="702" reactiontime="+83" swimtime="00:00:31.29" resultid="10284" heatid="14389" lane="9" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="10271">
              <RESULTS>
                <RESULT eventid="1058" points="613" reactiontime="+74" swimtime="00:00:30.77" resultid="10272" heatid="14140" lane="6" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1135" points="613" reactiontime="+64" swimtime="00:11:11.11" resultid="10273" heatid="14178" lane="7" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:17.86" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                    <SPLIT distance="200" swimtime="00:02:44.15" />
                    <SPLIT distance="250" swimtime="00:03:27.11" />
                    <SPLIT distance="300" swimtime="00:04:09.54" />
                    <SPLIT distance="350" swimtime="00:04:52.10" />
                    <SPLIT distance="400" swimtime="00:05:34.43" />
                    <SPLIT distance="450" swimtime="00:06:16.67" />
                    <SPLIT distance="500" swimtime="00:06:59.34" />
                    <SPLIT distance="550" swimtime="00:07:41.35" />
                    <SPLIT distance="600" swimtime="00:08:23.45" />
                    <SPLIT distance="650" swimtime="00:09:05.89" />
                    <SPLIT distance="700" swimtime="00:09:47.86" />
                    <SPLIT distance="750" swimtime="00:10:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="584" reactiontime="+69" swimtime="00:03:02.76" resultid="10274" heatid="14211" lane="7" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                    <SPLIT distance="150" swimtime="00:02:14.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="464" reactiontime="+85" swimtime="00:03:04.70" resultid="10275" heatid="14257" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:25.65" />
                    <SPLIT distance="150" swimtime="00:02:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="545" reactiontime="+67" swimtime="00:01:24.76" resultid="10276" heatid="14273" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="605" reactiontime="+90" swimtime="00:05:59.97" resultid="10277" heatid="14342" lane="1" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:02:12.61" />
                    <SPLIT distance="200" swimtime="00:02:59.12" />
                    <SPLIT distance="250" swimtime="00:03:47.50" />
                    <SPLIT distance="300" swimtime="00:04:37.03" />
                    <SPLIT distance="350" swimtime="00:05:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="493" reactiontime="+74" swimtime="00:00:39.68" resultid="10278" heatid="14376" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="8726" points="617" reactiontime="+81" swimtime="00:05:21.18" resultid="10279" heatid="14393" lane="1" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:15.52" />
                    <SPLIT distance="150" swimtime="00:01:56.87" />
                    <SPLIT distance="200" swimtime="00:02:38.07" />
                    <SPLIT distance="250" swimtime="00:03:18.92" />
                    <SPLIT distance="300" swimtime="00:04:00.19" />
                    <SPLIT distance="350" swimtime="00:04:41.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="10294">
              <RESULTS>
                <RESULT eventid="1075" points="673" reactiontime="+65" swimtime="00:00:25.25" resultid="10295" heatid="14159" lane="9" entrytime="00:00:25.65" entrycourse="SCM" />
                <RESULT eventid="8277" points="629" reactiontime="+63" swimtime="00:00:57.22" resultid="10296" heatid="14235" lane="9" entrytime="00:00:58.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="595" reactiontime="+74" swimtime="00:01:05.38" resultid="10297" heatid="14252" lane="4" entrytime="00:01:07.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="517" reactiontime="+71" swimtime="00:00:28.48" resultid="10298" heatid="14299" lane="7" entrytime="00:00:28.84" />
                <RESULT eventid="8518" points="520" reactiontime="+85" swimtime="00:02:12.46" resultid="10299" heatid="14330" lane="1" entrytime="00:02:17.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="8694" reactiontime="+64" status="DSQ" swimtime="00:00:33.84" resultid="10300" heatid="14386" lane="6" entrytime="00:00:35.53" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+85" swimtime="00:01:38.32" resultid="10309" heatid="14339" lane="4" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.54" />
                    <SPLIT distance="100" swimtime="00:00:49.76" />
                    <SPLIT distance="150" swimtime="00:01:13.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10301" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="10280" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="10285" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10294" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8373" reactiontime="+64" swimtime="00:01:49.20" resultid="10310" heatid="14268" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                    <SPLIT distance="150" swimtime="00:01:24.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10301" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="10280" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="10285" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="10294" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+63" swimtime="00:02:01.43" resultid="10311" heatid="14392" lane="3" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="100" swimtime="00:01:02.45" />
                    <SPLIT distance="150" swimtime="00:01:29.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10301" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="10259" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="10285" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="10264" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1120" reactiontime="+69" swimtime="00:01:48.11" resultid="10312" heatid="14177" lane="6" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="100" swimtime="00:00:49.86" />
                    <SPLIT distance="150" swimtime="00:01:17.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10301" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="10280" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10259" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10271" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="11914" name="KS Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem jacek" phone="502 499 565" state="WIE" street="osiedle Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="11954">
              <RESULTS>
                <RESULT eventid="1150" points="450" reactiontime="+107" swimtime="00:12:47.97" resultid="11955" heatid="14185" lane="6" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:16.32" />
                    <SPLIT distance="200" swimtime="00:03:04.98" />
                    <SPLIT distance="250" swimtime="00:03:53.35" />
                    <SPLIT distance="300" swimtime="00:04:43.83" />
                    <SPLIT distance="350" swimtime="00:05:33.22" />
                    <SPLIT distance="400" swimtime="00:06:23.24" />
                    <SPLIT distance="450" swimtime="00:07:11.88" />
                    <SPLIT distance="500" swimtime="00:08:00.61" />
                    <SPLIT distance="550" swimtime="00:08:49.89" />
                    <SPLIT distance="600" swimtime="00:09:39.42" />
                    <SPLIT distance="650" swimtime="00:10:28.17" />
                    <SPLIT distance="700" swimtime="00:11:16.50" />
                    <SPLIT distance="750" swimtime="00:12:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="449" reactiontime="+106" swimtime="00:03:12.69" resultid="11956" heatid="14260" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:32.62" />
                    <SPLIT distance="150" swimtime="00:02:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="447" reactiontime="+108" swimtime="00:00:37.29" resultid="11957" heatid="14293" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="8518" points="480" reactiontime="+109" swimtime="00:02:47.34" resultid="11958" heatid="14326" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:05.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="454" reactiontime="+106" swimtime="00:01:24.27" resultid="11959" heatid="14356" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-01" firstname="Natalia" gender="F" lastname="Wiśniewska" nation="POL" license="500115600544" athleteid="11915">
              <RESULTS>
                <RESULT eventid="1090" points="784" reactiontime="+85" swimtime="00:02:29.71" resultid="11916" heatid="14165" lane="3" entrytime="00:02:29.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="730" reactiontime="+83" swimtime="00:10:08.43" resultid="11917" heatid="14178" lane="6" entrytime="00:10:15.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:49.57" />
                    <SPLIT distance="200" swimtime="00:02:27.90" />
                    <SPLIT distance="250" swimtime="00:03:06.67" />
                    <SPLIT distance="300" swimtime="00:03:44.77" />
                    <SPLIT distance="350" swimtime="00:04:23.52" />
                    <SPLIT distance="400" swimtime="00:05:02.03" />
                    <SPLIT distance="450" swimtime="00:05:40.80" />
                    <SPLIT distance="500" swimtime="00:06:19.59" />
                    <SPLIT distance="550" swimtime="00:06:58.48" />
                    <SPLIT distance="600" swimtime="00:07:37.05" />
                    <SPLIT distance="650" swimtime="00:08:15.50" />
                    <SPLIT distance="700" swimtime="00:08:53.92" />
                    <SPLIT distance="750" swimtime="00:09:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="796" reactiontime="+82" swimtime="00:02:43.86" resultid="11918" heatid="14211" lane="4" entrytime="00:02:44.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="746" reactiontime="+81" swimtime="00:01:09.65" resultid="11919" heatid="14243" lane="6" entrytime="00:01:09.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="840" reactiontime="+84" swimtime="00:01:14.94" resultid="11920" heatid="14274" lane="4" entrytime="00:01:15.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="812" reactiontime="+88" swimtime="00:05:23.28" resultid="11921" heatid="14342" lane="3" entrytime="00:05:25.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                    <SPLIT distance="200" swimtime="00:02:35.52" />
                    <SPLIT distance="250" swimtime="00:03:19.14" />
                    <SPLIT distance="300" swimtime="00:04:03.59" />
                    <SPLIT distance="350" swimtime="00:04:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="746" reactiontime="+78" swimtime="00:01:08.50" resultid="11922" heatid="14352" lane="5" entrytime="00:01:09.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="845" reactiontime="+78" swimtime="00:00:34.73" resultid="11923" heatid="14378" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="11924">
              <RESULTS>
                <RESULT eventid="1075" points="753" reactiontime="+84" swimtime="00:00:27.93" resultid="11925" heatid="14154" lane="1" entrytime="00:00:27.95" />
                <RESULT eventid="1150" points="656" reactiontime="+95" swimtime="00:10:18.67" resultid="11926" heatid="14182" lane="0" entrytime="00:10:15.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:49.68" />
                    <SPLIT distance="200" swimtime="00:02:28.15" />
                    <SPLIT distance="250" swimtime="00:03:06.69" />
                    <SPLIT distance="300" swimtime="00:03:45.37" />
                    <SPLIT distance="350" swimtime="00:04:24.27" />
                    <SPLIT distance="400" swimtime="00:05:03.67" />
                    <SPLIT distance="450" swimtime="00:05:42.93" />
                    <SPLIT distance="500" swimtime="00:06:22.67" />
                    <SPLIT distance="550" swimtime="00:07:02.67" />
                    <SPLIT distance="600" swimtime="00:07:42.32" />
                    <SPLIT distance="650" swimtime="00:08:22.07" />
                    <SPLIT distance="700" swimtime="00:09:01.84" />
                    <SPLIT distance="750" swimtime="00:09:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="785" reactiontime="+66" swimtime="00:00:31.71" resultid="11927" heatid="14205" lane="5" entrytime="00:00:31.40" />
                <RESULT eventid="8486" points="751" reactiontime="+90" swimtime="00:01:10.00" resultid="11928" heatid="14314" lane="8" entrytime="00:01:09.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="701" reactiontime="+95" swimtime="00:02:20.20" resultid="11929" heatid="14330" lane="0" entrytime="00:02:18.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="721" reactiontime="+85" swimtime="00:02:35.14" resultid="11930" heatid="14370" lane="1" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="668" reactiontime="+90" swimtime="00:04:57.92" resultid="11931" heatid="14400" lane="7" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:49.10" />
                    <SPLIT distance="200" swimtime="00:02:27.27" />
                    <SPLIT distance="250" swimtime="00:03:05.58" />
                    <SPLIT distance="300" swimtime="00:03:44.15" />
                    <SPLIT distance="350" swimtime="00:04:22.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-31" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" license="500115700461" athleteid="11977">
              <RESULTS>
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="11978" heatid="14217" lane="9" entrytime="00:02:42.14" />
                <RESULT eventid="8406" points="794" reactiontime="+72" swimtime="00:01:10.84" resultid="11979" heatid="14283" lane="6" entrytime="00:01:11.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Szymon" gender="M" lastname="Wieja" nation="POL" license="500115700467" athleteid="11932">
              <RESULTS>
                <RESULT eventid="1075" points="751" reactiontime="+71" swimtime="00:00:26.13" resultid="11933" heatid="14159" lane="1" entrytime="00:00:25.40" />
                <RESULT eventid="1105" points="707" reactiontime="+73" swimtime="00:02:23.54" resultid="11934" heatid="14173" lane="3" entrytime="00:02:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="696" reactiontime="+78" swimtime="00:00:30.63" resultid="11935" heatid="14207" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="8277" points="757" reactiontime="+81" swimtime="00:00:57.12" resultid="11936" heatid="14236" lane="0" entrytime="00:00:57.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="700" reactiontime="+76" swimtime="00:01:06.51" resultid="11937" heatid="14314" lane="7" entrytime="00:01:08.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="11938" heatid="14348" lane="0" entrytime="00:05:21.30" />
                <RESULT eventid="8662" points="711" reactiontime="+71" swimtime="00:02:26.13" resultid="11939" heatid="14370" lane="5" entrytime="00:02:29.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="577" reactiontime="+68" swimtime="00:04:49.03" resultid="11940" heatid="14399" lane="8" entrytime="00:04:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                    <SPLIT distance="150" swimtime="00:01:46.26" />
                    <SPLIT distance="200" swimtime="00:02:23.79" />
                    <SPLIT distance="250" swimtime="00:03:01.17" />
                    <SPLIT distance="300" swimtime="00:03:38.29" />
                    <SPLIT distance="350" swimtime="00:04:15.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-12" firstname="Marcin" gender="M" lastname="Szymkowiak" nation="POL" license="500115700523" athleteid="11941">
              <RESULTS>
                <RESULT eventid="1075" points="723" reactiontime="+75" swimtime="00:00:25.62" resultid="11942" heatid="14159" lane="8" entrytime="00:00:25.40" />
                <RESULT eventid="1105" points="719" reactiontime="+80" swimtime="00:02:22.07" resultid="11943" heatid="14173" lane="6" entrytime="00:02:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="772" reactiontime="+73" swimtime="00:02:33.20" resultid="11944" heatid="14217" lane="6" entrytime="00:02:33.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8406" points="861" reactiontime="+81" swimtime="00:01:07.28" resultid="11945" heatid="14284" lane="0" entrytime="00:01:06.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="703" reactiontime="+79" swimtime="00:00:27.98" resultid="11946" heatid="14300" lane="3" entrytime="00:00:27.50" />
                <RESULT comment="Rekord Polski" eventid="8694" points="875" reactiontime="+70" swimtime="00:00:30.18" resultid="11947" heatid="14389" lane="8" entrytime="00:00:29.99" />
                <RESULT eventid="8742" points="631" reactiontime="+65" swimtime="00:04:42.47" resultid="11948" heatid="14399" lane="5" entrytime="00:04:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:41.70" />
                    <SPLIT distance="200" swimtime="00:02:17.89" />
                    <SPLIT distance="250" swimtime="00:02:54.75" />
                    <SPLIT distance="300" swimtime="00:03:31.41" />
                    <SPLIT distance="350" swimtime="00:04:07.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-17" firstname="Magdalena" gender="F" lastname="Zajączek" nation="POL" license="500115600524" athleteid="11989">
              <RESULTS>
                <RESULT eventid="1058" points="148" swimtime="00:00:51.32" resultid="11990" heatid="14135" lane="7" entrytime="00:00:53.93" />
                <RESULT eventid="8229" points="246" swimtime="00:04:24.96" resultid="11991" heatid="14209" lane="0" entrytime="00:04:17.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.70" />
                    <SPLIT distance="100" swimtime="00:02:08.14" />
                    <SPLIT distance="150" swimtime="00:03:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="213" swimtime="00:02:06.69" resultid="11992" heatid="14270" lane="6" entrytime="00:02:03.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="198" swimtime="00:00:58.89" resultid="11993" heatid="14373" lane="1" entrytime="00:00:58.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-05" firstname="Filip" gender="M" lastname="Piotrowski" nation="POL" license="500115700522" athleteid="11949">
              <RESULTS>
                <RESULT eventid="1075" points="645" reactiontime="+90" swimtime="00:00:27.49" resultid="11950" heatid="14159" lane="0" entrytime="00:00:25.40" />
                <RESULT eventid="8277" points="643" reactiontime="+65" swimtime="00:01:00.30" resultid="11951" heatid="14236" lane="9" entrytime="00:00:57.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="571" reactiontime="+77" swimtime="00:00:30.29" resultid="11952" heatid="14300" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="8630" points="631" reactiontime="+62" swimtime="00:01:06.00" resultid="11953" heatid="14359" lane="3" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" license="500115600462" athleteid="11980">
              <RESULTS>
                <RESULT eventid="1090" points="324" swimtime="00:03:55.76" resultid="11981" heatid="14163" lane="0" entrytime="00:03:56.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                    <SPLIT distance="100" swimtime="00:01:55.00" />
                    <SPLIT distance="150" swimtime="00:02:59.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="293" reactiontime="+105" swimtime="00:15:17.25" resultid="11982" heatid="14180" lane="2" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:38.60" />
                    <SPLIT distance="200" swimtime="00:03:36.96" />
                    <SPLIT distance="250" swimtime="00:04:35.42" />
                    <SPLIT distance="300" swimtime="00:05:34.05" />
                    <SPLIT distance="350" swimtime="00:06:34.18" />
                    <SPLIT distance="400" swimtime="00:07:34.11" />
                    <SPLIT distance="450" swimtime="00:08:32.19" />
                    <SPLIT distance="500" swimtime="00:09:30.82" />
                    <SPLIT distance="550" swimtime="00:10:28.69" />
                    <SPLIT distance="600" swimtime="00:11:26.33" />
                    <SPLIT distance="650" swimtime="00:12:24.65" />
                    <SPLIT distance="700" swimtime="00:13:23.45" />
                    <SPLIT distance="750" swimtime="00:14:21.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="410" reactiontime="+91" swimtime="00:04:09.24" resultid="11983" heatid="14209" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.69" />
                    <SPLIT distance="100" swimtime="00:01:57.56" />
                    <SPLIT distance="150" swimtime="00:03:03.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="290" reactiontime="+115" swimtime="00:04:27.83" resultid="11984" heatid="14256" lane="2" entrytime="00:04:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                    <SPLIT distance="100" swimtime="00:02:05.13" />
                    <SPLIT distance="150" swimtime="00:03:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="488" reactiontime="+106" swimtime="00:01:46.28" resultid="11985" heatid="14270" lane="4" entrytime="00:02:01.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="432" swimtime="00:08:09.09" resultid="11986" heatid="14340" lane="3" entrytime="00:08:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:02:04.62" />
                    <SPLIT distance="150" swimtime="00:03:07.09" />
                    <SPLIT distance="200" swimtime="00:04:07.40" />
                    <SPLIT distance="250" swimtime="00:05:12.00" />
                    <SPLIT distance="300" swimtime="00:06:16.33" />
                    <SPLIT distance="350" swimtime="00:07:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="257" swimtime="00:02:03.62" resultid="11987" heatid="14350" lane="7" entrytime="00:01:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="335" reactiontime="+113" swimtime="00:03:56.76" resultid="11988" heatid="14363" lane="8" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:55.61" />
                    <SPLIT distance="150" swimtime="00:02:57.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" license="500115600525" athleteid="12029">
              <RESULTS>
                <RESULT eventid="1058" points="115" reactiontime="+112" swimtime="00:00:55.79" resultid="12030" heatid="14135" lane="8" entrytime="00:00:57.00" />
                <RESULT eventid="8229" points="244" reactiontime="+126" swimtime="00:04:25.68" resultid="12031" heatid="14208" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.19" />
                    <SPLIT distance="100" swimtime="00:02:06.70" />
                    <SPLIT distance="150" swimtime="00:03:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="87" reactiontime="+117" swimtime="00:02:14.06" resultid="12032" heatid="14218" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="212" reactiontime="+110" swimtime="00:02:06.90" resultid="12033" heatid="14270" lane="3" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="217" reactiontime="+110" swimtime="00:00:57.13" resultid="12034" heatid="14373" lane="5" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" license="500115600520" athleteid="12009">
              <RESULTS>
                <RESULT eventid="1058" points="398" reactiontime="+116" swimtime="00:00:43.81" resultid="12010" heatid="14136" lane="9" entrytime="00:00:46.00" />
                <RESULT eventid="8229" points="575" reactiontime="+109" swimtime="00:04:01.41" resultid="12011" heatid="14209" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.49" />
                    <SPLIT distance="100" swimtime="00:01:54.14" />
                    <SPLIT distance="150" swimtime="00:02:58.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="333" reactiontime="+120" swimtime="00:01:42.34" resultid="12012" heatid="14219" lane="0" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="547" reactiontime="+116" swimtime="00:01:51.39" resultid="12013" heatid="14271" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="387" reactiontime="+124" swimtime="00:03:44.96" resultid="12014" heatid="14317" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:01:49.99" />
                    <SPLIT distance="150" swimtime="00:02:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="533" reactiontime="+117" swimtime="00:00:50.84" resultid="12015" heatid="14374" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-08" firstname="Błażej" gender="M" lastname="Wachowski" nation="POL" license="100115700545" athleteid="12023">
              <RESULTS>
                <RESULT eventid="1150" points="507" reactiontime="+99" swimtime="00:10:43.50" resultid="12024" heatid="14182" lane="9" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:01:55.31" />
                    <SPLIT distance="200" swimtime="00:02:36.44" />
                    <SPLIT distance="250" swimtime="00:03:17.39" />
                    <SPLIT distance="300" swimtime="00:03:58.56" />
                    <SPLIT distance="350" swimtime="00:04:39.12" />
                    <SPLIT distance="400" swimtime="00:05:20.13" />
                    <SPLIT distance="450" swimtime="00:06:01.43" />
                    <SPLIT distance="500" swimtime="00:06:42.17" />
                    <SPLIT distance="550" swimtime="00:07:22.74" />
                    <SPLIT distance="600" swimtime="00:08:03.40" />
                    <SPLIT distance="650" swimtime="00:08:44.30" />
                    <SPLIT distance="700" swimtime="00:09:25.22" />
                    <SPLIT distance="750" swimtime="00:10:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="412" reactiontime="+108" swimtime="00:02:50.09" resultid="12025" heatid="14261" lane="0" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:02.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="463" reactiontime="+93" swimtime="00:02:24.02" resultid="12026" heatid="14329" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="428" reactiontime="+96" swimtime="00:01:13.20" resultid="12027" heatid="14356" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="467" reactiontime="+105" swimtime="00:05:12.33" resultid="12028" heatid="14400" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:54.60" />
                    <SPLIT distance="200" swimtime="00:02:34.66" />
                    <SPLIT distance="250" swimtime="00:03:15.30" />
                    <SPLIT distance="300" swimtime="00:03:54.92" />
                    <SPLIT distance="350" swimtime="00:04:34.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-11" firstname="Piotr" gender="M" lastname="Witt" nation="POL" license="500115700548" athleteid="12016">
              <RESULTS>
                <RESULT eventid="1075" points="749" reactiontime="+79" swimtime="00:00:25.15" resultid="12017" heatid="14160" lane="2" entrytime="00:00:24.40" />
                <RESULT eventid="8213" points="597" reactiontime="+84" swimtime="00:00:29.75" resultid="12018" heatid="14206" lane="7" entrytime="00:00:30.59" />
                <RESULT eventid="8277" points="725" reactiontime="+71" swimtime="00:00:54.07" resultid="12019" heatid="14237" lane="8" entrytime="00:00:54.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="607" reactiontime="+74" swimtime="00:00:27.98" resultid="12020" heatid="14300" lane="4" entrytime="00:00:27.49" />
                <RESULT eventid="8518" points="680" reactiontime="+70" swimtime="00:02:07.97" resultid="12021" heatid="14332" lane="8" entrytime="00:02:08.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                    <SPLIT distance="150" swimtime="00:01:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="566" reactiontime="+75" swimtime="00:01:05.19" resultid="12022" heatid="14359" lane="9" entrytime="00:01:05.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" license="100115600353" athleteid="11969">
              <RESULTS>
                <RESULT eventid="1135" points="335" reactiontime="+109" swimtime="00:17:18.49" resultid="11970" heatid="14180" lane="8" entrytime="00:18:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:49.33" />
                    <SPLIT distance="400" swimtime="00:08:26.64" />
                    <SPLIT distance="650" swimtime="00:14:03.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="298" reactiontime="+124" swimtime="00:04:40.51" resultid="11971" heatid="14208" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.86" />
                    <SPLIT distance="100" swimtime="00:02:09.70" />
                    <SPLIT distance="150" swimtime="00:03:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="302" reactiontime="+124" swimtime="00:01:46.39" resultid="11972" heatid="14218" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="11973" heatid="14270" lane="5" entrytime="00:02:02.00" />
                <RESULT eventid="8502" points="273" reactiontime="+129" swimtime="00:04:04.78" resultid="11974" heatid="14317" lane="7" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.09" />
                    <SPLIT distance="100" swimtime="00:01:53.37" />
                    <SPLIT distance="150" swimtime="00:02:59.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="11975" heatid="14362" lane="5" entrytime="00:04:55.00" />
                <RESULT eventid="8678" points="319" reactiontime="+113" swimtime="00:00:56.12" resultid="11976" heatid="14373" lane="6" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="12000">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="12001" heatid="14174" lane="7" entrytime="00:02:20.00" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="12002" heatid="14182" lane="5" entrytime="00:09:10.00" />
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="12003" heatid="14217" lane="2" entrytime="00:02:34.00" />
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="12004" heatid="14262" lane="7" entrytime="00:02:20.00" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="12005" heatid="14332" lane="5" entrytime="00:02:06.00" />
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="12006" heatid="14348" lane="6" entrytime="00:05:00.00" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="12007" heatid="14360" lane="1" entrytime="00:01:02.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="11961">
              <RESULTS>
                <RESULT eventid="1135" points="396" swimtime="00:13:16.26" resultid="11962" heatid="14179" lane="8" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:28.25" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                    <SPLIT distance="200" swimtime="00:03:06.39" />
                    <SPLIT distance="250" swimtime="00:03:55.28" />
                    <SPLIT distance="300" swimtime="00:04:45.47" />
                    <SPLIT distance="350" swimtime="00:05:35.77" />
                    <SPLIT distance="400" swimtime="00:06:26.89" />
                    <SPLIT distance="450" swimtime="00:07:18.29" />
                    <SPLIT distance="500" swimtime="00:08:09.78" />
                    <SPLIT distance="550" swimtime="00:09:01.11" />
                    <SPLIT distance="600" swimtime="00:09:51.85" />
                    <SPLIT distance="650" swimtime="00:10:42.39" />
                    <SPLIT distance="700" swimtime="00:11:34.13" />
                    <SPLIT distance="750" swimtime="00:12:26.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="350" reactiontime="+124" swimtime="00:00:47.11" resultid="11963" heatid="14194" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="8261" points="397" swimtime="00:01:24.24" resultid="11964" heatid="14219" lane="5" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="353" reactiontime="+116" swimtime="00:01:42.15" resultid="11965" heatid="14305" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" status="DNS" swimtime="00:00:00.00" resultid="11966" heatid="14318" lane="5" entrytime="00:03:10.00" />
                <RESULT eventid="8646" points="411" reactiontime="+132" swimtime="00:03:31.69" resultid="11967" heatid="14363" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:43.44" />
                    <SPLIT distance="150" swimtime="00:02:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="388" swimtime="00:06:32.43" resultid="11968" heatid="14395" lane="0" entrytime="00:06:21.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.46" />
                    <SPLIT distance="250" swimtime="00:03:59.17" />
                    <SPLIT distance="300" swimtime="00:04:50.78" />
                    <SPLIT distance="350" swimtime="00:05:41.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" license="500115700493" athleteid="11994">
              <RESULTS>
                <RESULT eventid="1058" points="628" reactiontime="+96" swimtime="00:00:36.21" resultid="11995" heatid="14138" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="8229" points="737" reactiontime="+89" swimtime="00:03:27.46" resultid="11996" heatid="14210" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="704" reactiontime="+88" swimtime="00:01:28.88" resultid="11997" heatid="14240" lane="8" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="739" reactiontime="+98" swimtime="00:01:35.00" resultid="11998" heatid="14272" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="706" reactiontime="+85" swimtime="00:00:43.10" resultid="11999" heatid="14377" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="SZYMKOWIAK TEAM" number="4">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+93" swimtime="00:01:57.77" resultid="12038" heatid="14268" lane="1" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:02.66" />
                    <SPLIT distance="150" swimtime="00:01:31.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11924" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="11941" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="11949" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="11932" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="OD A DO Z" number="5">
              <RESULTS>
                <RESULT eventid="8373" status="DNS" swimtime="00:00:00.00" resultid="12039" heatid="14266" lane="5" entrytime="00:02:12.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12016" number="1" />
                    <RELAYPOSITION athleteid="11977" number="2" />
                    <RELAYPOSITION athleteid="12023" number="3" />
                    <RELAYPOSITION athleteid="11954" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="ASY SPRINTU" number="7">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+77" swimtime="00:01:43.02" resultid="12042" heatid="14339" lane="2" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.91" />
                    <SPLIT distance="100" swimtime="00:00:50.90" />
                    <SPLIT distance="150" swimtime="00:01:17.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12016" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="11932" number="2" reactiontime="+17" />
                    <RELAYPOSITION athleteid="11949" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="11941" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="PANIE ZMIENNE" number="3">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+113" swimtime="00:03:04.68" resultid="12037" heatid="14263" lane="6" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:30.73" />
                    <SPLIT distance="150" swimtime="00:02:19.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11961" number="1" reactiontime="+113" />
                    <RELAYPOSITION athleteid="11994" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="11980" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="12009" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="GWIAZDY" number="6">
              <RESULTS>
                <RESULT eventid="8534" status="DNS" swimtime="00:00:00.00" resultid="12040" heatid="14334" lane="4" entrytime="00:02:35.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11961" number="1" />
                    <RELAYPOSITION athleteid="11994" number="2" />
                    <RELAYPOSITION athleteid="12009" number="3" />
                    <RELAYPOSITION athleteid="11980" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="ANIA TEAM" number="1">
              <RESULTS>
                <RESULT eventid="1120" swimtime="00:02:11.44" resultid="12035" heatid="14176" lane="8" entrytime="00:02:06.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:06.43" />
                    <SPLIT distance="150" swimtime="00:01:42.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11961" number="1" />
                    <RELAYPOSITION athleteid="11949" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="11994" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="11924" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="THIEM TEAM" number="2">
              <RESULTS>
                <RESULT eventid="1120" swimtime="00:02:40.28" resultid="12036" heatid="14175" lane="1" entrytime="00:02:53.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11989" number="1" />
                    <RELAYPOSITION athleteid="12023" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="11969" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="11954" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="MASA KRYTYCZNA" number="8">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8710" reactiontime="+95" status="DSQ" swimtime="00:02:38.44" resultid="12041" heatid="14390" lane="3" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="100" swimtime="00:01:44.75" />
                    <SPLIT distance="150" swimtime="00:02:13.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11980" number="1" reactiontime="+95" status="DSQ" />
                    <RELAYPOSITION athleteid="12029" number="2" reactiontime="+80" status="DSQ" />
                    <RELAYPOSITION athleteid="11949" number="3" reactiontime="-4" status="DSQ" />
                    <RELAYPOSITION athleteid="12016" number="4" reactiontime="+38" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="9085" name="KS_Niezrzeszeni_pl">
          <CONTACT name="KS_Niezrzeszeni_pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="9086">
              <RESULTS>
                <RESULT eventid="1075" points="433" reactiontime="+94" swimtime="00:00:34.46" resultid="9087" heatid="14146" lane="7" entrytime="00:00:35.32" />
                <RESULT eventid="1150" points="469" reactiontime="+125" swimtime="00:12:37.83" resultid="9088" heatid="14185" lane="1" entrytime="00:13:08.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:18.37" />
                    <SPLIT distance="200" swimtime="00:03:06.91" />
                    <SPLIT distance="250" swimtime="00:03:55.80" />
                    <SPLIT distance="300" swimtime="00:04:44.19" />
                    <SPLIT distance="350" swimtime="00:05:32.69" />
                    <SPLIT distance="400" swimtime="00:06:21.53" />
                    <SPLIT distance="450" swimtime="00:07:10.28" />
                    <SPLIT distance="500" swimtime="00:07:58.54" />
                    <SPLIT distance="550" swimtime="00:08:46.57" />
                    <SPLIT distance="600" swimtime="00:09:34.88" />
                    <SPLIT distance="650" swimtime="00:10:23.09" />
                    <SPLIT distance="700" swimtime="00:11:10.95" />
                    <SPLIT distance="750" swimtime="00:11:57.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="346" reactiontime="+111" swimtime="00:01:33.63" resultid="9089" heatid="14244" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="288" reactiontime="+110" swimtime="00:00:43.16" resultid="9090" heatid="14292" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="8486" points="358" reactiontime="+80" swimtime="00:01:31.15" resultid="9091" heatid="14311" lane="6" entrytime="00:01:27.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="429" reactiontime="+75" swimtime="00:03:09.89" resultid="9092" heatid="14366" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.82" />
                    <SPLIT distance="100" swimtime="00:02:22.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="430" reactiontime="+106" swimtime="00:06:15.47" resultid="9093" heatid="14404" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:28.51" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                    <SPLIT distance="200" swimtime="00:03:05.83" />
                    <SPLIT distance="250" swimtime="00:03:55.08" />
                    <SPLIT distance="300" swimtime="00:04:44.19" />
                    <SPLIT distance="350" swimtime="00:05:32.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="WIE" clubid="10916" name="KU AZS UAM Poznań">
          <CONTACT email="swimteamuam@gmail.com" name="Sterczyński" phone="693840114" />
          <ATHLETES>
            <ATHLETE birthdate="1981-06-05" firstname="Marek" gender="M" lastname="Serafin" nation="POL" athleteid="10952">
              <RESULTS>
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="10953" heatid="14228" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="10954" heatid="14292" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="10955" heatid="14326" lane="4" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-27" firstname="Bartosz" gender="M" lastname="Kaczmarek" nation="POL" athleteid="10968">
              <RESULTS>
                <RESULT eventid="1075" points="492" reactiontime="+67" swimtime="00:00:29.13" resultid="10969" heatid="14152" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="8277" points="474" reactiontime="+71" swimtime="00:01:05.92" resultid="10970" heatid="14229" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="325" reactiontime="+78" swimtime="00:01:22.53" resultid="10971" heatid="14248" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="347" reactiontime="+80" swimtime="00:02:38.53" resultid="10972" heatid="14328" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:57.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" license="103315200006" athleteid="10946">
              <RESULTS>
                <RESULT eventid="1075" points="752" reactiontime="+66" swimtime="00:00:25.11" resultid="10947" heatid="14161" lane="6" entrytime="00:00:23.40" />
                <RESULT eventid="8213" points="808" reactiontime="+67" swimtime="00:00:26.89" resultid="10948" heatid="14207" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10949" heatid="14255" lane="7" entrytime="00:00:59.00" />
                <RESULT comment="Rekord Polski" eventid="8454" points="901" swimtime="00:00:24.53" resultid="10950" heatid="14302" lane="5" entrytime="00:00:24.50" />
                <RESULT eventid="8630" points="863" reactiontime="+65" swimtime="00:00:56.64" resultid="10951" heatid="14361" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-19" firstname="Damian" gender="M" lastname="Kowalik" nation="POL" license="103315200009" athleteid="10941">
              <RESULTS>
                <RESULT eventid="1075" points="802" reactiontime="+69" swimtime="00:00:24.69" resultid="10942" heatid="14161" lane="1" entrytime="00:00:23.73" />
                <RESULT eventid="8277" points="753" reactiontime="+66" swimtime="00:00:55.68" resultid="10943" heatid="14236" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="880" swimtime="00:00:25.83" resultid="10944" heatid="14302" lane="6" entrytime="00:00:25.00" />
                <RESULT eventid="8630" points="747" reactiontime="+63" swimtime="00:00:59.85" resultid="10945" heatid="14361" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-01" firstname="Dariusz" gender="M" lastname="Perkowski" nation="POL" athleteid="10917">
              <RESULTS>
                <RESULT eventid="1075" points="396" reactiontime="+69" swimtime="00:00:32.35" resultid="10918" heatid="14150" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="8277" points="285" reactiontime="+82" swimtime="00:01:19.07" resultid="10919" heatid="14228" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="222" reactiontime="+77" swimtime="00:01:38.76" resultid="10920" heatid="14247" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="294" reactiontime="+66" swimtime="00:00:37.79" resultid="10921" heatid="14294" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="10936">
              <RESULTS>
                <RESULT eventid="1075" points="484" reactiontime="+90" swimtime="00:00:29.29" resultid="10937" heatid="14152" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="8277" points="470" reactiontime="+78" swimtime="00:01:06.11" resultid="10938" heatid="14230" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="423" reactiontime="+88" swimtime="00:01:15.62" resultid="10939" heatid="14248" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="395" reactiontime="+88" swimtime="00:00:33.90" resultid="10940" heatid="14294" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-20" firstname="Krzysztof" gender="M" lastname="Strzelczyk" nation="POL" athleteid="10922">
              <RESULTS>
                <RESULT eventid="1075" points="330" reactiontime="+90" swimtime="00:00:34.38" resultid="10923" heatid="14146" lane="5" entrytime="00:00:34.88" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="10924" heatid="14185" lane="8" entrytime="00:13:30.00" />
                <RESULT eventid="8277" points="302" reactiontime="+89" swimtime="00:01:17.60" resultid="10925" heatid="14226" lane="6" entrytime="00:01:22.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="244" reactiontime="+98" swimtime="00:01:35.62" resultid="10926" heatid="14246" lane="5" entrytime="00:01:38.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="242" reactiontime="+80" swimtime="00:00:40.32" resultid="10927" heatid="14292" lane="8" entrytime="00:00:43.62" />
                <RESULT eventid="8518" points="265" reactiontime="+94" swimtime="00:02:55.95" resultid="10928" heatid="14325" lane="0" entrytime="00:03:09.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:10.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-13" firstname="Kamil" gender="M" lastname="Bernaś" nation="POL" athleteid="10930">
              <RESULTS>
                <RESULT eventid="1075" points="532" reactiontime="+74" swimtime="00:00:27.31" resultid="10931" heatid="14154" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="8277" points="488" reactiontime="+72" swimtime="00:01:02.28" resultid="10932" heatid="14231" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="407" reactiontime="+74" swimtime="00:01:14.19" resultid="10933" heatid="14248" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="432" reactiontime="+70" swimtime="00:00:30.25" resultid="10934" heatid="14298" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="8630" points="301" reactiontime="+70" swimtime="00:01:18.49" resultid="10935" heatid="14358" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="10963">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="10964" heatid="14173" lane="8" entrytime="00:02:30.00" />
                <RESULT eventid="8309" points="616" reactiontime="+69" swimtime="00:01:04.62" resultid="10965" heatid="14254" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="528" reactiontime="+70" swimtime="00:00:28.28" resultid="10966" heatid="14299" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="8630" points="535" reactiontime="+73" swimtime="00:01:04.83" resultid="10967" heatid="14359" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Sterczyńska" nation="POL" athleteid="10957">
              <RESULTS>
                <RESULT eventid="1058" points="830" reactiontime="+80" swimtime="00:00:27.40" resultid="10958" heatid="14141" lane="5" entrytime="00:00:27.58" />
                <RESULT eventid="8261" points="830" reactiontime="+81" swimtime="00:00:59.71" resultid="10959" heatid="14223" lane="6" entrytime="00:01:00.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="850" reactiontime="+81" swimtime="00:01:08.87" resultid="10960" heatid="14243" lane="7" entrytime="00:01:10.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="755" reactiontime="+83" swimtime="00:00:30.81" resultid="10961" heatid="14289" lane="6" entrytime="00:00:30.70" />
                <RESULT eventid="8678" points="671" reactiontime="+77" swimtime="00:00:36.07" resultid="10962" heatid="14378" lane="1" entrytime="00:00:35.91" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+82" swimtime="00:01:46.73" resultid="10974" heatid="14338" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:00:56.42" />
                    <SPLIT distance="150" swimtime="00:01:22.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10936" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="10930" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="10963" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="10946" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8373" reactiontime="+71" swimtime="00:01:59.22" resultid="10975" heatid="14268" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:59.54" />
                    <SPLIT distance="150" swimtime="00:01:30.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10946" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="10963" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="10930" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="10936" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="8550" swimtime="00:01:59.97" resultid="10976" heatid="14337" lane="7" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:30.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10922" number="1" />
                    <RELAYPOSITION athleteid="10917" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="10941" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10968" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8373" reactiontime="+89" swimtime="00:02:18.81" resultid="10977" heatid="14266" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:21.37" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10968" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="10922" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="10941" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="10917" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="8860" name="Kúpele Piešťany">
          <ATHLETES>
            <ATHLETE birthdate="1961-04-20" firstname="Anna" gender="F" lastname="Kičínová" nation="SVK" athleteid="9042">
              <RESULTS>
                <RESULT eventid="8678" points="631" reactiontime="+81" swimtime="00:00:43.78" resultid="9043" heatid="14375" lane="2" entrytime="00:00:43.70" />
                <RESULT eventid="8404" points="674" reactiontime="+97" swimtime="00:01:35.42" resultid="9044" heatid="14272" lane="2" entrytime="00:01:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="714" reactiontime="+98" swimtime="00:03:27.25" resultid="9045" heatid="14210" lane="2" entrytime="00:03:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:38.93" />
                    <SPLIT distance="150" swimtime="00:02:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="533" reactiontime="+95" swimtime="00:00:40.38" resultid="9046" heatid="14287" lane="1" entrytime="00:00:38.20" />
                <RESULT eventid="8613" points="726" reactiontime="+90" swimtime="00:01:27.53" resultid="9047" heatid="14351" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="673" reactiontime="+91" swimtime="00:03:22.29" resultid="9048" heatid="14257" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="541" reactiontime="+92" swimtime="00:03:18.91" resultid="9049" heatid="14163" lane="3" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:01:32.33" />
                    <SPLIT distance="150" swimtime="00:02:26.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-11-28" firstname="Karol" gender="M" lastname="Kantek" nation="SVK" athleteid="8861">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1075" reactiontime="+69" status="DSQ" swimtime="00:00:31.92" resultid="8862" heatid="14148" lane="5" entrytime="00:00:31.94" />
                <RESULT eventid="8213" points="658" reactiontime="+72" swimtime="00:00:39.87" resultid="8863" heatid="14202" lane="8" entrytime="00:00:40.20" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="8864" heatid="14294" lane="9" entrytime="00:00:35.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol" gender="M" lastname="Škodný" nation="SVK" athleteid="9050">
              <RESULTS>
                <RESULT eventid="8213" points="584" reactiontime="+79" swimtime="00:00:33.33" resultid="9051" heatid="14204" lane="7" entrytime="00:00:33.20" />
                <RESULT eventid="8486" points="544" reactiontime="+104" swimtime="00:01:12.85" resultid="9052" heatid="14313" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="678" reactiontime="+83" swimtime="00:02:35.09" resultid="9053" heatid="14370" lane="8" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="699" reactiontime="+91" swimtime="00:02:32.38" resultid="9054" heatid="14172" lane="7" entrytime="00:02:35.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="622" reactiontime="+98" swimtime="00:05:38.49" resultid="9055" heatid="14347" lane="6" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:59.75" />
                    <SPLIT distance="200" swimtime="00:02:42.49" />
                    <SPLIT distance="250" swimtime="00:03:30.82" />
                    <SPLIT distance="300" swimtime="00:04:20.78" />
                    <SPLIT distance="350" swimtime="00:05:00.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="499" reactiontime="+100" swimtime="00:02:45.90" resultid="9056" heatid="14261" lane="9" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="558" reactiontime="+110" swimtime="00:10:31.17" resultid="9057" heatid="14183" lane="2" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                    <SPLIT distance="200" swimtime="00:02:31.41" />
                    <SPLIT distance="250" swimtime="00:03:11.57" />
                    <SPLIT distance="300" swimtime="00:03:51.84" />
                    <SPLIT distance="350" swimtime="00:04:32.20" />
                    <SPLIT distance="400" swimtime="00:05:12.76" />
                    <SPLIT distance="450" swimtime="00:05:53.26" />
                    <SPLIT distance="500" swimtime="00:06:34.08" />
                    <SPLIT distance="550" swimtime="00:07:14.44" />
                    <SPLIT distance="600" swimtime="00:07:55.34" />
                    <SPLIT distance="650" swimtime="00:08:36.26" />
                    <SPLIT distance="700" swimtime="00:09:16.59" />
                    <SPLIT distance="750" swimtime="00:09:55.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-12" firstname="Zuzana " gender="F" lastname="Matúšová" nation="SVK" athleteid="9058">
              <RESULTS>
                <RESULT eventid="1058" points="695" reactiontime="+89" swimtime="00:00:30.07" resultid="9059" heatid="14141" lane="0" entrytime="00:00:29.80" />
                <RESULT eventid="8261" points="692" reactiontime="+79" swimtime="00:01:05.33" resultid="9060" heatid="14222" lane="4" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="723" reactiontime="+83" swimtime="00:00:32.75" resultid="9061" heatid="14289" lane="2" entrytime="00:00:31.10" />
                <RESULT eventid="8196" points="615" reactiontime="+77" swimtime="00:00:37.47" resultid="9062" heatid="14196" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="8678" points="787" reactiontime="+76" swimtime="00:00:36.70" resultid="9063" heatid="14377" lane="3" entrytime="00:00:37.50" />
                <RESULT eventid="8293" points="769" reactiontime="+84" swimtime="00:01:13.92" resultid="9064" heatid="14242" lane="4" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="728" reactiontime="+90" swimtime="00:02:41.47" resultid="9065" heatid="14165" lane="0" entrytime="00:02:42.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:02:03.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+104" swimtime="00:02:06.91" resultid="9070" heatid="14175" lane="4" entrytime="00:02:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:38.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8861" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="9042" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="9058" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="9050" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+87" swimtime="00:02:19.12" resultid="9113" heatid="14391" lane="9" entrytime="00:02:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="150" swimtime="00:01:48.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9050" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="9042" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="9058" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="8861" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9131" name="Legia Warszawa">
          <CONTACT city="Warszawa" email="twilczega@gmail.com" name="Tomasz Wilczęga" phone="+48531984974" />
          <ATHLETES>
            <ATHLETE birthdate="1976-11-12" firstname="Marcin" gender="M" lastname="Podhorecki" nation="POL" athleteid="9183">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9184" heatid="14147" lane="0" entrytime="00:00:34.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-21" firstname="Piotr" gender="M" lastname="Ciałkowski" nation="POL" athleteid="9181" />
            <ATHLETE birthdate="1966-08-13" firstname="Roman" gender="M" lastname="Kozłowski" nation="POL" athleteid="9948">
              <RESULTS>
                <RESULT eventid="1075" points="736" reactiontime="+84" swimtime="00:00:28.14" resultid="9949" heatid="14151" lane="2" entrytime="00:00:29.51" />
                <RESULT eventid="8309" points="810" reactiontime="+75" swimtime="00:01:09.87" resultid="9950" heatid="14250" lane="5" entrytime="00:01:13.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="822" reactiontime="+88" swimtime="00:01:14.24" resultid="9951" heatid="14280" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="710" reactiontime="+88" swimtime="00:00:30.68" resultid="9952" heatid="14296" lane="0" entrytime="00:00:31.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-09" firstname="Jakub" gender="M" lastname="Dobies" nation="POL" athleteid="9177">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9178" heatid="14147" lane="9" entrytime="00:00:34.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-02" firstname="Władysław" gender="M" lastname="Surała" nation="POL" athleteid="9182" />
            <ATHLETE birthdate="1976-01-04" firstname="Hubert" gender="M" lastname="Markowski" nation="POL" athleteid="9160">
              <RESULTS>
                <RESULT eventid="1105" points="546" reactiontime="+91" swimtime="00:02:36.42" resultid="9161" heatid="14171" lane="3" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="485" reactiontime="+76" swimtime="00:00:34.55" resultid="9162" heatid="14204" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="8341" points="532" reactiontime="+87" swimtime="00:02:35.49" resultid="9163" heatid="14261" lane="7" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:55.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="9164" heatid="14313" lane="9" entrytime="00:01:14.00" />
                <RESULT eventid="8582" points="478" reactiontime="+92" swimtime="00:05:46.59" resultid="9165" heatid="14347" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:17.91" />
                    <SPLIT distance="150" swimtime="00:02:03.53" />
                    <SPLIT distance="200" swimtime="00:02:47.13" />
                    <SPLIT distance="250" swimtime="00:03:37.14" />
                    <SPLIT distance="300" swimtime="00:04:26.85" />
                    <SPLIT distance="350" swimtime="00:05:08.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="598" reactiontime="+86" swimtime="00:01:07.20" resultid="9166" heatid="14358" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="558" reactiontime="+61" swimtime="00:02:38.44" resultid="9167" heatid="14369" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:01:59.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="9144">
              <RESULTS>
                <RESULT eventid="1075" points="758" reactiontime="+76" swimtime="00:00:25.05" resultid="9145" heatid="14159" lane="3" entrytime="00:00:25.10" />
                <RESULT eventid="8309" points="761" reactiontime="+76" swimtime="00:01:00.45" resultid="9146" heatid="14255" lane="1" entrytime="00:00:59.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="909" reactiontime="+76" swimtime="00:01:04.02" resultid="9147" heatid="14284" lane="2" entrytime="00:01:04.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="671" swimtime="00:00:27.07" resultid="9148" heatid="14302" lane="9" entrytime="00:00:25.99" />
                <RESULT eventid="8694" points="941" reactiontime="+68" swimtime="00:00:28.83" resultid="9149" heatid="14389" lane="6" entrytime="00:00:28.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-16" firstname="Jacek" gender="M" lastname="Kaczyński" nation="POL" athleteid="9141">
              <RESULTS>
                <RESULT eventid="1075" points="769" reactiontime="+82" swimtime="00:00:24.15" resultid="9142" heatid="14160" lane="4" entrytime="00:00:24.00" />
                <RESULT eventid="8454" points="692" swimtime="00:00:25.85" resultid="9143" heatid="14302" lane="8" entrytime="00:00:25.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-05" firstname="Karolina" gender="F" lastname="Modzelan" nation="POL" athleteid="9199">
              <RESULTS>
                <RESULT eventid="1058" points="632" reactiontime="+74" swimtime="00:00:30.45" resultid="9200" heatid="14140" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="8229" status="DNS" swimtime="00:00:00.00" resultid="9201" heatid="14211" lane="1" entrytime="00:03:10.00" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="9202" heatid="14222" lane="5" entrytime="00:01:09.00" />
                <RESULT eventid="8293" status="DNS" swimtime="00:00:00.00" resultid="9203" heatid="14242" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="9204" heatid="14273" lane="6" entrytime="00:01:28.00" />
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="9205" heatid="14376" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-23" firstname="Katarzyna" gender="F" lastname="Żołnowska" nation="POL" athleteid="9192">
              <RESULTS>
                <RESULT eventid="1090" points="977" reactiontime="+81" swimtime="00:02:24.24" resultid="9193" heatid="14165" lane="5" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="984" reactiontime="+83" swimtime="00:17:59.31" resultid="9194" heatid="14187" lane="5" entrytime="00:19:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                    <SPLIT distance="150" swimtime="00:01:42.16" />
                    <SPLIT distance="200" swimtime="00:02:17.51" />
                    <SPLIT distance="250" swimtime="00:02:53.33" />
                    <SPLIT distance="300" swimtime="00:03:29.48" />
                    <SPLIT distance="350" swimtime="00:04:05.69" />
                    <SPLIT distance="400" swimtime="00:04:42.20" />
                    <SPLIT distance="450" swimtime="00:05:18.19" />
                    <SPLIT distance="500" swimtime="00:05:54.32" />
                    <SPLIT distance="550" swimtime="00:06:30.38" />
                    <SPLIT distance="600" swimtime="00:07:06.43" />
                    <SPLIT distance="650" swimtime="00:07:42.37" />
                    <SPLIT distance="700" swimtime="00:08:18.67" />
                    <SPLIT distance="750" swimtime="00:08:54.90" />
                    <SPLIT distance="800" swimtime="00:09:31.23" />
                    <SPLIT distance="850" swimtime="00:10:07.71" />
                    <SPLIT distance="900" swimtime="00:10:44.20" />
                    <SPLIT distance="950" swimtime="00:11:20.36" />
                    <SPLIT distance="1000" swimtime="00:11:56.73" />
                    <SPLIT distance="1050" swimtime="00:12:33.31" />
                    <SPLIT distance="1100" swimtime="00:13:09.25" />
                    <SPLIT distance="1150" swimtime="00:13:45.71" />
                    <SPLIT distance="1200" swimtime="00:14:21.96" />
                    <SPLIT distance="1250" swimtime="00:14:58.68" />
                    <SPLIT distance="1300" swimtime="00:15:35.47" />
                    <SPLIT distance="1350" swimtime="00:16:12.04" />
                    <SPLIT distance="1400" swimtime="00:16:48.70" />
                    <SPLIT distance="1450" swimtime="00:17:25.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="819" reactiontime="+86" swimtime="00:00:31.68" resultid="9195" heatid="14197" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="8261" points="810" reactiontime="+82" swimtime="00:01:00.18" resultid="9196" heatid="14223" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="907" reactiontime="+89" swimtime="00:02:09.16" resultid="9197" heatid="14321" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="150" swimtime="00:01:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="9198" heatid="14365" lane="4" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="9137">
              <RESULTS>
                <RESULT eventid="1075" points="710" reactiontime="+81" swimtime="00:00:25.77" resultid="9138" heatid="14156" lane="3" entrytime="00:00:26.62" />
                <RESULT eventid="8277" points="716" reactiontime="+74" swimtime="00:00:57.48" resultid="9139" heatid="14234" lane="6" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="601" reactiontime="+77" swimtime="00:00:29.48" resultid="9140" heatid="14299" lane="1" entrytime="00:00:28.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-25" firstname="Adrian" gender="M" lastname="Jagodziński" nation="POL" athleteid="9179">
              <RESULTS>
                <RESULT eventid="1075" points="441" reactiontime="+91" swimtime="00:00:29.07" resultid="9180" heatid="14151" lane="8" entrytime="00:00:29.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-08-19" firstname="Paweł" gender="M" lastname="Filipowski" nation="POL" athleteid="9185">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9186" heatid="14147" lane="1" entrytime="00:00:34.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="9154">
              <RESULTS>
                <RESULT eventid="1075" points="1008" reactiontime="+70" swimtime="00:00:23.69" resultid="9155" heatid="14160" lane="7" entrytime="00:00:24.63" />
                <RESULT comment="Rekord Polski, Rekord Europy" eventid="8213" points="1168" reactiontime="+71" swimtime="00:00:25.78" resultid="9156" heatid="14207" lane="5" entrytime="00:00:26.17" />
                <RESULT eventid="8454" points="1048" reactiontime="+72" swimtime="00:00:24.74" resultid="9157" heatid="14290" lane="5" />
                <RESULT comment="Rekord Polski" eventid="8486" points="1095" reactiontime="+80" swimtime="00:00:57.30" resultid="9158" heatid="14315" lane="5" entrytime="00:00:57.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9159" heatid="14361" lane="9" entrytime="00:00:59.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-22" firstname="Mariusz" gender="M" lastname="Mikołajewski" nation="POL" athleteid="9150">
              <RESULTS>
                <RESULT eventid="1075" points="834" reactiontime="+79" swimtime="00:00:24.26" resultid="9151" heatid="14160" lane="3" entrytime="00:00:24.00" />
                <RESULT eventid="8309" points="841" reactiontime="+82" swimtime="00:00:58.47" resultid="9152" heatid="14255" lane="2" entrytime="00:00:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="9153" heatid="14284" lane="9" entrytime="00:01:07.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-04" firstname="Marcin" gender="M" lastname="Walkowicz" nation="POL" athleteid="9187">
              <RESULTS>
                <RESULT eventid="1075" points="394" reactiontime="+72" swimtime="00:00:32.41" resultid="9188" heatid="14147" lane="8" entrytime="00:00:34.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-01" firstname="Stanisław" gender="M" lastname="Fluder" nation="POL" athleteid="9168">
              <RESULTS>
                <RESULT eventid="1075" points="545" reactiontime="+83" swimtime="00:00:27.09" resultid="9169" heatid="14158" lane="9" entrytime="00:00:26.15" />
                <RESULT eventid="1150" points="636" reactiontime="+90" swimtime="00:09:40.22" resultid="9170" heatid="14182" lane="8" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:46.76" />
                    <SPLIT distance="200" swimtime="00:02:23.80" />
                    <SPLIT distance="250" swimtime="00:03:01.20" />
                    <SPLIT distance="300" swimtime="00:03:38.47" />
                    <SPLIT distance="350" swimtime="00:04:15.22" />
                    <SPLIT distance="400" swimtime="00:04:51.83" />
                    <SPLIT distance="450" swimtime="00:05:28.65" />
                    <SPLIT distance="500" swimtime="00:06:05.40" />
                    <SPLIT distance="550" swimtime="00:06:42.11" />
                    <SPLIT distance="600" swimtime="00:07:18.27" />
                    <SPLIT distance="650" swimtime="00:07:54.46" />
                    <SPLIT distance="700" swimtime="00:08:30.51" />
                    <SPLIT distance="750" swimtime="00:09:06.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="542" reactiontime="+83" swimtime="00:00:32.49" resultid="9171" heatid="14205" lane="4" entrytime="00:00:31.20" />
                <RESULT eventid="8277" points="593" reactiontime="+85" swimtime="00:00:58.35" resultid="9172" heatid="14236" lane="2" entrytime="00:00:56.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="459" reactiontime="+87" swimtime="00:00:29.63" resultid="9173" heatid="14300" lane="0" entrytime="00:00:28.10" />
                <RESULT eventid="8518" points="578" reactiontime="+80" swimtime="00:02:07.87" resultid="9174" heatid="14332" lane="7" entrytime="00:02:07.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="9206">
              <RESULTS>
                <RESULT eventid="1058" points="723" reactiontime="+88" swimtime="00:00:29.12" resultid="9207" heatid="14141" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1090" points="779" reactiontime="+85" swimtime="00:02:35.42" resultid="9208" heatid="14165" lane="6" entrytime="00:02:32.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="838" reactiontime="+125" swimtime="00:00:32.20" resultid="9209" heatid="14197" lane="5" entrytime="00:00:31.90" />
                <RESULT eventid="8293" points="757" reactiontime="+91" swimtime="00:01:11.13" resultid="9210" heatid="14243" lane="2" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="854" reactiontime="+87" swimtime="00:01:10.11" resultid="9211" heatid="14307" lane="3" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="9212" heatid="14342" lane="2" entrytime="00:05:35.00" />
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="9213" heatid="14365" lane="3" entrytime="00:02:32.00" />
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="9214" heatid="14377" lane="5" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-15" firstname="Aleksandra" gender="F" lastname="Marianek" nation="POL" athleteid="9189">
              <RESULTS>
                <RESULT eventid="8229" points="470" reactiontime="+86" swimtime="00:03:17.57" resultid="9190" heatid="14210" lane="5" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:01:34.05" />
                    <SPLIT distance="150" swimtime="00:02:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="9191" heatid="14272" lane="5" entrytime="00:01:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Patryk" gender="M" lastname="Wakuła" nation="POL" athleteid="9175">
              <RESULTS>
                <RESULT eventid="1075" points="650" reactiontime="+73" swimtime="00:00:25.54" resultid="9176" heatid="14159" lane="7" entrytime="00:00:25.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-26" firstname="Tomasz" gender="M" lastname="Wilczęga" nation="POL" athleteid="9132">
              <RESULTS>
                <RESULT eventid="1075" points="688" reactiontime="+79" swimtime="00:00:25.06" resultid="9133" heatid="14159" lane="2" entrytime="00:00:25.39" />
                <RESULT eventid="8277" points="696" reactiontime="+77" swimtime="00:00:55.32" resultid="9134" heatid="14224" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="546" reactiontime="+79" swimtime="00:01:07.29" resultid="9135" heatid="14253" lane="2" entrytime="00:01:06.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="584" reactiontime="+80" swimtime="00:00:27.36" resultid="9136" heatid="14300" lane="2" entrytime="00:00:27.69" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+74" swimtime="00:01:38.58" resultid="9217" heatid="14339" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="150" swimtime="00:01:15.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9132" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="9175" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="9144" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="9150" number="4" reactiontime="+7" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+72" swimtime="00:01:37.98" resultid="9218" heatid="14339" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                    <SPLIT distance="100" swimtime="00:00:50.25" />
                    <SPLIT distance="150" swimtime="00:01:15.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9154" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9168" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="9137" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="9141" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8550" status="DSQ" swimtime="00:02:18.95" resultid="9219" heatid="14337" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="150" swimtime="00:01:29.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9179" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="9182" number="2" reactiontime="+87" status="DSQ" />
                    <RELAYPOSITION athleteid="9177" number="3" reactiontime="-5" status="DSQ" />
                    <RELAYPOSITION athleteid="9181" number="4" reactiontime="+57" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+72" swimtime="00:02:22.48" resultid="9220" heatid="14266" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:26.91" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9177" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="9181" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="9175" number="3" reactiontime="+87" />
                    <RELAYPOSITION athleteid="9179" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT comment="Rekord Europy, Rekord Polski, pierwsza zmiana, kat.40-44" eventid="8373" reactiontime="+66" swimtime="00:01:55.01" resultid="9221" heatid="14268" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.54" />
                    <SPLIT distance="100" swimtime="00:00:57.61" />
                    <SPLIT distance="150" swimtime="00:01:27.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9154" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="9137" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="9160" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="9168" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+68" swimtime="00:01:46.23" resultid="9222" heatid="14268" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="100" swimtime="00:00:56.37" />
                    <SPLIT distance="150" swimtime="00:01:21.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9150" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="9144" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="9141" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="9132" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="9">
              <RESULTS>
                <RESULT eventid="8534" status="DNS" swimtime="00:00:00.00" resultid="9223" heatid="14335" lane="5" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9206" number="1" />
                    <RELAYPOSITION athleteid="9189" number="2" />
                    <RELAYPOSITION athleteid="9199" number="3" />
                    <RELAYPOSITION athleteid="9192" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="10">
              <RESULTS>
                <RESULT comment="Rekord Polski , pierwsza zmiana" eventid="8357" reactiontime="+76" swimtime="00:02:26.00" resultid="9224" heatid="14264" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:01:53.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9206" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="9189" number="2" reactiontime="+123" />
                    <RELAYPOSITION athleteid="9192" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="9199" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="9215" heatid="14176" lane="2" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9144" number="1" />
                    <RELAYPOSITION athleteid="9199" number="2" />
                    <RELAYPOSITION athleteid="9150" number="3" />
                    <RELAYPOSITION athleteid="9189" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+90" swimtime="00:01:43.14" resultid="9216" heatid="14176" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="100" swimtime="00:00:56.45" />
                    <SPLIT distance="150" swimtime="00:01:19.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9141" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="9192" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="9206" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="9154" number="4" reactiontime="-3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="11">
              <RESULTS>
                <RESULT eventid="8710" status="DNS" swimtime="00:00:00.00" resultid="9225" heatid="14392" lane="2" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9154" number="1" />
                    <RELAYPOSITION athleteid="9144" number="2" />
                    <RELAYPOSITION athleteid="9206" number="3" />
                    <RELAYPOSITION athleteid="9192" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9458" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="DM" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="9459">
              <RESULTS>
                <RESULT eventid="1165" points="740" reactiontime="+90" swimtime="00:20:29.41" resultid="9460" heatid="14187" lane="3" entrytime="00:19:46.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:12.99" />
                    <SPLIT distance="150" swimtime="00:01:52.46" />
                    <SPLIT distance="200" swimtime="00:02:32.35" />
                    <SPLIT distance="250" swimtime="00:03:12.13" />
                    <SPLIT distance="300" swimtime="00:03:52.20" />
                    <SPLIT distance="350" swimtime="00:04:32.45" />
                    <SPLIT distance="400" swimtime="00:05:12.91" />
                    <SPLIT distance="450" swimtime="00:05:53.12" />
                    <SPLIT distance="500" swimtime="00:06:33.74" />
                    <SPLIT distance="550" swimtime="00:07:14.38" />
                    <SPLIT distance="600" swimtime="00:07:55.05" />
                    <SPLIT distance="650" swimtime="00:08:36.08" />
                    <SPLIT distance="700" swimtime="00:09:17.30" />
                    <SPLIT distance="750" swimtime="00:09:58.80" />
                    <SPLIT distance="800" swimtime="00:10:40.23" />
                    <SPLIT distance="850" swimtime="00:11:22.18" />
                    <SPLIT distance="900" swimtime="00:12:04.11" />
                    <SPLIT distance="950" swimtime="00:12:45.77" />
                    <SPLIT distance="1000" swimtime="00:13:28.13" />
                    <SPLIT distance="1050" swimtime="00:14:10.11" />
                    <SPLIT distance="1100" swimtime="00:14:52.77" />
                    <SPLIT distance="1150" swimtime="00:15:34.85" />
                    <SPLIT distance="1200" swimtime="00:16:17.36" />
                    <SPLIT distance="1250" swimtime="00:16:59.69" />
                    <SPLIT distance="1300" swimtime="00:17:42.58" />
                    <SPLIT distance="1350" swimtime="00:18:24.90" />
                    <SPLIT distance="1400" swimtime="00:19:06.75" />
                    <SPLIT distance="1450" swimtime="00:19:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="694" reactiontime="+77" swimtime="00:01:05.25" resultid="9461" heatid="14223" lane="8" entrytime="00:01:05.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="729" reactiontime="+89" swimtime="00:02:22.32" resultid="9462" heatid="14321" lane="7" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="735" reactiontime="+86" swimtime="00:05:02.61" resultid="9463" heatid="14393" lane="6" entrytime="00:04:56.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                    <SPLIT distance="150" swimtime="00:01:51.58" />
                    <SPLIT distance="200" swimtime="00:02:30.30" />
                    <SPLIT distance="250" swimtime="00:03:09.47" />
                    <SPLIT distance="300" swimtime="00:03:48.17" />
                    <SPLIT distance="350" swimtime="00:04:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="9464">
              <RESULTS>
                <RESULT eventid="1105" points="411" reactiontime="+97" swimtime="00:03:11.40" resultid="9465" heatid="14169" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:27.12" />
                    <SPLIT distance="150" swimtime="00:02:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="428" reactiontime="+95" swimtime="00:03:25.32" resultid="9466" heatid="14214" lane="8" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:36.19" />
                    <SPLIT distance="150" swimtime="00:02:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8341" reactiontime="+71" status="DSQ" swimtime="00:03:41.97" resultid="9467" heatid="14259" lane="3" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:45.61" />
                    <SPLIT distance="150" swimtime="00:02:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="9468" heatid="14278" lane="7" entrytime="00:01:33.00" />
                <RESULT eventid="8582" points="365" reactiontime="+115" swimtime="00:07:11.30" resultid="9469" heatid="14345" lane="2" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:45.61" />
                    <SPLIT distance="150" swimtime="00:02:39.95" />
                    <SPLIT distance="200" swimtime="00:03:33.55" />
                    <SPLIT distance="250" swimtime="00:04:33.00" />
                    <SPLIT distance="300" swimtime="00:05:34.23" />
                    <SPLIT distance="350" swimtime="00:06:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="384" reactiontime="+92" swimtime="00:03:11.30" resultid="9470" heatid="14369" lane="9" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:30.81" />
                    <SPLIT distance="150" swimtime="00:02:21.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="9471" heatid="14383" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="RZ" clubid="10236" name="Masters Ikar Mielec">
          <CONTACT city="MIELEC" email="sebastianboicetta@gmail.com" name="SEBASTIAN BOICETTA" phone="501072284" state="PODKA" street="WARSZAWSKA 6/41" zip="39-300" />
          <ATHLETES>
            <ATHLETE birthdate="1988-06-09" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" license="503208700002" athleteid="10237">
              <RESULTS>
                <RESULT eventid="8179" points="631" reactiontime="+84" swimtime="00:19:18.12" resultid="10238" heatid="14189" lane="5" entrytime="00:17:52.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:43.76" />
                    <SPLIT distance="200" swimtime="00:02:20.73" />
                    <SPLIT distance="250" swimtime="00:02:58.51" />
                    <SPLIT distance="300" swimtime="00:03:36.46" />
                    <SPLIT distance="350" swimtime="00:04:15.02" />
                    <SPLIT distance="400" swimtime="00:04:53.97" />
                    <SPLIT distance="450" swimtime="00:05:33.03" />
                    <SPLIT distance="500" swimtime="00:06:11.82" />
                    <SPLIT distance="550" swimtime="00:06:51.95" />
                    <SPLIT distance="600" swimtime="00:07:31.28" />
                    <SPLIT distance="650" swimtime="00:08:10.40" />
                    <SPLIT distance="700" swimtime="00:08:49.59" />
                    <SPLIT distance="750" swimtime="00:09:29.34" />
                    <SPLIT distance="800" swimtime="00:10:09.07" />
                    <SPLIT distance="850" swimtime="00:10:48.80" />
                    <SPLIT distance="900" swimtime="00:11:28.42" />
                    <SPLIT distance="950" swimtime="00:12:07.96" />
                    <SPLIT distance="1000" swimtime="00:12:47.61" />
                    <SPLIT distance="1050" swimtime="00:13:27.10" />
                    <SPLIT distance="1100" swimtime="00:14:06.76" />
                    <SPLIT distance="1150" swimtime="00:14:46.32" />
                    <SPLIT distance="1200" swimtime="00:15:25.47" />
                    <SPLIT distance="1250" swimtime="00:16:05.59" />
                    <SPLIT distance="1300" swimtime="00:16:44.97" />
                    <SPLIT distance="1350" swimtime="00:17:23.36" />
                    <SPLIT distance="1400" swimtime="00:18:01.41" />
                    <SPLIT distance="1450" swimtime="00:18:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="10239" heatid="14262" lane="5" entrytime="00:02:14.24" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASKRAS" nation="POL" region="LBL" clubid="9390" name="Masters Kraśnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.com" name="Michalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 1" zip="23-204" />
          <ATHLETES>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="9403">
              <RESULTS>
                <RESULT eventid="1105" points="297" reactiontime="+94" swimtime="00:03:54.36" resultid="9404" heatid="14168" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="100" swimtime="00:01:53.98" />
                    <SPLIT distance="150" swimtime="00:03:03.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="314" reactiontime="+94" swimtime="00:00:46.74" resultid="9405" heatid="14200" lane="2" entrytime="00:00:51.00" />
                <RESULT eventid="8486" points="339" reactiontime="+99" swimtime="00:01:43.46" resultid="9406" heatid="14310" lane="7" entrytime="00:01:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="312" reactiontime="+125" swimtime="00:08:20.53" resultid="9407" heatid="14344" lane="2" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.20" />
                    <SPLIT distance="100" swimtime="00:02:04.31" />
                    <SPLIT distance="150" swimtime="00:03:10.43" />
                    <SPLIT distance="200" swimtime="00:04:11.80" />
                    <SPLIT distance="250" swimtime="00:05:23.65" />
                    <SPLIT distance="300" swimtime="00:06:34.08" />
                    <SPLIT distance="350" swimtime="00:07:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9408" heatid="14354" lane="5" entrytime="00:01:50.35" />
                <RESULT eventid="8662" points="353" reactiontime="+87" swimtime="00:03:44.36" resultid="9409" heatid="14367" lane="5" entrytime="00:04:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.37" />
                    <SPLIT distance="100" swimtime="00:01:49.93" />
                    <SPLIT distance="150" swimtime="00:02:49.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-04" firstname="Zdzisław" gender="M" lastname="Bąk" nation="POL" athleteid="9398">
              <RESULTS>
                <RESULT eventid="1075" points="485" reactiontime="+77" swimtime="00:00:33.19" resultid="9399" heatid="14147" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="8277" points="460" reactiontime="+101" swimtime="00:01:15.16" resultid="9400" heatid="14226" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="462" reactiontime="+139" swimtime="00:02:49.49" resultid="9401" heatid="14325" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="480" reactiontime="+88" swimtime="00:06:01.99" resultid="9402" heatid="14402" lane="7" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:02:06.38" />
                    <SPLIT distance="200" swimtime="00:02:53.38" />
                    <SPLIT distance="250" swimtime="00:03:41.04" />
                    <SPLIT distance="300" swimtime="00:04:29.18" />
                    <SPLIT distance="350" swimtime="00:05:17.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-17" firstname="Jacek" gender="M" lastname="Janik" nation="POL" athleteid="9391">
              <RESULTS>
                <RESULT eventid="1075" points="331" reactiontime="+94" swimtime="00:00:36.72" resultid="9392" heatid="14146" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="8245" points="317" reactiontime="+129" swimtime="00:03:46.94" resultid="9393" heatid="14213" lane="0" entrytime="00:03:50.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.08" />
                    <SPLIT distance="100" swimtime="00:01:46.87" />
                    <SPLIT distance="150" swimtime="00:02:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="292" reactiontime="+110" swimtime="00:01:25.04" resultid="9394" heatid="14226" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="346" reactiontime="+92" swimtime="00:01:39.02" resultid="9395" heatid="14277" lane="8" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="260" reactiontime="+114" swimtime="00:03:14.92" resultid="9396" heatid="14324" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:01:31.15" />
                    <SPLIT distance="150" swimtime="00:02:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="316" reactiontime="+96" swimtime="00:00:45.14" resultid="9397" heatid="14381" lane="6" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="9410">
              <RESULTS>
                <RESULT eventid="1075" points="258" reactiontime="+99" swimtime="00:00:42.16" resultid="9411" heatid="14143" lane="3" entrytime="00:00:50.28" />
                <RESULT eventid="8213" points="184" reactiontime="+96" swimtime="00:00:55.88" resultid="9412" heatid="14199" lane="4" entrytime="00:00:58.32" />
                <RESULT eventid="8309" points="267" reactiontime="+99" swimtime="00:01:49.99" resultid="9413" heatid="14245" lane="5" entrytime="00:01:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="189" reactiontime="+96" swimtime="00:00:50.78" resultid="9414" heatid="14291" lane="8" entrytime="00:00:59.20" />
                <RESULT eventid="8630" points="130" reactiontime="+99" swimtime="00:02:12.79" resultid="9415" heatid="14354" lane="0" entrytime="00:02:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBL" clubid="9255" name="Masters Lublin">
          <CONTACT city="LUBLIN" email="masters_lublin@wp.pl" name="WÓJCICKI" phone="+48501794954" state="LUB" street="STANISŁAWA LEMA 18" zip="20-445" />
          <ATHLETES>
            <ATHLETE birthdate="1975-11-07" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" license="103503700005" athleteid="9256">
              <RESULTS>
                <RESULT eventid="8309" points="517" reactiontime="+84" swimtime="00:01:14.50" resultid="9257" heatid="14249" lane="6" entrytime="00:01:15.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="399" reactiontime="+98" swimtime="00:02:33.50" resultid="9258" heatid="14327" lane="3" entrytime="00:02:35.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:12.96" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="346" reactiontime="+99" swimtime="00:05:42.59" resultid="9259" heatid="14401" lane="9" entrytime="00:05:40.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:02:01.76" />
                    <SPLIT distance="200" swimtime="00:02:45.78" />
                    <SPLIT distance="250" swimtime="00:03:30.02" />
                    <SPLIT distance="300" swimtime="00:04:15.96" />
                    <SPLIT distance="350" swimtime="00:05:00.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-10-21" firstname="Adam" gender="M" lastname="Pietrzak" nation="POL" license="103503700011" athleteid="9271">
              <RESULTS>
                <RESULT eventid="1075" points="357" reactiontime="+100" swimtime="00:00:31.17" resultid="9272" heatid="14149" lane="5" entrytime="00:00:30.38" entrycourse="SCM" />
                <RESULT eventid="8213" points="374" reactiontime="+79" swimtime="00:00:36.75" resultid="9273" heatid="14203" lane="7" entrytime="00:00:35.87" entrycourse="SCM" />
                <RESULT eventid="8309" points="348" reactiontime="+97" swimtime="00:01:18.17" resultid="9274" heatid="14249" lane="3" entrytime="00:01:15.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="393" reactiontime="+96" swimtime="00:01:23.72" resultid="9275" heatid="14281" lane="2" entrytime="00:01:20.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="357" reactiontime="+91" swimtime="00:01:21.12" resultid="9276" heatid="14312" lane="9" entrytime="00:01:20.72" entrycourse="SCM" />
                <RESULT eventid="8662" points="304" reactiontime="+84" swimtime="00:02:53.35" resultid="9277" heatid="14370" lane="3" entrytime="00:02:30.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:01:25.97" />
                    <SPLIT distance="150" swimtime="00:02:09.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="382" reactiontime="+82" swimtime="00:00:38.30" resultid="9278" heatid="14384" lane="1" entrytime="00:00:38.11" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-28" firstname="Rafał" gender="M" lastname="Wójcicki" nation="POL" license="103503700001" athleteid="9267">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9268" heatid="14153" lane="2" entrytime="00:00:28.35" entrycourse="SCM" />
                <RESULT eventid="8213" points="361" reactiontime="+70" swimtime="00:00:38.11" resultid="9269" heatid="14203" lane="9" entrytime="00:00:36.81" entrycourse="SCM" />
                <RESULT eventid="8486" points="377" reactiontime="+83" swimtime="00:01:21.71" resultid="9270" heatid="14312" lane="3" entrytime="00:01:17.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-06" firstname="Marek" gender="M" lastname="Walencik" nation="POL" license="103503700010" athleteid="9279">
              <RESULTS>
                <RESULT eventid="8213" points="629" reactiontime="+88" swimtime="00:00:31.68" resultid="9280" heatid="14204" lane="4" entrytime="00:00:32.82" entrycourse="SCM" />
                <RESULT eventid="8309" points="655" reactiontime="+93" swimtime="00:01:08.88" resultid="9281" heatid="14249" lane="4" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="668" reactiontime="+88" swimtime="00:01:15.06" resultid="9282" heatid="14282" lane="2" entrytime="00:01:17.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="577" reactiontime="+104" swimtime="00:01:10.94" resultid="9283" heatid="14313" lane="8" entrytime="00:01:12.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="699" reactiontime="+75" swimtime="00:00:33.22" resultid="9284" heatid="14387" lane="6" entrytime="00:00:34.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-28" firstname="Anna" gender="F" lastname="Michalska" nation="POL" license="103503600002" athleteid="9260">
              <RESULTS>
                <RESULT eventid="1090" points="522" reactiontime="+103" swimtime="00:03:02.32" resultid="9261" heatid="14164" lane="8" entrytime="00:03:10.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                    <SPLIT distance="150" swimtime="00:02:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="554" reactiontime="+99" swimtime="00:00:37.19" resultid="9262" heatid="14196" lane="0" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="8293" points="591" reactiontime="+84" swimtime="00:01:21.18" resultid="9263" heatid="14241" lane="8" entrytime="00:01:26.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="596" reactiontime="+87" swimtime="00:01:20.72" resultid="9264" heatid="14306" lane="3" entrytime="00:01:22.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="588" reactiontime="+75" swimtime="00:02:58.25" resultid="9265" heatid="14364" lane="4" entrytime="00:03:07.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="524" reactiontime="+105" swimtime="00:00:42.59" resultid="9266" heatid="14376" lane="7" entrytime="00:00:40.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+80" swimtime="00:02:12.45" resultid="9285" heatid="14267" lane="9" entrytime="00:02:10.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:01:44.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9279" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="9271" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="9267" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="9256" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+88" swimtime="00:01:57.63" resultid="9286" heatid="14338" lane="7" entrytime="00:01:52.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:28.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9279" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="9271" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="9267" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="9256" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12385" name="Masters Rzeszów">
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="12386">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="12387" heatid="14148" lane="7" entrytime="00:00:32.20" />
                <RESULT eventid="8179" points="516" reactiontime="+104" swimtime="00:24:25.05" resultid="12388" heatid="14191" lane="4" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:27.24" />
                    <SPLIT distance="150" swimtime="00:02:14.62" />
                    <SPLIT distance="200" swimtime="00:03:02.43" />
                    <SPLIT distance="250" swimtime="00:08:43.48" />
                    <SPLIT distance="300" swimtime="00:09:32.58" />
                    <SPLIT distance="350" swimtime="00:10:21.48" />
                    <SPLIT distance="400" swimtime="00:11:11.90" />
                    <SPLIT distance="450" swimtime="00:12:01.58" />
                    <SPLIT distance="500" swimtime="00:14:28.47" />
                    <SPLIT distance="550" swimtime="00:16:07.79" />
                    <SPLIT distance="600" swimtime="00:17:46.65" />
                    <SPLIT distance="650" swimtime="00:18:36.89" />
                    <SPLIT distance="700" swimtime="00:19:26.45" />
                    <SPLIT distance="750" swimtime="00:21:10.75" />
                    <SPLIT distance="800" swimtime="00:22:00.70" />
                    <SPLIT distance="1250" swimtime="00:23:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="513" reactiontime="+83" swimtime="00:01:14.76" resultid="12389" heatid="14228" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="12390" heatid="14247" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="8454" points="353" reactiontime="+97" swimtime="00:00:41.21" resultid="12391" heatid="14293" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="8518" points="540" reactiontime="+100" swimtime="00:02:47.56" resultid="12392" heatid="14326" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:06.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="525" reactiontime="+105" swimtime="00:06:05.70" resultid="12393" heatid="14402" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:12.98" />
                    <SPLIT distance="200" swimtime="00:03:00.70" />
                    <SPLIT distance="250" swimtime="00:03:47.62" />
                    <SPLIT distance="300" swimtime="00:04:34.21" />
                    <SPLIT distance="350" swimtime="00:05:21.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="9303" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="9327">
              <RESULTS>
                <RESULT eventid="1058" points="263" reactiontime="+121" swimtime="00:00:48.34" resultid="9328" heatid="14135" lane="5" entrytime="00:00:48.00" entrycourse="SCM" />
                <RESULT eventid="1090" points="261" reactiontime="+115" swimtime="00:04:36.11" resultid="9329" heatid="14162" lane="5" entrytime="00:04:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.15" />
                    <SPLIT distance="100" swimtime="00:02:14.80" />
                    <SPLIT distance="150" swimtime="00:03:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="305" reactiontime="+95" swimtime="00:00:57.18" resultid="9330" heatid="14193" lane="3" entrytime="00:00:57.30" entrycourse="SCM" />
                <RESULT eventid="8261" points="294" reactiontime="+103" swimtime="00:01:47.36" resultid="9331" heatid="14219" lane="9" entrytime="00:01:48.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="282" reactiontime="+82" swimtime="00:02:07.81" resultid="9332" heatid="14304" lane="6" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="286" reactiontime="+126" swimtime="00:04:00.92" resultid="9333" heatid="14317" lane="2" entrytime="00:04:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:01:54.77" />
                    <SPLIT distance="150" swimtime="00:03:00.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="191" reactiontime="+96" swimtime="00:02:21.30" resultid="9334" heatid="14349" lane="4" entrytime="00:02:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="279" reactiontime="+89" swimtime="00:04:39.92" resultid="9335" heatid="14363" lane="9" entrytime="00:04:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.55" />
                    <SPLIT distance="100" swimtime="00:02:14.58" />
                    <SPLIT distance="150" swimtime="00:03:29.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="9345">
              <RESULTS>
                <RESULT eventid="8277" points="467" reactiontime="+84" swimtime="00:01:08.18" resultid="9346" heatid="14230" lane="1" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="521" reactiontime="+70" swimtime="00:00:32.85" resultid="9347" heatid="14295" lane="9" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="8518" points="370" reactiontime="+112" swimtime="00:02:39.80" resultid="9348" heatid="14327" lane="2" entrytime="00:02:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="351" reactiontime="+74" swimtime="00:01:23.31" resultid="9349" heatid="14356" lane="2" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="9304">
              <RESULTS>
                <RESULT eventid="1075" points="526" reactiontime="+119" swimtime="00:00:48.07" resultid="9305" heatid="14143" lane="6" entrytime="00:00:51.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="465" reactiontime="+136" swimtime="00:05:03.54" resultid="9306" heatid="14167" lane="1" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.10" />
                    <SPLIT distance="100" swimtime="00:02:38.39" />
                    <SPLIT distance="150" swimtime="00:04:01.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="446" reactiontime="+102" swimtime="00:01:01.70" resultid="9307" heatid="14199" lane="5" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="457" reactiontime="+123" swimtime="00:01:53.02" resultid="9308" heatid="14225" lane="9" entrytime="00:01:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="354" reactiontime="+124" swimtime="00:02:26.57" resultid="9309" heatid="14276" lane="6" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="487" reactiontime="+117" swimtime="00:04:07.35" resultid="9310" heatid="14323" lane="5" entrytime="00:04:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:57.49" />
                    <SPLIT distance="150" swimtime="00:03:02.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="421" reactiontime="+124" swimtime="00:01:03.37" resultid="9311" heatid="14380" lane="2" entrytime="00:01:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="9350">
              <RESULTS>
                <RESULT eventid="8277" points="168" reactiontime="+102" swimtime="00:01:50.57" resultid="9351" heatid="14224" lane="5" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="136" reactiontime="+128" swimtime="00:02:23.37" resultid="9352" heatid="14245" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="200" reactiontime="+79" swimtime="00:02:03.71" resultid="9353" heatid="14309" lane="5" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="183" reactiontime="+97" swimtime="00:04:11.20" resultid="9354" heatid="14323" lane="6" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.92" />
                    <SPLIT distance="100" swimtime="00:01:59.44" />
                    <SPLIT distance="150" swimtime="00:03:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="215" reactiontime="+79" swimtime="00:04:22.88" resultid="9355" heatid="14367" lane="7" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:03:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="173" reactiontime="+104" swimtime="00:09:11.15" resultid="9356" heatid="14404" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="100" swimtime="00:02:03.05" />
                    <SPLIT distance="150" swimtime="00:03:11.75" />
                    <SPLIT distance="200" swimtime="00:04:22.23" />
                    <SPLIT distance="250" swimtime="00:05:33.85" />
                    <SPLIT distance="300" swimtime="00:06:46.45" />
                    <SPLIT distance="350" swimtime="00:07:58.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="9318">
              <RESULTS>
                <RESULT eventid="1075" points="210" reactiontime="+95" swimtime="00:00:39.97" resultid="9319" heatid="14144" lane="7" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="128" reactiontime="+103" swimtime="00:04:13.47" resultid="9320" heatid="14167" lane="4" entrytime="00:04:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.57" />
                    <SPLIT distance="100" swimtime="00:02:01.66" />
                    <SPLIT distance="150" swimtime="00:03:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="125" reactiontime="+92" swimtime="00:00:54.17" resultid="9321" heatid="14200" lane="8" entrytime="00:00:55.00" entrycourse="SCM" />
                <RESULT eventid="8309" points="139" reactiontime="+106" swimtime="00:01:55.26" resultid="9322" heatid="14245" lane="4" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="155" reactiontime="+100" swimtime="00:02:02.05" resultid="9323" heatid="14276" lane="7" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="95" reactiontime="+93" swimtime="00:02:09.38" resultid="9324" heatid="14309" lane="6" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="73" reactiontime="+108" swimtime="00:02:15.27" resultid="9325" heatid="14354" lane="1" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="131" reactiontime="+96" swimtime="00:00:58.00" resultid="9326" heatid="14380" lane="5" entrytime="00:00:54.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" license="501806600049" athleteid="9336">
              <RESULTS>
                <RESULT eventid="1090" points="1005" reactiontime="+82" swimtime="00:02:22.91" resultid="9337" heatid="14165" lane="4" entrytime="00:02:21.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="799" reactiontime="+83" swimtime="00:19:17.17" resultid="9338" heatid="14187" lane="6" entrytime="00:20:35.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:08.23" />
                    <SPLIT distance="150" swimtime="00:01:44.04" />
                    <SPLIT distance="200" swimtime="00:02:20.67" />
                    <SPLIT distance="250" swimtime="00:02:58.27" />
                    <SPLIT distance="300" swimtime="00:03:36.07" />
                    <SPLIT distance="350" swimtime="00:04:14.16" />
                    <SPLIT distance="400" swimtime="00:04:52.65" />
                    <SPLIT distance="450" swimtime="00:05:31.55" />
                    <SPLIT distance="500" swimtime="00:06:10.65" />
                    <SPLIT distance="550" swimtime="00:06:49.28" />
                    <SPLIT distance="600" swimtime="00:07:28.02" />
                    <SPLIT distance="650" swimtime="00:08:06.83" />
                    <SPLIT distance="700" swimtime="00:08:45.75" />
                    <SPLIT distance="750" swimtime="00:09:24.71" />
                    <SPLIT distance="800" swimtime="00:10:03.71" />
                    <SPLIT distance="850" swimtime="00:10:43.36" />
                    <SPLIT distance="900" swimtime="00:11:22.89" />
                    <SPLIT distance="950" swimtime="00:12:02.40" />
                    <SPLIT distance="1000" swimtime="00:12:41.67" />
                    <SPLIT distance="1050" swimtime="00:13:21.23" />
                    <SPLIT distance="1100" swimtime="00:14:00.64" />
                    <SPLIT distance="1150" swimtime="00:14:40.16" />
                    <SPLIT distance="1200" swimtime="00:15:19.62" />
                    <SPLIT distance="1250" swimtime="00:15:59.43" />
                    <SPLIT distance="1300" swimtime="00:16:39.40" />
                    <SPLIT distance="1350" swimtime="00:17:18.81" />
                    <SPLIT distance="1400" swimtime="00:17:58.23" />
                    <SPLIT distance="1450" swimtime="00:18:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="848" reactiontime="+82" swimtime="00:00:59.28" resultid="9339" heatid="14223" lane="4" entrytime="00:00:58.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="909" reactiontime="+81" swimtime="00:01:07.36" resultid="9340" heatid="14243" lane="4" entrytime="00:01:07.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="905" reactiontime="+91" swimtime="00:02:09.27" resultid="9341" heatid="14321" lane="4" entrytime="00:02:06.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:01.97" />
                    <SPLIT distance="150" swimtime="00:01:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="908" reactiontime="+84" swimtime="00:05:10.01" resultid="9342" heatid="14342" lane="4" entrytime="00:04:59.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:11.09" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                    <SPLIT distance="200" swimtime="00:02:31.29" />
                    <SPLIT distance="250" swimtime="00:03:15.12" />
                    <SPLIT distance="300" swimtime="00:03:59.02" />
                    <SPLIT distance="350" swimtime="00:04:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="758" reactiontime="+75" swimtime="00:00:34.64" resultid="9343" heatid="14378" lane="4" entrytime="00:00:33.99" entrycourse="SCM" />
                <RESULT eventid="8726" points="851" reactiontime="+78" swimtime="00:04:42.64" resultid="9344" heatid="14393" lane="4" entrytime="00:04:31.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                    <SPLIT distance="150" swimtime="00:01:43.15" />
                    <SPLIT distance="200" swimtime="00:02:19.74" />
                    <SPLIT distance="250" swimtime="00:02:55.54" />
                    <SPLIT distance="300" swimtime="00:03:31.60" />
                    <SPLIT distance="350" swimtime="00:04:07.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-11" firstname="García Rodríguez" gender="M" lastname="Alberto" nation="POL" athleteid="9312">
              <RESULTS>
                <RESULT eventid="1075" points="563" reactiontime="+86" swimtime="00:00:26.80" resultid="9313" heatid="14158" lane="0" entrytime="00:00:26.11" entrycourse="SCM" />
                <RESULT eventid="1105" points="514" reactiontime="+81" swimtime="00:02:27.39" resultid="9314" heatid="14174" lane="8" entrytime="00:02:22.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="583" reactiontime="+80" swimtime="00:00:58.69" resultid="9315" heatid="14235" lane="6" entrytime="00:00:57.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="573" reactiontime="+86" swimtime="00:02:08.20" resultid="9316" heatid="14333" lane="2" entrytime="00:02:03.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:01.49" />
                    <SPLIT distance="150" swimtime="00:01:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="661" reactiontime="+80" swimtime="00:04:35.73" resultid="9317" heatid="14398" lane="6" entrytime="00:04:23.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:38.91" />
                    <SPLIT distance="200" swimtime="00:02:14.10" />
                    <SPLIT distance="250" swimtime="00:02:49.29" />
                    <SPLIT distance="300" swimtime="00:03:25.34" />
                    <SPLIT distance="350" swimtime="00:04:00.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-08-12" firstname="Konrad" gender="M" lastname="Plutecki" nation="POL" athleteid="9357">
              <RESULTS>
                <RESULT eventid="1075" points="695" reactiontime="+81" swimtime="00:00:25.89" resultid="9358" heatid="14155" lane="2" entrytime="00:00:27.27" entrycourse="SCM" />
                <RESULT eventid="1150" points="504" reactiontime="+87" swimtime="00:10:34.51" resultid="9359" heatid="14183" lane="3" entrytime="00:10:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.05" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                    <SPLIT distance="200" swimtime="00:02:30.57" />
                    <SPLIT distance="250" swimtime="00:03:10.22" />
                    <SPLIT distance="300" swimtime="00:03:49.96" />
                    <SPLIT distance="350" swimtime="00:04:30.58" />
                    <SPLIT distance="400" swimtime="00:05:10.86" />
                    <SPLIT distance="450" swimtime="00:05:51.30" />
                    <SPLIT distance="500" swimtime="00:06:31.97" />
                    <SPLIT distance="550" swimtime="00:07:13.46" />
                    <SPLIT distance="600" swimtime="00:07:55.23" />
                    <SPLIT distance="650" swimtime="00:08:36.03" />
                    <SPLIT distance="700" swimtime="00:09:17.14" />
                    <SPLIT distance="750" swimtime="00:09:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="452" reactiontime="+75" swimtime="00:00:33.76" resultid="9360" heatid="14203" lane="4" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="8277" points="672" reactiontime="+81" swimtime="00:00:57.81" resultid="9361" heatid="14235" lane="3" entrytime="00:00:57.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="506" reactiontime="+75" swimtime="00:01:17.45" resultid="9362" heatid="14282" lane="8" entrytime="00:01:18.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="559" reactiontime="+71" swimtime="00:02:13.56" resultid="9363" heatid="14329" lane="6" entrytime="00:02:20.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:03.94" />
                    <SPLIT distance="150" swimtime="00:01:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="546" reactiontime="+54" swimtime="00:02:33.13" resultid="9364" heatid="14369" lane="4" entrytime="00:02:38.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="566" reactiontime="+77" swimtime="00:04:56.54" resultid="9365" heatid="14400" lane="6" entrytime="00:05:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:46.87" />
                    <SPLIT distance="200" swimtime="00:02:25.40" />
                    <SPLIT distance="250" swimtime="00:03:04.00" />
                    <SPLIT distance="300" swimtime="00:03:42.93" />
                    <SPLIT distance="350" swimtime="00:04:21.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9583" name="Masters Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1970-03-11" firstname="ANNA" gender="F" lastname="GŁOWIAK" nation="POL" athleteid="9584">
              <RESULTS>
                <RESULT eventid="1058" points="558" reactiontime="+87" swimtime="00:00:33.17" resultid="9585" heatid="14139" lane="6" entrytime="00:00:32.39" />
                <RESULT eventid="1090" points="536" reactiontime="+81" swimtime="00:03:04.77" resultid="9586" heatid="14164" lane="1" entrytime="00:03:10.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:28.40" />
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="466" reactiontime="+93" swimtime="00:00:39.76" resultid="9587" heatid="14195" lane="4" entrytime="00:00:39.69" />
                <RESULT eventid="8261" points="563" swimtime="00:01:12.21" resultid="9588" heatid="14221" lane="5" entrytime="00:01:13.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="590" reactiontime="+63" swimtime="00:01:32.74" resultid="9589" heatid="14273" lane="9" entrytime="00:01:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="533" reactiontime="+99" swimtime="00:02:40.86" resultid="9590" heatid="14320" lane="3" entrytime="00:02:39.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="555" reactiontime="+67" swimtime="00:00:42.77" resultid="9591" heatid="14376" lane="8" entrytime="00:00:40.93" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12357" name="MASTERS Zdzieszowice">
          <CONTACT email="dejot.swim@gmail.com" name="Jajuga Dawid" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-12" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="12371">
              <RESULTS>
                <RESULT eventid="8293" points="583" reactiontime="+94" swimtime="00:01:22.87" resultid="12372" heatid="14241" lane="6" entrytime="00:01:22.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="632" reactiontime="+77" swimtime="00:01:21.53" resultid="12373" heatid="14306" lane="5" entrytime="00:01:22.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="570" reactiontime="+100" swimtime="00:06:29.93" resultid="12374" heatid="14341" lane="4" entrytime="00:06:40.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:20.12" />
                    <SPLIT distance="200" swimtime="00:03:08.11" />
                    <SPLIT distance="250" swimtime="00:04:04.86" />
                    <SPLIT distance="300" swimtime="00:05:02.17" />
                    <SPLIT distance="350" swimtime="00:05:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="657" reactiontime="+79" swimtime="00:02:56.80" resultid="12375" heatid="14365" lane="8" entrytime="00:02:54.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="528" reactiontime="+100" swimtime="00:05:51.01" resultid="12376" heatid="14394" lane="7" entrytime="00:05:54.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:08.35" />
                    <SPLIT distance="200" swimtime="00:02:53.76" />
                    <SPLIT distance="250" swimtime="00:03:39.34" />
                    <SPLIT distance="300" swimtime="00:04:24.44" />
                    <SPLIT distance="350" swimtime="00:05:08.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-21" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="12377">
              <RESULTS>
                <RESULT eventid="8229" status="DNS" swimtime="00:00:00.00" resultid="12378" heatid="14209" lane="5" entrytime="00:03:41.33" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="12379" heatid="14221" lane="9" entrytime="00:01:16.21" />
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="12380" heatid="14272" lane="8" entrytime="00:01:38.76" />
                <RESULT eventid="8502" status="DNS" swimtime="00:00:00.00" resultid="12381" heatid="14319" lane="4" entrytime="00:02:52.11" />
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="12382" heatid="14341" lane="7" entrytime="00:07:06.43" />
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="12383" heatid="14374" lane="3" entrytime="00:00:45.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="12364">
              <RESULTS>
                <RESULT eventid="8277" points="661" reactiontime="+84" swimtime="00:00:56.27" resultid="12365" heatid="14236" lane="5" entrytime="00:00:55.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="757" reactiontime="+88" swimtime="00:02:16.04" resultid="12366" heatid="14262" lane="2" entrytime="00:02:18.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                    <SPLIT distance="150" swimtime="00:01:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="12367" heatid="14301" lane="0" entrytime="00:00:27.11" />
                <RESULT eventid="8582" points="710" reactiontime="+75" swimtime="00:04:59.30" resultid="12368" heatid="14348" lane="7" entrytime="00:05:05.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:06.86" />
                    <SPLIT distance="150" swimtime="00:01:46.67" />
                    <SPLIT distance="200" swimtime="00:02:25.63" />
                    <SPLIT distance="250" swimtime="00:03:08.65" />
                    <SPLIT distance="300" swimtime="00:03:52.03" />
                    <SPLIT distance="350" swimtime="00:04:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="651" reactiontime="+74" swimtime="00:01:00.70" resultid="12369" heatid="14360" lane="7" entrytime="00:01:00.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="12370" heatid="14388" lane="4" entrytime="00:00:31.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-23" firstname="Szymon" gender="M" lastname="Paciej" nation="POL" athleteid="12358">
              <RESULTS>
                <RESULT eventid="8213" points="583" reactiontime="+91" swimtime="00:00:31.72" resultid="12359" heatid="14205" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="8245" points="574" reactiontime="+94" swimtime="00:02:49.01" resultid="12360" heatid="14216" lane="3" entrytime="00:02:46.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:02:04.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="593" reactiontime="+108" swimtime="00:01:08.52" resultid="12361" heatid="14314" lane="1" entrytime="00:01:08.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="539" reactiontime="+89" swimtime="00:05:28.01" resultid="12362" heatid="14347" lane="3" entrytime="00:05:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:59.22" />
                    <SPLIT distance="200" swimtime="00:02:41.99" />
                    <SPLIT distance="250" swimtime="00:03:28.86" />
                    <SPLIT distance="300" swimtime="00:04:16.33" />
                    <SPLIT distance="350" swimtime="00:04:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="465" reactiontime="+43" swimtime="00:02:30.55" resultid="12363" heatid="14371" lane="0" entrytime="00:02:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:51.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9971" name="MASTERS Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="9972">
              <RESULTS>
                <RESULT eventid="1075" points="679" reactiontime="+66" swimtime="00:00:26.16" resultid="9973" heatid="14157" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="8277" points="722" reactiontime="+87" swimtime="00:00:57.32" resultid="9974" heatid="14234" lane="7" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="507" reactiontime="+100" swimtime="00:02:38.73" resultid="9975" heatid="14260" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="646" reactiontime="+77" swimtime="00:00:28.77" resultid="9976" heatid="14298" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="8630" points="650" reactiontime="+81" swimtime="00:01:03.70" resultid="9977" heatid="14359" lane="0" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-01" firstname="Marek" gender="M" lastname="Gurbski" nation="POL" athleteid="9995">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1075" reactiontime="+43" status="DSQ" swimtime="00:00:28.43" resultid="9996" heatid="14149" lane="4" entrytime="00:00:30.36" />
                <RESULT eventid="8213" points="503" reactiontime="+75" swimtime="00:00:34.13" resultid="9997" heatid="14203" lane="1" entrytime="00:00:36.02" />
                <RESULT eventid="8277" points="526" reactiontime="+100" swimtime="00:01:04.50" resultid="9998" heatid="14228" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="455" reactiontime="+100" swimtime="00:00:32.66" resultid="9999" heatid="14294" lane="7" entrytime="00:00:33.34" />
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="10000" heatid="14312" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="8694" points="465" reactiontime="+102" swimtime="00:00:38.06" resultid="10001" heatid="14383" lane="1" entrytime="00:00:40.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-18" firstname="Paweł" gender="M" lastname="Lipka" nation="POL" athleteid="10035">
              <RESULTS>
                <RESULT eventid="1105" points="231" reactiontime="+92" swimtime="00:03:27.24" resultid="10036" heatid="14166" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:33.23" />
                    <SPLIT distance="150" swimtime="00:02:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="258" reactiontime="+90" swimtime="00:01:29.17" resultid="10037" heatid="14245" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="10075">
              <RESULTS>
                <RESULT eventid="1075" points="381" reactiontime="+80" swimtime="00:00:31.72" resultid="10076" heatid="14149" lane="7" entrytime="00:00:30.78" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10077" heatid="14248" lane="9" entrytime="00:01:22.66" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="10078" heatid="14279" lane="3" entrytime="00:01:28.46" />
                <RESULT eventid="8694" points="370" reactiontime="+84" swimtime="00:00:40.20" resultid="10079" heatid="14383" lane="4" entrytime="00:00:39.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-02" firstname="Ksawery" gender="M" lastname="Wiaderek" nation="POL" athleteid="10068">
              <RESULTS>
                <RESULT eventid="1075" points="547" reactiontime="+83" swimtime="00:00:27.05" resultid="10069" heatid="14156" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="8277" points="473" reactiontime="+94" swimtime="00:01:02.93" resultid="10070" heatid="14232" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="456" reactiontime="+81" swimtime="00:00:29.70" resultid="10071" heatid="14298" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-14" firstname="Anna" gender="F" lastname="Ostrowska" nation="POL" athleteid="10057">
              <RESULTS>
                <RESULT eventid="1058" points="667" reactiontime="+83" swimtime="00:00:31.10" resultid="10058" heatid="14140" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="8261" points="606" reactiontime="+84" swimtime="00:01:10.20" resultid="10059" heatid="14222" lane="9" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="591" reactiontime="+82" swimtime="00:00:35.59" resultid="10060" heatid="14287" lane="4" entrytime="00:00:37.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="10046">
              <RESULTS>
                <RESULT eventid="1075" points="518" reactiontime="+91" swimtime="00:00:29.57" resultid="10047" heatid="14151" lane="0" entrytime="00:00:29.99" />
                <RESULT eventid="1150" points="425" reactiontime="+92" swimtime="00:11:20.56" resultid="10048" heatid="14184" lane="7" entrytime="00:11:57.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:54.55" />
                    <SPLIT distance="200" swimtime="00:02:34.97" />
                    <SPLIT distance="250" swimtime="00:03:16.77" />
                    <SPLIT distance="300" swimtime="00:03:59.92" />
                    <SPLIT distance="350" swimtime="00:04:43.63" />
                    <SPLIT distance="400" swimtime="00:05:27.34" />
                    <SPLIT distance="450" swimtime="00:06:11.91" />
                    <SPLIT distance="500" swimtime="00:06:56.67" />
                    <SPLIT distance="550" swimtime="00:07:41.68" />
                    <SPLIT distance="600" swimtime="00:08:26.24" />
                    <SPLIT distance="650" swimtime="00:09:10.30" />
                    <SPLIT distance="700" swimtime="00:09:55.13" />
                    <SPLIT distance="750" swimtime="00:10:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="364" reactiontime="+101" swimtime="00:00:38.01" resultid="10049" heatid="14204" lane="1" entrytime="00:00:33.79" />
                <RESULT eventid="8277" points="478" reactiontime="+102" swimtime="00:01:06.58" resultid="10050" heatid="14231" lane="1" entrytime="00:01:04.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="442" reactiontime="+98" swimtime="00:02:28.32" resultid="10051" heatid="14328" lane="5" entrytime="00:02:25.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="9986">
              <RESULTS>
                <RESULT eventid="1075" points="675" reactiontime="+83" swimtime="00:00:27.08" resultid="9987" heatid="14156" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="1105" points="656" reactiontime="+81" swimtime="00:02:27.15" resultid="9988" heatid="14173" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="9989" heatid="14233" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="8309" points="713" reactiontime="+90" swimtime="00:01:06.93" resultid="9990" heatid="14251" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="614" reactiontime="+90" swimtime="00:00:29.56" resultid="9991" heatid="14297" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="8518" points="601" reactiontime="+93" swimtime="00:02:13.89" resultid="9992" heatid="14331" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="576" reactiontime="+84" swimtime="00:01:08.03" resultid="9993" heatid="14357" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Monika" gender="F" lastname="Klarecka" nation="POL" athleteid="10026">
              <RESULTS>
                <RESULT comment="przekroczony limit czasu" eventid="1135" reactiontime="+112" status="DSQ" swimtime="00:15:38.28" resultid="10027" heatid="14180" lane="9" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                    <SPLIT distance="100" swimtime="00:01:42.27" />
                    <SPLIT distance="150" swimtime="00:02:39.31" />
                    <SPLIT distance="200" swimtime="00:03:36.87" />
                    <SPLIT distance="250" swimtime="00:04:35.27" />
                    <SPLIT distance="300" swimtime="00:05:34.27" />
                    <SPLIT distance="350" swimtime="00:06:33.60" />
                    <SPLIT distance="400" swimtime="00:07:33.13" />
                    <SPLIT distance="450" swimtime="00:08:32.87" />
                    <SPLIT distance="500" swimtime="00:09:31.24" />
                    <SPLIT distance="550" swimtime="00:10:31.42" />
                    <SPLIT distance="600" swimtime="00:11:31.56" />
                    <SPLIT distance="650" swimtime="00:12:33.66" />
                    <SPLIT distance="700" swimtime="00:13:35.67" />
                    <SPLIT distance="750" swimtime="00:14:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="262" reactiontime="+113" swimtime="00:04:19.62" resultid="10028" heatid="14209" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.79" />
                    <SPLIT distance="100" swimtime="00:02:02.73" />
                    <SPLIT distance="150" swimtime="00:03:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="210" reactiontime="+128" swimtime="00:00:50.23" resultid="10029" heatid="14286" lane="0" entrytime="00:00:54.00" />
                <RESULT eventid="8502" points="204" reactiontime="+117" swimtime="00:03:39.47" resultid="10030" heatid="14318" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                    <SPLIT distance="150" swimtime="00:02:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="239" reactiontime="+146" swimtime="00:07:25.81" resultid="10031" heatid="14396" lane="6" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:36.26" />
                    <SPLIT distance="200" swimtime="00:03:33.39" />
                    <SPLIT distance="250" swimtime="00:04:31.92" />
                    <SPLIT distance="300" swimtime="00:05:29.99" />
                    <SPLIT distance="350" swimtime="00:06:29.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="10061">
              <RESULTS>
                <RESULT eventid="1075" points="524" reactiontime="+78" swimtime="00:00:28.52" resultid="10062" heatid="14153" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="10063" heatid="14215" lane="9" entrytime="00:03:10.00" />
                <RESULT eventid="8309" points="504" reactiontime="+76" swimtime="00:01:11.34" resultid="10064" heatid="14250" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="583" reactiontime="+80" swimtime="00:01:16.63" resultid="10065" heatid="14281" lane="8" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="540" reactiontime="+86" swimtime="00:00:30.55" resultid="10066" heatid="14296" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="8694" points="619" reactiontime="+79" swimtime="00:00:33.87" resultid="10067" heatid="14387" lane="2" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-11" firstname="Przemysław" gender="M" lastname="Michniewski" nation="POL" athleteid="10038">
              <RESULTS>
                <RESULT eventid="1075" points="662" reactiontime="+80" swimtime="00:00:26.39" resultid="10039" heatid="14157" lane="9" entrytime="00:00:26.50" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="10040" heatid="14170" lane="4" entrytime="00:02:45.00" />
                <RESULT eventid="8245" points="618" reactiontime="+88" swimtime="00:02:45.00" resultid="10041" heatid="14216" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                    <SPLIT distance="150" swimtime="00:02:01.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="689" reactiontime="+97" swimtime="00:01:04.29" resultid="10042" heatid="14253" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="716" reactiontime="+81" swimtime="00:01:11.56" resultid="10043" heatid="14283" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="673" reactiontime="+80" swimtime="00:00:28.39" resultid="10044" heatid="14299" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="8694" points="749" reactiontime="+84" swimtime="00:00:31.79" resultid="10045" heatid="14387" lane="3" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="9978">
              <RESULTS>
                <RESULT eventid="1105" points="696" reactiontime="+82" swimtime="00:02:23.65" resultid="9979" heatid="14170" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="688" reactiontime="+78" swimtime="00:00:29.52" resultid="9980" heatid="14203" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="8341" points="493" reactiontime="+103" swimtime="00:02:40.22" resultid="9981" heatid="14259" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="150" swimtime="00:01:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="704" reactiontime="+90" swimtime="00:01:11.94" resultid="9982" heatid="14279" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="693" reactiontime="+75" swimtime="00:01:03.78" resultid="9983" heatid="14312" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="572" reactiontime="+74" swimtime="00:02:26.42" resultid="9984" heatid="14369" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="706" reactiontime="+78" swimtime="00:00:32.42" resultid="9985" heatid="14383" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-30" firstname="Monika" gender="F" lastname="Kurstak-Jagiełło" nation="POL" athleteid="10032">
              <RESULTS>
                <RESULT eventid="1058" points="627" reactiontime="+86" swimtime="00:00:31.12" resultid="10033" heatid="14140" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="8196" points="539" reactiontime="+94" swimtime="00:00:39.15" resultid="10034" heatid="14196" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-08" firstname="Michał" gender="M" lastname="Olkowicz" nation="POL" athleteid="10053">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="10054" heatid="14145" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="10055" heatid="14202" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="8694" points="279" reactiontime="+87" swimtime="00:00:44.14" resultid="10056" heatid="14382" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Joanna" gender="F" lastname="Wilińska-Nowak" nation="POL" athleteid="10072">
              <RESULTS>
                <RESULT eventid="8325" points="715" reactiontime="+99" swimtime="00:02:45.63" resultid="10073" heatid="14257" lane="3" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="690" reactiontime="+94" swimtime="00:01:13.76" resultid="10074" heatid="14352" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-10-05" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" athleteid="10008">
              <RESULTS>
                <RESULT eventid="1075" points="556" reactiontime="+91" swimtime="00:00:27.96" resultid="10009" heatid="14154" lane="2" entrytime="00:00:27.77" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="10010" heatid="14184" lane="2" entrytime="00:11:57.77" />
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="10011" heatid="14215" lane="8" entrytime="00:03:07.77" />
                <RESULT eventid="8309" points="447" reactiontime="+84" swimtime="00:01:14.25" resultid="10012" heatid="14250" lane="3" entrytime="00:01:13.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="494" reactiontime="+78" swimtime="00:00:31.47" resultid="10013" heatid="14296" lane="9" entrytime="00:00:31.77" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="10014" heatid="14329" lane="2" entrytime="00:02:21.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-14" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="10023">
              <RESULTS>
                <RESULT eventid="1075" points="417" reactiontime="+94" swimtime="00:00:30.78" resultid="10024" heatid="14150" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="8213" points="380" swimtime="00:00:35.98" resultid="10025" heatid="14203" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="10015">
              <RESULTS>
                <RESULT eventid="1075" points="523" reactiontime="+92" swimtime="00:00:28.54" resultid="10016" heatid="14144" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1105" points="361" reactiontime="+106" swimtime="00:02:58.79" resultid="10017" heatid="14169" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="384" reactiontime="+96" swimtime="00:01:18.09" resultid="10018" heatid="14246" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="307" reactiontime="+108" swimtime="00:01:23.63" resultid="10019" heatid="14310" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="278" reactiontime="+103" swimtime="00:06:58.04" resultid="10020" heatid="14343" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:03:22.70" />
                    <SPLIT distance="200" swimtime="00:04:20.51" />
                    <SPLIT distance="250" swimtime="00:05:20.16" />
                    <SPLIT distance="300" swimtime="00:06:09.98" />
                    <SPLIT distance="350" swimtime="00:06:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="296" reactiontime="+83" swimtime="00:03:02.27" resultid="10021" heatid="14368" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:27.12" />
                    <SPLIT distance="150" swimtime="00:02:16.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="428" reactiontime="+87" swimtime="00:00:38.29" resultid="10022" heatid="14382" lane="6" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+81" swimtime="00:01:56.70" resultid="10082" heatid="14267" lane="3" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:01.46" />
                    <SPLIT distance="150" swimtime="00:01:29.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9978" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="10038" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="9972" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="10068" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+93" swimtime="00:02:09.10" resultid="10083" heatid="14267" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:42.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10015" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="10061" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="10008" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="9986" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+82" swimtime="00:02:21.28" resultid="10084" heatid="14266" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="150" swimtime="00:01:52.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10023" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="10035" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="10046" number="3" />
                    <RELAYPOSITION athleteid="9995" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+80" swimtime="00:01:45.41" resultid="10086" heatid="14339" lane="8" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:00:52.81" />
                    <SPLIT distance="150" swimtime="00:01:18.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9986" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="10038" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="9972" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="10068" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8550" reactiontime="+69" status="DSQ" swimtime="00:01:53.83" resultid="10087" heatid="14338" lane="6" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:00:57.80" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10008" number="1" reactiontime="+69" status="DSQ" />
                    <RELAYPOSITION athleteid="10061" number="2" reactiontime="+41" status="DSQ" />
                    <RELAYPOSITION athleteid="10046" number="3" reactiontime="+26" status="DSQ" />
                    <RELAYPOSITION athleteid="9978" number="4" reactiontime="+50" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="8550" swimtime="00:02:06.36" resultid="10088" heatid="14337" lane="6" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="150" swimtime="00:01:32.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9995" number="1" />
                    <RELAYPOSITION athleteid="10075" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10023" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="10035" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="8357" status="DNS" swimtime="00:00:00.00" resultid="10081" heatid="14264" lane="0" entrytime="00:02:33.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10057" number="1" />
                    <RELAYPOSITION athleteid="10026" number="2" />
                    <RELAYPOSITION athleteid="10072" number="3" />
                    <RELAYPOSITION athleteid="10032" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="6">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8534" reactiontime="+82" status="DSQ" swimtime="00:02:15.42" resultid="10085" heatid="14335" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10057" number="1" reactiontime="+82" status="DSQ" />
                    <RELAYPOSITION athleteid="10026" number="2" reactiontime="+97" status="DSQ" />
                    <RELAYPOSITION athleteid="10072" number="3" reactiontime="-54" status="DSQ" />
                    <RELAYPOSITION athleteid="10032" number="4" reactiontime="+27" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+87" swimtime="00:01:53.84" resultid="10080" heatid="14177" lane="8" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:02.43" />
                    <SPLIT distance="150" swimtime="00:01:27.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10057" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="10032" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="9972" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="10068" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="10">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+77" swimtime="00:02:10.91" resultid="10089" heatid="14392" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:39.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10032" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="10038" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="9972" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="10057" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="13280" name="Masters Ślęza">
          <CONTACT name="Masters Ślęza" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="13290">
              <RESULTS>
                <RESULT eventid="1058" points="470" reactiontime="+83" swimtime="00:00:38.02" resultid="13291" heatid="14136" lane="4" entrytime="00:00:38.60" />
                <RESULT eventid="8229" points="528" reactiontime="+84" swimtime="00:03:49.08" resultid="13292" heatid="14209" lane="2" entrytime="00:03:51.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.96" />
                    <SPLIT distance="100" swimtime="00:01:47.81" />
                    <SPLIT distance="150" swimtime="00:02:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="417" reactiontime="+83" swimtime="00:01:40.58" resultid="13293" heatid="14239" lane="6" entrytime="00:01:39.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="536" reactiontime="+80" swimtime="00:01:42.99" resultid="13294" heatid="14271" lane="6" entrytime="00:01:44.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="559" reactiontime="+79" swimtime="00:00:45.59" resultid="13295" heatid="14374" lane="1" entrytime="00:00:47.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-11" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="13281">
              <RESULTS>
                <RESULT eventid="1058" points="552" reactiontime="+90" swimtime="00:00:33.30" resultid="13282" heatid="14138" lane="7" entrytime="00:00:34.34" />
                <RESULT eventid="1090" points="486" reactiontime="+94" swimtime="00:03:10.88" resultid="13283" heatid="14165" lane="9" entrytime="00:02:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:29.41" />
                    <SPLIT distance="150" swimtime="00:02:23.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="482" reactiontime="+93" swimtime="00:01:16.05" resultid="13284" heatid="14220" lane="8" entrytime="00:01:19.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="521" reactiontime="+99" swimtime="00:01:26.05" resultid="13285" heatid="14241" lane="9" entrytime="00:01:28.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="525" reactiontime="+91" swimtime="00:00:37.19" resultid="13286" heatid="14287" lane="9" entrytime="00:00:39.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-11" firstname="Marta" gender="F" lastname="Burandt" nation="POL" athleteid="13287">
              <RESULTS>
                <RESULT eventid="1165" points="434" reactiontime="+123" swimtime="00:25:37.57" resultid="13288" heatid="14188" lane="5" entrytime="00:26:05.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:14.87" />
                    <SPLIT distance="200" swimtime="00:03:04.38" />
                    <SPLIT distance="250" swimtime="00:03:55.10" />
                    <SPLIT distance="300" swimtime="00:04:46.06" />
                    <SPLIT distance="350" swimtime="00:05:37.27" />
                    <SPLIT distance="400" swimtime="00:06:28.81" />
                    <SPLIT distance="450" swimtime="00:07:20.79" />
                    <SPLIT distance="500" swimtime="00:08:12.76" />
                    <SPLIT distance="550" swimtime="00:09:05.11" />
                    <SPLIT distance="600" swimtime="00:09:57.73" />
                    <SPLIT distance="650" swimtime="00:10:50.30" />
                    <SPLIT distance="700" swimtime="00:11:43.28" />
                    <SPLIT distance="750" swimtime="00:12:35.30" />
                    <SPLIT distance="800" swimtime="00:13:27.97" />
                    <SPLIT distance="850" swimtime="00:14:20.41" />
                    <SPLIT distance="900" swimtime="00:15:12.55" />
                    <SPLIT distance="950" swimtime="00:16:04.59" />
                    <SPLIT distance="1000" swimtime="00:16:56.87" />
                    <SPLIT distance="1050" swimtime="00:17:48.88" />
                    <SPLIT distance="1100" swimtime="00:18:40.93" />
                    <SPLIT distance="1150" swimtime="00:19:32.48" />
                    <SPLIT distance="1200" swimtime="00:20:24.06" />
                    <SPLIT distance="1250" swimtime="00:21:16.32" />
                    <SPLIT distance="1300" swimtime="00:22:09.25" />
                    <SPLIT distance="1350" swimtime="00:23:01.74" />
                    <SPLIT distance="1400" swimtime="00:23:53.93" />
                    <SPLIT distance="1450" swimtime="00:24:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="403" reactiontime="+96" swimtime="00:01:33.68" resultid="13289" heatid="14240" lane="9" entrytime="00:01:35.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="SZ" clubid="9560" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="9568">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9569" heatid="14146" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="9570">
              <RESULTS>
                <RESULT eventid="1105" points="539" reactiontime="+84" swimtime="00:03:18.52" resultid="9571" heatid="14169" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:32.38" />
                    <SPLIT distance="150" swimtime="00:02:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="634" reactiontime="+101" swimtime="00:03:31.98" resultid="9572" heatid="14213" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:44.15" />
                    <SPLIT distance="150" swimtime="00:02:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="9573" heatid="14275" lane="3" />
                <RESULT eventid="8454" points="560" reactiontime="+97" swimtime="00:00:37.07" resultid="9574" heatid="14293" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="8694" points="636" reactiontime="+85" swimtime="00:00:40.57" resultid="9575" heatid="14382" lane="3" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="9561">
              <RESULTS>
                <RESULT eventid="8196" points="826" reactiontime="+93" swimtime="00:00:41.02" resultid="9562" heatid="14195" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="8261" points="734" reactiontime="+108" swimtime="00:01:19.13" resultid="9563" heatid="14220" lane="1" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="892" reactiontime="+86" swimtime="00:01:27.14" resultid="9564" heatid="14305" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="781" reactiontime="+124" swimtime="00:02:52.55" resultid="9565" heatid="14319" lane="2" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="981" reactiontime="+91" swimtime="00:03:04.07" resultid="9566" heatid="14364" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:17.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="861" reactiontime="+91" swimtime="00:06:08.02" resultid="9567" heatid="14395" lane="3" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:02:14.18" />
                    <SPLIT distance="150" swimtime="00:03:48.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06611" nation="POL" region="SLA" clubid="10590" name="MKP Wodnik 29 Tychy">
          <CONTACT city="Tychy" email="marekmrozw29@gmail.com" internet="https://www.facebook.com/wodnik29tychy/" name="Marek Mróz" phone="782985239" state="SLA" street="Damrota 170" zip="43-100" />
          <ATHLETES>
            <ATHLETE birthdate="1995-07-13" firstname="Szymon" gender="M" lastname="Warwas" nation="POL" license="106611700009" athleteid="10591">
              <RESULTS>
                <RESULT eventid="1075" points="852" reactiontime="+78" swimtime="00:00:24.19" resultid="10592" heatid="14161" lane="0" entrytime="00:00:23.80" />
                <RESULT eventid="8213" points="761" reactiontime="+72" swimtime="00:00:28.37" resultid="10593" heatid="14207" lane="7" entrytime="00:00:28.30" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="10594" heatid="14237" lane="9" entrytime="00:00:55.00" />
                <RESULT eventid="8309" points="690" reactiontime="+75" swimtime="00:01:03.62" resultid="10595" heatid="14254" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="818" reactiontime="+68" swimtime="00:00:26.47" resultid="10596" heatid="14301" lane="3" entrytime="00:00:26.20" />
                <RESULT eventid="8486" points="638" reactiontime="+79" swimtime="00:01:04.07" resultid="10597" heatid="14315" lane="7" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="ZAC" clubid="10470" name="MKS Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1973-02-20" firstname="Mariusz" gender="M" lastname="Chrzan" nation="POL" athleteid="10471">
              <RESULTS>
                <RESULT eventid="1075" points="701" reactiontime="+99" swimtime="00:00:26.86" resultid="10472" heatid="14158" lane="8" entrytime="00:00:26.10" />
                <RESULT eventid="1105" points="834" reactiontime="+83" swimtime="00:02:23.70" resultid="10473" heatid="14173" lane="2" entrytime="00:02:26.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="782" reactiontime="+80" swimtime="00:00:30.24" resultid="10474" heatid="14206" lane="6" entrytime="00:00:30.45" />
                <RESULT eventid="8309" points="805" reactiontime="+75" swimtime="00:01:04.55" resultid="10475" heatid="14253" lane="4" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="827" reactiontime="+69" swimtime="00:00:28.16" resultid="10476" heatid="14300" lane="9" entrytime="00:00:28.20" />
                <RESULT eventid="8486" points="788" reactiontime="+96" swimtime="00:01:04.37" resultid="10477" heatid="14315" lane="9" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="885" reactiontime="+82" swimtime="00:02:21.94" resultid="10478" heatid="14371" lane="1" entrytime="00:02:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="150" swimtime="00:01:46.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" region="DOL" clubid="9576" name="MKS Swim Academy Termy Jakuba Oława" shortname="MKS Swim Academy Termy Jakuba ">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOL" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-27" firstname="Magdalena" gender="F" lastname="Mruk" nation="POL" license="104501600044" athleteid="9577">
              <RESULTS>
                <RESULT eventid="8229" points="673" reactiontime="+107" swimtime="00:03:09.49" resultid="9578" heatid="14211" lane="2" entrytime="00:03:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="687" reactiontime="+92" swimtime="00:01:17.19" resultid="9579" heatid="14242" lane="7" entrytime="00:01:19.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="723" reactiontime="+105" swimtime="00:01:24.30" resultid="9580" heatid="14274" lane="0" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="641" reactiontime="+92" swimtime="00:00:34.63" resultid="9581" heatid="14289" lane="0" entrytime="00:00:32.80" />
                <RESULT eventid="8678" points="745" reactiontime="+82" swimtime="00:00:37.87" resultid="9582" heatid="14377" lane="8" entrytime="00:00:38.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="PDK" clubid="9592" name="Motyl MOSIR Stalowa Wola">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="600831914" street="Hutnicza 15" zip="37=450" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="9601">
              <RESULTS>
                <RESULT eventid="1058" points="510" reactiontime="+99" swimtime="00:00:35.66" resultid="9602" heatid="14137" lane="1" entrytime="00:00:37.01" />
                <RESULT eventid="1090" points="564" reactiontime="+96" swimtime="00:03:07.97" resultid="9603" heatid="14163" lane="4" entrytime="00:03:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:31.10" />
                    <SPLIT distance="150" swimtime="00:02:24.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="556" reactiontime="+102" swimtime="00:03:35.80" resultid="9604" heatid="14210" lane="1" entrytime="00:03:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:44.37" />
                    <SPLIT distance="150" swimtime="00:02:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="571" reactiontime="+95" swimtime="00:01:26.34" resultid="9605" heatid="14240" lane="4" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="482" reactiontime="+95" swimtime="00:01:42.30" resultid="9606" heatid="14271" lane="3" entrytime="00:01:42.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="491" reactiontime="+104" swimtime="00:00:39.48" resultid="9607" heatid="14287" lane="0" entrytime="00:00:39.10" />
                <RESULT eventid="8613" points="405" reactiontime="+91" swimtime="00:01:35.60" resultid="9608" heatid="14350" lane="5" entrytime="00:01:36.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="513" reactiontime="+92" swimtime="00:00:45.58" resultid="9609" heatid="14374" lane="7" entrytime="00:00:47.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" athleteid="9626">
              <RESULTS>
                <RESULT eventid="8179" points="668" reactiontime="+84" swimtime="00:18:16.83" resultid="9627" heatid="14189" lane="8" entrytime="00:19:02.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:43.61" />
                    <SPLIT distance="200" swimtime="00:02:20.04" />
                    <SPLIT distance="250" swimtime="00:02:56.42" />
                    <SPLIT distance="300" swimtime="00:03:32.90" />
                    <SPLIT distance="350" swimtime="00:04:09.49" />
                    <SPLIT distance="400" swimtime="00:04:46.06" />
                    <SPLIT distance="450" swimtime="00:05:22.73" />
                    <SPLIT distance="500" swimtime="00:05:59.45" />
                    <SPLIT distance="550" swimtime="00:06:35.93" />
                    <SPLIT distance="600" swimtime="00:07:13.06" />
                    <SPLIT distance="650" swimtime="00:07:49.27" />
                    <SPLIT distance="700" swimtime="00:08:26.19" />
                    <SPLIT distance="750" swimtime="00:09:02.57" />
                    <SPLIT distance="800" swimtime="00:09:39.58" />
                    <SPLIT distance="850" swimtime="00:10:16.57" />
                    <SPLIT distance="900" swimtime="00:10:53.37" />
                    <SPLIT distance="950" swimtime="00:11:30.53" />
                    <SPLIT distance="1000" swimtime="00:12:07.85" />
                    <SPLIT distance="1050" swimtime="00:12:44.97" />
                    <SPLIT distance="1100" swimtime="00:13:22.04" />
                    <SPLIT distance="1150" swimtime="00:13:59.22" />
                    <SPLIT distance="1200" swimtime="00:14:36.72" />
                    <SPLIT distance="1250" swimtime="00:15:14.09" />
                    <SPLIT distance="1300" swimtime="00:15:51.49" />
                    <SPLIT distance="1350" swimtime="00:16:28.79" />
                    <SPLIT distance="1400" swimtime="00:17:06.27" />
                    <SPLIT distance="1450" swimtime="00:17:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="557" reactiontime="+91" swimtime="00:02:31.64" resultid="9628" heatid="14261" lane="2" entrytime="00:02:35.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="625" reactiontime="+92" swimtime="00:02:08.63" resultid="9629" heatid="14331" lane="3" entrytime="00:02:12.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="599" reactiontime="+82" swimtime="00:05:18.20" resultid="9630" heatid="14348" lane="9" entrytime="00:05:22.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:51.82" />
                    <SPLIT distance="200" swimtime="00:02:32.08" />
                    <SPLIT distance="250" swimtime="00:03:19.95" />
                    <SPLIT distance="300" swimtime="00:04:07.79" />
                    <SPLIT distance="350" swimtime="00:04:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="640" reactiontime="+77" swimtime="00:02:25.17" resultid="9631" heatid="14370" lane="7" entrytime="00:02:32.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="753" reactiontime="+86" swimtime="00:04:29.72" resultid="9632" heatid="14399" lane="6" entrytime="00:04:38.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="150" swimtime="00:01:37.81" />
                    <SPLIT distance="200" swimtime="00:02:11.61" />
                    <SPLIT distance="250" swimtime="00:02:46.12" />
                    <SPLIT distance="300" swimtime="00:03:20.83" />
                    <SPLIT distance="350" swimtime="00:03:55.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="9610">
              <RESULTS>
                <RESULT eventid="1075" points="683" reactiontime="+85" swimtime="00:00:26.97" resultid="9611" heatid="14155" lane="4" entrytime="00:00:27.01" />
                <RESULT eventid="8213" points="745" reactiontime="+99" swimtime="00:00:29.94" resultid="9612" heatid="14206" lane="3" entrytime="00:00:30.27" />
                <RESULT eventid="8277" points="673" reactiontime="+83" swimtime="00:00:59.39" resultid="9613" heatid="14233" lane="8" entrytime="00:01:00.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="749" reactiontime="+95" swimtime="00:01:05.03" resultid="9614" heatid="14314" lane="6" entrytime="00:01:07.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="736" reactiontime="+86" swimtime="00:02:24.46" resultid="9615" heatid="14370" lane="2" entrytime="00:02:32.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="9616" heatid="14384" lane="7" entrytime="00:00:38.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="9633">
              <RESULTS>
                <RESULT eventid="1105" points="963" reactiontime="+86" swimtime="00:02:16.95" resultid="9634" heatid="14174" lane="2" entrytime="00:02:18.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                    <SPLIT distance="150" swimtime="00:01:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="842" reactiontime="+71" swimtime="00:00:56.03" resultid="9635" heatid="14236" lane="7" entrytime="00:00:56.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="871" reactiontime="+82" swimtime="00:01:02.90" resultid="9636" heatid="14254" lane="2" entrytime="00:01:03.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="789" reactiontime="+80" swimtime="00:02:04.11" resultid="9637" heatid="14333" lane="8" entrytime="00:02:04.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="100" swimtime="00:00:59.92" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="880" reactiontime="+86" swimtime="00:05:01.59" resultid="9638" heatid="14348" lane="2" entrytime="00:05:04.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:08.52" />
                    <SPLIT distance="150" swimtime="00:01:48.26" />
                    <SPLIT distance="200" swimtime="00:02:26.99" />
                    <SPLIT distance="250" swimtime="00:03:09.36" />
                    <SPLIT distance="300" swimtime="00:03:51.95" />
                    <SPLIT distance="350" swimtime="00:04:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="963" reactiontime="+74" swimtime="00:00:59.54" resultid="9639" heatid="14360" lane="6" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="772" reactiontime="+82" swimtime="00:04:27.95" resultid="9640" heatid="14398" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="150" swimtime="00:01:40.72" />
                    <SPLIT distance="200" swimtime="00:02:15.63" />
                    <SPLIT distance="250" swimtime="00:02:49.97" />
                    <SPLIT distance="300" swimtime="00:03:24.14" />
                    <SPLIT distance="350" swimtime="00:03:57.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="9617">
              <RESULTS>
                <RESULT eventid="1105" points="504" reactiontime="+93" swimtime="00:02:40.69" resultid="9618" heatid="14170" lane="2" entrytime="00:02:52.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:02:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="463" reactiontime="+87" swimtime="00:11:01.17" resultid="9619" heatid="14184" lane="6" entrytime="00:11:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                    <SPLIT distance="200" swimtime="00:02:40.01" />
                    <SPLIT distance="250" swimtime="00:03:21.39" />
                    <SPLIT distance="300" swimtime="00:04:03.49" />
                    <SPLIT distance="350" swimtime="00:04:45.45" />
                    <SPLIT distance="400" swimtime="00:05:27.37" />
                    <SPLIT distance="450" swimtime="00:06:08.94" />
                    <SPLIT distance="500" swimtime="00:06:50.65" />
                    <SPLIT distance="550" swimtime="00:07:32.92" />
                    <SPLIT distance="600" swimtime="00:08:14.92" />
                    <SPLIT distance="650" swimtime="00:08:57.28" />
                    <SPLIT distance="700" swimtime="00:09:39.32" />
                    <SPLIT distance="750" swimtime="00:10:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="9620" heatid="14205" lane="0" entrytime="00:00:32.51" />
                <RESULT eventid="8309" points="581" reactiontime="+85" swimtime="00:01:11.67" resultid="9621" heatid="14250" lane="4" entrytime="00:01:12.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="551" reactiontime="+94" swimtime="00:01:12.03" resultid="9622" heatid="14313" lane="7" entrytime="00:01:11.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="453" reactiontime="+84" swimtime="00:05:52.92" resultid="9623" heatid="14346" lane="6" entrytime="00:06:03.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:23.71" />
                    <SPLIT distance="150" swimtime="00:02:08.22" />
                    <SPLIT distance="200" swimtime="00:02:52.01" />
                    <SPLIT distance="250" swimtime="00:03:40.63" />
                    <SPLIT distance="300" swimtime="00:04:30.77" />
                    <SPLIT distance="350" swimtime="00:05:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" status="DNS" swimtime="00:00:00.00" resultid="9624" heatid="14369" lane="8" entrytime="00:03:01.50" />
                <RESULT eventid="8694" points="585" reactiontime="+79" swimtime="00:00:35.26" resultid="9625" heatid="14386" lane="2" entrytime="00:00:35.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="9593">
              <RESULTS>
                <RESULT eventid="1105" points="595" reactiontime="+86" swimtime="00:02:52.85" resultid="9594" heatid="14170" lane="8" entrytime="00:02:58.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:02:13.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="619" reactiontime="+98" swimtime="00:01:08.08" resultid="9595" heatid="14228" lane="4" entrytime="00:01:09.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="467" reactiontime="+98" swimtime="00:03:10.22" resultid="9596" heatid="14260" lane="0" entrytime="00:03:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:01:29.61" />
                    <SPLIT distance="150" swimtime="00:02:20.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="623" reactiontime="+159" swimtime="00:02:33.42" resultid="9597" heatid="14327" lane="6" entrytime="00:02:36.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:53.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="655" reactiontime="+84" swimtime="00:06:11.53" resultid="9598" heatid="14346" lane="7" entrytime="00:06:24.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="150" swimtime="00:02:13.71" />
                    <SPLIT distance="200" swimtime="00:02:59.20" />
                    <SPLIT distance="250" swimtime="00:03:54.91" />
                    <SPLIT distance="300" swimtime="00:04:48.77" />
                    <SPLIT distance="350" swimtime="00:05:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="558" reactiontime="+81" swimtime="00:02:53.98" resultid="9599" heatid="14368" lane="4" entrytime="00:03:02.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="622" reactiontime="+87" swimtime="00:05:32.13" resultid="9600" heatid="14402" lane="4" entrytime="00:05:58.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                    <SPLIT distance="200" swimtime="00:02:42.55" />
                    <SPLIT distance="250" swimtime="00:03:25.82" />
                    <SPLIT distance="300" swimtime="00:04:09.13" />
                    <SPLIT distance="350" swimtime="00:04:52.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" status="DNS" swimtime="00:00:00.00" resultid="10837" heatid="14265" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9610" number="1" />
                    <RELAYPOSITION athleteid="9617" number="2" />
                    <RELAYPOSITION athleteid="9633" number="3" />
                    <RELAYPOSITION athleteid="9593" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00403" nation="POL" region="03" clubid="8852" name="MUKS Lider Chełm">
          <ATHLETES>
            <ATHLETE birthdate="1941-11-10" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="8853">
              <RESULTS>
                <RESULT eventid="8245" points="441" reactiontime="+112" swimtime="00:04:16.89" resultid="8854" heatid="14212" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                    <SPLIT distance="100" swimtime="00:02:04.14" />
                    <SPLIT distance="150" swimtime="00:03:11.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="407" reactiontime="+131" swimtime="00:04:36.83" resultid="8855" heatid="14258" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.24" />
                    <SPLIT distance="100" swimtime="00:02:16.75" />
                    <SPLIT distance="150" swimtime="00:03:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="531" reactiontime="+122" swimtime="00:01:47.09" resultid="8856" heatid="14277" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="344" reactiontime="+117" swimtime="00:00:49.30" resultid="8857" heatid="14291" lane="6" entrytime="00:00:48.25" />
                <RESULT eventid="8630" points="405" reactiontime="+110" swimtime="00:01:54.97" resultid="8858" heatid="14354" lane="6" entrytime="00:01:55.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="632" reactiontime="+123" swimtime="00:00:45.67" resultid="8859" heatid="14382" lane="9" entrytime="00:00:45.35" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8782" name="Nabaiji Team Decathlon">
          <CONTACT email="rafal.liszewski@decathlon.com" name="Liszewski Rafal" phone="663643393" />
          <ATHLETES>
            <ATHLETE birthdate="1994-06-25" firstname="Filip" gender="M" lastname="Wasielewski" nation="POL" athleteid="10762">
              <RESULTS>
                <RESULT eventid="1075" points="592" reactiontime="+66" swimtime="00:00:27.31" resultid="10763" heatid="14155" lane="9" entrytime="00:00:27.50" />
                <RESULT eventid="8277" points="574" reactiontime="+72" swimtime="00:01:00.93" resultid="10764" heatid="14233" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="590" reactiontime="+69" swimtime="00:00:29.52" resultid="10765" heatid="14297" lane="7" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-11-23" firstname="Filip" gender="M" lastname="Kolodziejski" nation="POL" athleteid="10791">
              <RESULTS>
                <RESULT eventid="1075" points="913" reactiontime="+65" swimtime="00:00:23.64" resultid="10792" heatid="14161" lane="7" entrytime="00:00:23.50" />
                <RESULT eventid="8213" points="958" reactiontime="+75" swimtime="00:00:26.28" resultid="10793" heatid="14207" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="8277" points="958" reactiontime="+72" swimtime="00:00:51.39" resultid="10794" heatid="14237" lane="3" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="891" reactiontime="+77" swimtime="00:00:57.32" resultid="10795" heatid="14315" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="905" reactiontime="+65" swimtime="00:00:56.15" resultid="10796" heatid="14361" lane="5" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-08-24" firstname="Aleksandra" gender="F" lastname="Czechowicz" nation="POL" athleteid="10787">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="10788" heatid="14136" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="8261" points="211" reactiontime="+100" swimtime="00:01:37.20" resultid="10789" heatid="14219" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" status="DNS" swimtime="00:00:00.00" resultid="10790" heatid="14305" lane="9" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-20" firstname="Maciej" gender="M" lastname="Jekielek" nation="POL" athleteid="10797">
              <RESULTS>
                <RESULT eventid="1075" points="645" reactiontime="+74" swimtime="00:00:26.43" resultid="10798" heatid="14157" lane="7" entrytime="00:00:26.50" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10799" heatid="14252" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="8406" points="525" reactiontime="+92" swimtime="00:01:16.88" resultid="10800" heatid="14282" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="10801" heatid="14387" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-13" firstname="Agata" gender="F" lastname="Koc" nation="POL" athleteid="10807">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="10808" heatid="14140" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="10809" heatid="14222" lane="2" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-06" firstname="Pawel" gender="M" lastname="Bednarczyk" nation="POL" athleteid="10771">
              <RESULTS>
                <RESULT eventid="1075" points="822" reactiontime="+78" swimtime="00:00:24.48" resultid="10772" heatid="14160" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="8277" points="829" reactiontime="+73" swimtime="00:00:53.92" resultid="10773" heatid="14237" lane="7" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10774" heatid="14254" lane="4" entrytime="00:01:02.00" />
                <RESULT eventid="8454" points="870" swimtime="00:00:25.93" resultid="10775" heatid="14302" lane="3" entrytime="00:00:25.00" />
                <RESULT eventid="8630" points="671" reactiontime="+74" swimtime="00:01:02.02" resultid="10776" heatid="14361" lane="8" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="10746">
              <RESULTS>
                <RESULT eventid="1058" points="616" reactiontime="+86" swimtime="00:00:30.72" resultid="10747" heatid="14140" lane="3" entrytime="00:00:30.70" />
                <RESULT eventid="8261" points="605" reactiontime="+81" swimtime="00:01:07.92" resultid="10748" heatid="14222" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="596" reactiontime="+97" swimtime="00:02:29.57" resultid="10749" heatid="14320" lane="4" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:51.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-20" firstname="Rafal" gender="M" lastname="Liszewski" nation="POL" athleteid="10727">
              <RESULTS>
                <RESULT eventid="1075" points="570" reactiontime="+75" swimtime="00:00:26.68" resultid="10728" heatid="14156" lane="7" entrytime="00:00:26.80" entrycourse="SCM" />
                <RESULT eventid="8309" points="492" reactiontime="+78" swimtime="00:01:09.65" resultid="10729" heatid="14251" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="560" reactiontime="+79" swimtime="00:01:14.39" resultid="10730" heatid="14282" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="660" reactiontime="+79" swimtime="00:00:31.93" resultid="10731" heatid="14388" lane="1" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-03" firstname="Mateusz" gender="M" lastname="Turowski" nation="POL" athleteid="10758">
              <RESULTS>
                <RESULT eventid="1075" points="473" reactiontime="+101" swimtime="00:00:29.31" resultid="10759" heatid="14154" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="8277" points="358" reactiontime="+104" swimtime="00:01:08.39" resultid="10760" heatid="14233" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="378" reactiontime="+93" swimtime="00:00:32.75" resultid="10761" heatid="14297" lane="8" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-25" firstname="Mateusz" gender="M" lastname="Kołodziejski" nation="POL" athleteid="9026">
              <RESULTS>
                <RESULT eventid="1075" points="932" reactiontime="+73" swimtime="00:00:23.38" resultid="9027" heatid="14161" lane="2" entrytime="00:00:23.47" />
                <RESULT eventid="8309" points="867" reactiontime="+68" swimtime="00:00:57.88" resultid="9028" heatid="14255" lane="6" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="943" reactiontime="+70" swimtime="00:01:03.25" resultid="9029" heatid="14284" lane="5" entrytime="00:01:02.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="801" swimtime="00:00:25.51" resultid="9030" heatid="14302" lane="7" entrytime="00:00:25.22" />
                <RESULT eventid="8694" points="921" reactiontime="+64" swimtime="00:00:29.04" resultid="9031" heatid="14389" lane="4" entrytime="00:00:28.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-29" firstname="Kamil" gender="M" lastname="Ziemianin" nation="POL" athleteid="10780">
              <RESULTS>
                <RESULT eventid="8245" points="564" reactiontime="+95" swimtime="00:02:47.47" resultid="10781" heatid="14216" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:02:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="602" reactiontime="+92" swimtime="00:01:13.44" resultid="10782" heatid="14282" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="674" reactiontime="+81" swimtime="00:00:32.23" resultid="10783" heatid="14388" lane="8" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-18" firstname="EMIL" gender="M" lastname="STRUMIŃSKI" nation="POL" athleteid="9478">
              <RESULTS>
                <RESULT eventid="1075" points="576" reactiontime="+78" swimtime="00:00:26.59" resultid="9479" heatid="14158" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1105" points="510" reactiontime="+79" swimtime="00:02:27.77" resultid="9480" heatid="14173" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="603" reactiontime="+80" swimtime="00:00:58.04" resultid="9481" heatid="14235" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="9482" heatid="14250" lane="1" entrytime="00:01:15.00" />
                <RESULT eventid="8454" points="528" reactiontime="+79" swimtime="00:00:28.29" resultid="9483" heatid="14299" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="8518" points="513" reactiontime="+90" swimtime="00:02:13.02" resultid="9484" heatid="14331" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                    <SPLIT distance="150" swimtime="00:01:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9485" heatid="14357" lane="2" entrytime="00:01:11.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-07" firstname="Marzena" gender="F" lastname="Mikolajek" nation="POL" athleteid="10777">
              <RESULTS>
                <RESULT eventid="1058" points="431" reactiontime="+102" swimtime="00:00:34.08" resultid="10778" heatid="14137" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="8261" points="363" reactiontime="+106" swimtime="00:01:18.65" resultid="10779" heatid="14220" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-06" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="10738">
              <RESULTS>
                <RESULT eventid="1058" points="527" reactiontime="+84" swimtime="00:00:32.21" resultid="10739" heatid="14139" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="8293" points="458" reactiontime="+78" swimtime="00:01:21.92" resultid="10740" heatid="14241" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-13" firstname="Aleksander" gender="M" lastname="Zieminski" nation="POL" athleteid="10735">
              <RESULTS>
                <RESULT eventid="1075" points="255" reactiontime="+84" swimtime="00:00:36.14" resultid="10736" heatid="14146" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="8406" points="194" reactiontime="+97" swimtime="00:01:46.58" resultid="10737" heatid="14278" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-02-05" firstname="Ewelina" gender="F" lastname="Radonska" nation="POL" athleteid="10784">
              <RESULTS>
                <RESULT eventid="8196" points="339" reactiontime="+87" swimtime="00:00:41.99" resultid="10785" heatid="14196" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="8470" points="314" reactiontime="+93" swimtime="00:01:34.73" resultid="10786" heatid="14307" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-02" firstname="Karolina" gender="F" lastname="Mazurek-Swistak" nation="POL" athleteid="10741">
              <RESULTS>
                <RESULT eventid="8293" points="834" reactiontime="+87" swimtime="00:01:09.33" resultid="10742" heatid="14243" lane="3" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="656" reactiontime="+85" swimtime="00:01:21.27" resultid="10743" heatid="14274" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="729" reactiontime="+85" swimtime="00:00:31.17" resultid="10744" heatid="14289" lane="4" entrytime="00:00:29.20" />
                <RESULT eventid="8678" points="659" reactiontime="+80" swimtime="00:00:36.30" resultid="10745" heatid="14377" lane="6" entrytime="00:00:37.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-18" firstname="Krystian" gender="M" lastname="Lukaszewicz" nation="POL" athleteid="10750">
              <RESULTS>
                <RESULT eventid="1075" points="594" reactiontime="+84" swimtime="00:00:27.28" resultid="10751" heatid="14155" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="8277" points="583" reactiontime="+100" swimtime="00:01:00.63" resultid="10752" heatid="14233" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="464" reactiontime="+97" swimtime="00:00:31.98" resultid="10753" heatid="14297" lane="2" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-31" firstname="Agnieszka" gender="F" lastname="Dusza-Sabadasz" nation="POL" athleteid="10732">
              <RESULTS>
                <RESULT eventid="1058" points="380" reactiontime="+78" swimtime="00:00:37.52" resultid="10733" heatid="14137" lane="9" entrytime="00:00:38.55" />
                <RESULT eventid="8261" points="335" reactiontime="+103" swimtime="00:01:25.52" resultid="10734" heatid="14219" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-04" firstname="Tomasz" gender="M" lastname="Sabadasz" nation="POL" athleteid="8783">
              <RESULTS>
                <RESULT eventid="1075" points="414" reactiontime="+85" swimtime="00:00:31.87" resultid="8784" heatid="14148" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1105" points="309" reactiontime="+89" swimtime="00:03:09.01" resultid="8785" heatid="14169" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="341" reactiontime="+88" swimtime="00:01:14.51" resultid="8786" heatid="14227" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="311" reactiontime="+92" swimtime="00:01:28.24" resultid="8787" heatid="14247" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="290" reactiontime="+76" swimtime="00:00:37.96" resultid="8788" heatid="14293" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="8518" points="287" reactiontime="+83" swimtime="00:02:51.31" resultid="8789" heatid="14326" lane="9" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:22.65" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-09" firstname="Adam" gender="M" lastname="Marciszonek" nation="POL" athleteid="10802">
              <RESULTS>
                <RESULT eventid="1075" points="627" reactiontime="+77" swimtime="00:00:26.68" resultid="10803" heatid="14156" lane="4" entrytime="00:00:26.50" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10804" heatid="14252" lane="0" entrytime="00:01:10.00" />
                <RESULT eventid="8406" points="592" reactiontime="+79" swimtime="00:01:13.87" resultid="10805" heatid="14283" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="10806" heatid="14388" lane="3" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-05" firstname="Marta" gender="F" lastname="Mazur" nation="POL" athleteid="10766">
              <RESULTS>
                <RESULT eventid="8293" points="411" reactiontime="+94" swimtime="00:01:27.18" resultid="10767" heatid="14241" lane="7" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="399" reactiontime="+94" swimtime="00:01:34.05" resultid="10768" heatid="14272" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="428" reactiontime="+94" swimtime="00:00:37.40" resultid="10769" heatid="14287" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="8678" points="417" reactiontime="+90" swimtime="00:00:41.93" resultid="10770" heatid="14376" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Piotr" gender="M" lastname="Lawniczak" nation="POL" athleteid="10754">
              <RESULTS>
                <RESULT eventid="1075" points="502" reactiontime="+95" swimtime="00:00:28.72" resultid="10755" heatid="14155" lane="0" entrytime="00:00:27.50" />
                <RESULT eventid="8277" points="443" reactiontime="+83" swimtime="00:01:03.71" resultid="10756" heatid="14233" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="424" reactiontime="+91" swimtime="00:00:31.53" resultid="10757" heatid="14297" lane="1" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+77" swimtime="00:02:02.22" resultid="11182" heatid="14267" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="150" swimtime="00:01:30.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10727" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="10780" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="8783" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="9478" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+89" swimtime="00:01:51.47" resultid="11183" heatid="14338" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.88" />
                    <SPLIT distance="100" swimtime="00:00:54.29" />
                    <SPLIT distance="150" swimtime="00:01:25.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10727" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="8783" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9478" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="10780" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+72" swimtime="00:01:59.00" resultid="11184" heatid="14268" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:02.99" />
                    <SPLIT distance="150" swimtime="00:01:32.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10802" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="10754" number="2" reactiontime="+163" />
                    <RELAYPOSITION athleteid="10758" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="10797" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+69" swimtime="00:01:43.72" resultid="11185" heatid="14338" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                    <SPLIT distance="100" swimtime="00:00:54.71" />
                    <SPLIT distance="150" swimtime="00:01:17.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10797" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="9026" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="10802" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="10754" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+70" swimtime="00:01:56.64" resultid="11186" heatid="14268" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="100" swimtime="00:01:04.06" />
                    <SPLIT distance="150" swimtime="00:01:30.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10791" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="10750" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="10771" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="10762" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+72" swimtime="00:01:41.59" resultid="11187" heatid="14339" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                    <SPLIT distance="100" swimtime="00:00:48.25" />
                    <SPLIT distance="150" swimtime="00:01:14.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10771" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="10791" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="10750" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="10762" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+91" swimtime="00:02:26.61" resultid="11180" heatid="14264" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                    <SPLIT distance="150" swimtime="00:01:56.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10741" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="10766" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="10777" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="10746" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8534" reactiontime="+87" swimtime="00:02:10.99" resultid="11181" heatid="14335" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:40.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10746" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="10766" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="10741" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="10732" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="3">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8357" reactiontime="+92" status="DSQ" swimtime="00:02:50.41" resultid="11178" heatid="14264" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:30.06" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10787" number="1" reactiontime="+92" status="DSQ" />
                    <RELAYPOSITION athleteid="10738" number="2" reactiontime="+58" status="DSQ" />
                    <RELAYPOSITION athleteid="10732" number="3" reactiontime="-38" status="DSQ" />
                    <RELAYPOSITION athleteid="10784" number="4" reactiontime="+23" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+79" swimtime="00:02:02.09" resultid="11176" heatid="14392" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:38.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10741" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="10780" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="10746" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="9026" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+64" swimtime="00:01:52.55" resultid="11177" heatid="14177" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.24" />
                    <SPLIT distance="100" swimtime="00:00:55.96" />
                    <SPLIT distance="150" swimtime="00:01:26.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9026" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="10777" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="10746" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="10797" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+75" swimtime="00:02:02.30" resultid="11173" heatid="14176" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                    <SPLIT distance="150" swimtime="00:01:39.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10771" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="10787" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10738" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="10791" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8865" name="Niemaniemogę Sopot">
          <ATHLETES>
            <ATHLETE birthdate="1980-03-02" firstname="Radek" gender="M" lastname="Buszan" nation="POL" athleteid="8866">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="8867" heatid="14154" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="8868" heatid="14232" lane="2" entrytime="00:01:02.00" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="8869" heatid="14329" lane="4" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8765" name="Niezrzeszona Częstochowa">
          <ATHLETES>
            <ATHLETE birthdate="1951-06-06" firstname="Jolanta" gender="F" lastname="Lipińska" nation="POL" athleteid="8766">
              <RESULTS>
                <RESULT eventid="8229" points="132" reactiontime="+121" swimtime="00:06:33.54" resultid="8767" heatid="14208" lane="1" entrytime="00:06:17.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.72" />
                    <SPLIT distance="100" swimtime="00:03:16.73" />
                    <SPLIT distance="150" swimtime="00:04:59.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="78" swimtime="00:03:10.89" resultid="8768" heatid="14238" lane="5" entrytime="00:03:13.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="104" swimtime="00:03:13.70" resultid="8769" heatid="14270" lane="9" entrytime="00:02:55.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="107" reactiontime="+138" swimtime="00:03:04.16" resultid="8770" heatid="14304" lane="0" entrytime="00:02:52.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="126" reactiontime="+73" swimtime="00:06:15.09" resultid="8771" heatid="14362" lane="6" entrytime="00:06:11.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.38" />
                    <SPLIT distance="100" swimtime="00:03:04.39" />
                    <SPLIT distance="150" swimtime="00:04:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="129" swimtime="00:01:21.50" resultid="8772" heatid="14372" lane="5" entrytime="00:01:21.88" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9380" name="Niezrzeszona Kraków">
          <CONTACT name="Joanna Kwatera" />
          <ATHLETES>
            <ATHLETE birthdate="1996-04-04" firstname="Karolina" gender="F" lastname="Szkudlarek" nation="POL" athleteid="9381">
              <RESULTS>
                <RESULT eventid="1058" points="677" reactiontime="+86" swimtime="00:00:29.62" resultid="9382" heatid="14141" lane="2" entrytime="00:00:29.10" />
                <RESULT eventid="1135" points="612" reactiontime="+98" swimtime="00:10:45.06" resultid="9383" heatid="14178" lane="2" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:01:52.17" />
                    <SPLIT distance="200" swimtime="00:02:32.01" />
                    <SPLIT distance="250" swimtime="00:03:12.76" />
                    <SPLIT distance="300" swimtime="00:03:53.12" />
                    <SPLIT distance="350" swimtime="00:04:34.70" />
                    <SPLIT distance="400" swimtime="00:05:16.18" />
                    <SPLIT distance="450" swimtime="00:05:57.53" />
                    <SPLIT distance="500" swimtime="00:06:38.65" />
                    <SPLIT distance="550" swimtime="00:07:20.28" />
                    <SPLIT distance="600" swimtime="00:08:02.48" />
                    <SPLIT distance="650" swimtime="00:08:44.72" />
                    <SPLIT distance="700" swimtime="00:09:26.36" />
                    <SPLIT distance="750" swimtime="00:10:06.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="596" reactiontime="+76" swimtime="00:00:34.78" resultid="9384" heatid="14197" lane="8" entrytime="00:00:33.60" />
                <RESULT eventid="8261" points="737" reactiontime="+84" swimtime="00:01:04.04" resultid="9385" heatid="14223" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="608" reactiontime="+82" swimtime="00:01:15.97" resultid="9386" heatid="14307" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="626" reactiontime="+98" swimtime="00:02:23.97" resultid="9387" heatid="14321" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="529" reactiontime="+78" swimtime="00:02:42.86" resultid="9388" heatid="14365" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:21.14" />
                    <SPLIT distance="150" swimtime="00:02:03.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="573" reactiontime="+77" swimtime="00:05:09.14" resultid="9389" heatid="14393" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="150" swimtime="00:01:52.52" />
                    <SPLIT distance="200" swimtime="00:02:32.03" />
                    <SPLIT distance="250" swimtime="00:03:11.98" />
                    <SPLIT distance="300" swimtime="00:03:52.19" />
                    <SPLIT distance="350" swimtime="00:04:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11408" name="Niezrzeszona Piaseczno">
          <ATHLETES>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="11409">
              <RESULTS>
                <RESULT eventid="1090" points="643" reactiontime="+84" swimtime="00:03:24.48" resultid="11410" heatid="14163" lane="8" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:37.02" />
                    <SPLIT distance="150" swimtime="00:02:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="621" reactiontime="+84" swimtime="00:01:32.67" resultid="11411" heatid="14240" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="599" swimtime="00:01:41.86" resultid="11412" heatid="14271" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="546" reactiontime="+87" swimtime="00:00:40.88" resultid="11413" heatid="14286" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="8678" points="620" reactiontime="+86" swimtime="00:00:45.00" resultid="11414" heatid="14374" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="13206" name="Niezrzeszona Siewierz">
          <ATHLETES>
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="13207">
              <RESULTS>
                <RESULT eventid="1058" points="571" reactiontime="+86" swimtime="00:00:32.75" resultid="13208" heatid="14139" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="8261" points="537" reactiontime="+88" swimtime="00:01:13.11" resultid="13209" heatid="14221" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="493" reactiontime="+97" swimtime="00:01:35.77" resultid="13210" heatid="14272" lane="0" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="425" reactiontime="+79" swimtime="00:00:39.72" resultid="13211" heatid="14287" lane="8" entrytime="00:00:38.30" />
                <RESULT eventid="8678" points="571" reactiontime="+80" swimtime="00:00:41.38" resultid="13212" heatid="14376" lane="0" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8797" name="Niezrzeszona Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1991-02-25" firstname="JOANNA" gender="F" lastname="GRZESZCZUK" nation="POL" athleteid="9009">
              <RESULTS>
                <RESULT eventid="8404" points="775" reactiontime="+71" swimtime="00:01:16.90" resultid="9010" heatid="14274" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="743" reactiontime="+72" swimtime="00:00:30.98" resultid="9011" heatid="14289" lane="7" entrytime="00:00:31.41" />
                <RESULT eventid="8678" points="796" reactiontime="+73" swimtime="00:00:34.08" resultid="9012" heatid="14378" lane="6" entrytime="00:00:34.56" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="8798">
              <RESULTS>
                <RESULT eventid="8261" points="656" reactiontime="+86" swimtime="00:01:08.38" resultid="8799" heatid="14222" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="652" reactiontime="+92" swimtime="00:01:18.56" resultid="8800" heatid="14241" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-04-09" firstname="ANNA" gender="F" lastname="BŁAZUCKA" nation="POL" athleteid="12456">
              <RESULTS>
                <RESULT eventid="1058" points="178" reactiontime="+113" swimtime="00:00:55.07" resultid="12457" heatid="14135" lane="2" entrytime="00:00:52.54" />
                <RESULT eventid="8196" points="117" reactiontime="+97" swimtime="00:01:18.51" resultid="12458" heatid="14193" lane="0" entrytime="00:01:22.15" />
                <RESULT eventid="8293" points="127" reactiontime="+94" swimtime="00:02:37.18" resultid="12459" heatid="14238" lane="4" entrytime="00:02:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="129" reactiontime="+90" swimtime="00:02:49.80" resultid="12460" heatid="14270" lane="0" entrytime="00:02:36.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="180" reactiontime="+113" swimtime="00:04:41.43" resultid="12461" heatid="14317" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.92" />
                    <SPLIT distance="100" swimtime="00:02:15.60" />
                    <SPLIT distance="150" swimtime="00:03:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="155" reactiontime="+82" swimtime="00:01:11.37" resultid="12462" heatid="14372" lane="4" entrytime="00:01:09.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9071" name="Niezrzeszona Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1995-04-25" firstname="Adriana" gender="F" lastname="Hofman" nation="POL" athleteid="9299">
              <RESULTS>
                <RESULT eventid="8404" points="692" reactiontime="+86" swimtime="00:01:19.96" resultid="9300" heatid="14274" lane="2" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="707" reactiontime="+77" swimtime="00:00:36.86" resultid="9301" heatid="14378" lane="7" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-13" firstname="Małgorzata" gender="F" lastname="Bołtuć" nation="POL" athleteid="9072">
              <RESULTS>
                <RESULT eventid="1165" points="451" swimtime="00:24:10.33" resultid="9073" heatid="14187" lane="0" entrytime="00:24:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:17.46" />
                    <SPLIT distance="200" swimtime="00:03:04.72" />
                    <SPLIT distance="250" swimtime="00:03:52.61" />
                    <SPLIT distance="300" swimtime="00:04:41.42" />
                    <SPLIT distance="350" swimtime="00:05:29.88" />
                    <SPLIT distance="400" swimtime="00:06:17.91" />
                    <SPLIT distance="450" swimtime="00:07:06.36" />
                    <SPLIT distance="500" swimtime="00:07:54.65" />
                    <SPLIT distance="550" swimtime="00:08:43.02" />
                    <SPLIT distance="600" swimtime="00:09:31.43" />
                    <SPLIT distance="650" swimtime="00:10:20.12" />
                    <SPLIT distance="700" swimtime="00:11:09.17" />
                    <SPLIT distance="750" swimtime="00:11:57.77" />
                    <SPLIT distance="800" swimtime="00:12:46.49" />
                    <SPLIT distance="850" swimtime="00:13:35.40" />
                    <SPLIT distance="900" swimtime="00:14:24.40" />
                    <SPLIT distance="950" swimtime="00:15:13.19" />
                    <SPLIT distance="1000" swimtime="00:16:02.55" />
                    <SPLIT distance="1050" swimtime="00:16:51.73" />
                    <SPLIT distance="1100" swimtime="00:17:40.59" />
                    <SPLIT distance="1150" swimtime="00:18:29.89" />
                    <SPLIT distance="1200" swimtime="00:19:18.99" />
                    <SPLIT distance="1250" swimtime="00:20:08.07" />
                    <SPLIT distance="1300" swimtime="00:20:56.01" />
                    <SPLIT distance="1350" swimtime="00:21:44.98" />
                    <SPLIT distance="1400" swimtime="00:22:33.94" />
                    <SPLIT distance="1450" swimtime="00:23:22.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="316" swimtime="00:01:24.82" resultid="9074" heatid="14220" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="327" swimtime="00:01:38.25" resultid="9075" heatid="14238" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="328" reactiontime="+127" swimtime="00:01:35.58" resultid="9076" heatid="14305" lane="7" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="351" swimtime="00:03:01.49" resultid="9077" heatid="14319" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:02:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="361" reactiontime="+113" swimtime="00:03:20.54" resultid="9078" heatid="14364" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.65" />
                    <SPLIT distance="100" swimtime="00:01:40.46" />
                    <SPLIT distance="150" swimtime="00:02:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="390" swimtime="00:06:13.69" resultid="9079" heatid="14395" lane="2" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="300" swimtime="00:04:38.35" />
                    <SPLIT distance="350" swimtime="00:05:25.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-25" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="12463">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="12464" heatid="14163" lane="7" entrytime="00:03:31.00" />
                <RESULT eventid="1135" points="346" swimtime="00:13:38.91" resultid="12465" heatid="14180" lane="4" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:32.31" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                    <SPLIT distance="200" swimtime="00:03:16.20" />
                    <SPLIT distance="250" swimtime="00:04:08.38" />
                    <SPLIT distance="300" swimtime="00:04:59.80" />
                    <SPLIT distance="350" swimtime="00:05:52.10" />
                    <SPLIT distance="400" swimtime="00:06:44.39" />
                    <SPLIT distance="450" swimtime="00:07:37.48" />
                    <SPLIT distance="500" swimtime="00:08:29.38" />
                    <SPLIT distance="550" swimtime="00:09:21.82" />
                    <SPLIT distance="600" swimtime="00:10:13.94" />
                    <SPLIT distance="650" swimtime="00:11:07.14" />
                    <SPLIT distance="700" swimtime="00:11:59.31" />
                    <SPLIT distance="750" swimtime="00:12:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="349" reactiontime="+94" swimtime="00:00:43.37" resultid="12466" heatid="14194" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="8293" points="329" reactiontime="+112" swimtime="00:01:38.65" resultid="12467" heatid="14239" lane="3" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="295" reactiontime="+95" swimtime="00:01:41.98" resultid="12468" heatid="14306" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="313" reactiontime="+125" swimtime="00:03:10.36" resultid="12469" heatid="14318" lane="3" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="221" reactiontime="+116" swimtime="00:01:49.28" resultid="12470" heatid="14349" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="301" reactiontime="+64" swimtime="00:03:42.72" resultid="12471" heatid="14364" lane="0" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                    <SPLIT distance="100" swimtime="00:01:49.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9032" name="Niezrzeszony Białystok">
          <ATHLETES>
            <ATHLETE birthdate="1943-01-01" firstname="Edward" gender="M" lastname="DZIEKOŃSKI" nation="POL" athleteid="11154">
              <RESULTS>
                <RESULT eventid="1075" points="411" reactiontime="+124" swimtime="00:00:42.07" resultid="11155" heatid="14145" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1150" points="487" reactiontime="+135" swimtime="00:15:29.75" resultid="11156" heatid="14186" lane="3" entrytime="00:15:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                    <SPLIT distance="100" swimtime="00:01:48.71" />
                    <SPLIT distance="150" swimtime="00:02:46.48" />
                    <SPLIT distance="200" swimtime="00:03:44.11" />
                    <SPLIT distance="250" swimtime="00:04:42.54" />
                    <SPLIT distance="300" swimtime="00:05:41.45" />
                    <SPLIT distance="350" swimtime="00:06:40.99" />
                    <SPLIT distance="400" swimtime="00:07:41.05" />
                    <SPLIT distance="450" swimtime="00:08:39.26" />
                    <SPLIT distance="500" swimtime="00:09:39.38" />
                    <SPLIT distance="550" swimtime="00:10:39.90" />
                    <SPLIT distance="600" swimtime="00:11:39.50" />
                    <SPLIT distance="650" swimtime="00:12:38.14" />
                    <SPLIT distance="700" swimtime="00:13:37.02" />
                    <SPLIT distance="750" swimtime="00:14:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="359" reactiontime="+101" swimtime="00:00:53.31" resultid="11157" heatid="14200" lane="7" entrytime="00:00:51.50" />
                <RESULT eventid="8277" points="453" reactiontime="+119" swimtime="00:01:32.63" resultid="11158" heatid="14225" lane="3" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="409" reactiontime="+129" swimtime="00:00:46.55" resultid="11159" heatid="14292" lane="0" entrytime="00:00:44.50" />
                <RESULT eventid="8486" points="322" reactiontime="+129" swimtime="00:02:01.66" resultid="11160" heatid="14310" lane="8" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="346" reactiontime="+113" swimtime="00:02:01.14" resultid="11161" heatid="14354" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="469" reactiontime="+126" swimtime="00:07:34.27" resultid="11162" heatid="14403" lane="1" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                    <SPLIT distance="100" swimtime="00:01:47.35" />
                    <SPLIT distance="150" swimtime="00:02:45.37" />
                    <SPLIT distance="200" swimtime="00:03:43.87" />
                    <SPLIT distance="250" swimtime="00:04:41.55" />
                    <SPLIT distance="300" swimtime="00:05:39.54" />
                    <SPLIT distance="350" swimtime="00:06:36.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="9033">
              <RESULTS>
                <RESULT eventid="1075" points="822" reactiontime="+80" swimtime="00:00:27.84" resultid="9034" heatid="14154" lane="8" entrytime="00:00:27.95" />
                <RESULT eventid="1105" points="833" reactiontime="+93" swimtime="00:02:34.58" resultid="9035" heatid="14171" lane="4" entrytime="00:02:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                    <SPLIT distance="150" swimtime="00:01:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="843" reactiontime="+81" swimtime="00:01:01.42" resultid="9036" heatid="14232" lane="7" entrytime="00:01:02.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="801" reactiontime="+90" swimtime="00:01:10.82" resultid="9037" heatid="14251" lane="1" entrytime="00:01:11.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="854" reactiontime="+79" swimtime="00:00:30.05" resultid="9038" heatid="14297" lane="9" entrytime="00:00:30.55" />
                <RESULT eventid="8486" points="680" reactiontime="+87" swimtime="00:01:13.62" resultid="9039" heatid="14312" lane="5" entrytime="00:01:15.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="832" reactiontime="+82" swimtime="00:01:08.84" resultid="9040" heatid="14357" lane="3" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="585" reactiontime="+88" swimtime="00:00:36.46" resultid="9041" heatid="14385" lane="1" entrytime="00:00:37.25" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9019" name="Niezrzeszony Bydgoszcz">
          <ATHLETES>
            <ATHLETE birthdate="1978-01-05" firstname="Maciej" gender="M" lastname="Lubas" nation="POL" athleteid="10660">
              <RESULTS>
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="10661" heatid="14216" lane="1" entrytime="00:02:55.00" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10662" heatid="14250" lane="6" entrytime="00:01:14.00" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="10663" heatid="14282" lane="7" entrytime="00:01:18.00" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="10664" heatid="14386" lane="5" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-07" firstname="Michał " gender="M" lastname="Urbański" nation="POL" athleteid="9020">
              <RESULTS>
                <RESULT eventid="8179" points="751" reactiontime="+80" swimtime="00:17:35.07" resultid="9021" heatid="14189" lane="6" entrytime="00:18:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:05.23" />
                    <SPLIT distance="150" swimtime="00:01:39.99" />
                    <SPLIT distance="200" swimtime="00:02:15.10" />
                    <SPLIT distance="250" swimtime="00:02:50.28" />
                    <SPLIT distance="300" swimtime="00:03:25.71" />
                    <SPLIT distance="350" swimtime="00:04:01.19" />
                    <SPLIT distance="400" swimtime="00:04:37.05" />
                    <SPLIT distance="450" swimtime="00:05:12.37" />
                    <SPLIT distance="500" swimtime="00:05:47.59" />
                    <SPLIT distance="550" swimtime="00:06:23.18" />
                    <SPLIT distance="600" swimtime="00:06:58.46" />
                    <SPLIT distance="650" swimtime="00:07:34.08" />
                    <SPLIT distance="700" swimtime="00:08:09.67" />
                    <SPLIT distance="750" swimtime="00:08:45.18" />
                    <SPLIT distance="800" swimtime="00:09:20.69" />
                    <SPLIT distance="850" swimtime="00:09:56.06" />
                    <SPLIT distance="900" swimtime="00:10:31.25" />
                    <SPLIT distance="950" swimtime="00:11:06.72" />
                    <SPLIT distance="1000" swimtime="00:11:42.01" />
                    <SPLIT distance="1050" swimtime="00:12:17.57" />
                    <SPLIT distance="1100" swimtime="00:12:52.79" />
                    <SPLIT distance="1150" swimtime="00:13:28.46" />
                    <SPLIT distance="1200" swimtime="00:14:04.09" />
                    <SPLIT distance="1250" swimtime="00:14:39.12" />
                    <SPLIT distance="1300" swimtime="00:15:14.54" />
                    <SPLIT distance="1350" swimtime="00:15:49.86" />
                    <SPLIT distance="1400" swimtime="00:16:25.43" />
                    <SPLIT distance="1450" swimtime="00:17:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="783" reactiontime="+65" swimtime="00:02:28.69" resultid="9022" heatid="14217" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="9023" heatid="14333" lane="9" entrytime="00:02:05.00" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="9024" heatid="14389" lane="0" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9080" name="Niezrzeszony Gdańsk">
          <ATHLETES>
            <ATHLETE birthdate="1961-01-18" firstname="Wojciech" gender="M" lastname="Warchoł" nation="POL" athleteid="9081">
              <RESULTS>
                <RESULT eventid="8518" points="715" reactiontime="+113" swimtime="00:02:26.54" resultid="9082" heatid="14327" lane="1" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:12.16" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="720" reactiontime="+100" swimtime="00:05:59.99" resultid="9083" heatid="14346" lane="0" entrytime="00:06:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:02:09.24" />
                    <SPLIT distance="200" swimtime="00:02:56.79" />
                    <SPLIT distance="250" swimtime="00:03:48.32" />
                    <SPLIT distance="300" swimtime="00:04:41.30" />
                    <SPLIT distance="350" swimtime="00:05:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="674" reactiontime="+91" swimtime="00:05:23.43" resultid="15631" heatid="14403" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                    <SPLIT distance="200" swimtime="00:02:39.63" />
                    <SPLIT distance="250" swimtime="00:03:20.67" />
                    <SPLIT distance="300" swimtime="00:04:01.84" />
                    <SPLIT distance="350" swimtime="00:04:43.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8870" name="Niezrzeszony Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="8871">
              <RESULTS>
                <RESULT eventid="1105" points="205" reactiontime="+109" swimtime="00:05:01.37" resultid="8872" heatid="14166" lane="4" entrytime="00:05:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.38" />
                    <SPLIT distance="100" swimtime="00:02:24.44" />
                    <SPLIT distance="150" swimtime="00:03:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="190" reactiontime="+105" swimtime="00:05:22.17" resultid="8873" heatid="14212" lane="8" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.12" />
                    <SPLIT distance="100" swimtime="00:02:38.02" />
                    <SPLIT distance="150" swimtime="00:04:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="215" reactiontime="+114" swimtime="00:05:25.60" resultid="8874" heatid="14258" lane="7" entrytime="00:05:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.14" />
                    <SPLIT distance="100" swimtime="00:02:32.41" />
                    <SPLIT distance="150" swimtime="00:04:00.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="212" reactiontime="+109" swimtime="00:00:54.23" resultid="8875" heatid="14291" lane="1" entrytime="00:00:56.00" />
                <RESULT eventid="8518" points="159" reactiontime="+109" swimtime="00:04:37.55" resultid="8876" heatid="14323" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                    <SPLIT distance="100" swimtime="00:02:12.93" />
                    <SPLIT distance="150" swimtime="00:03:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="184" reactiontime="+113" swimtime="00:02:21.89" resultid="8877" heatid="14353" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="169" reactiontime="+116" swimtime="00:10:04.54" resultid="8878" heatid="14404" lane="3" entrytime="00:10:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.76" />
                    <SPLIT distance="100" swimtime="00:02:24.02" />
                    <SPLIT distance="150" swimtime="00:06:20.32" />
                    <SPLIT distance="200" swimtime="00:07:38.10" />
                    <SPLIT distance="250" swimtime="00:08:53.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9121" name="Niezrzeszony Kalisz">
          <ATHLETES>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="9122">
              <RESULTS>
                <RESULT eventid="1075" points="553" reactiontime="+90" swimtime="00:00:32.69" resultid="9123" heatid="14148" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1105" points="637" reactiontime="+83" swimtime="00:03:01.76" resultid="9124" heatid="14169" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:15.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="586" reactiontime="+89" swimtime="00:03:18.21" resultid="9125" heatid="14214" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="100" swimtime="00:01:34.05" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="677" reactiontime="+82" swimtime="00:01:20.71" resultid="9126" heatid="14248" lane="0" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="575" reactiontime="+80" swimtime="00:01:28.80" resultid="9127" heatid="14278" lane="5" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="589" reactiontime="+93" swimtime="00:01:26.10" resultid="9128" heatid="14312" lane="0" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="443" reactiontime="+75" swimtime="00:01:28.40" resultid="9129" heatid="14356" lane="9" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="551" reactiontime="+78" swimtime="00:00:39.92" resultid="9130" heatid="14383" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9646" name="Niezrzeszony Koszalin">
          <ATHLETES>
            <ATHLETE birthdate="1990-11-16" firstname="Dawid" gender="M" lastname="Wróblewski" nation="POL" athleteid="9647">
              <RESULTS>
                <RESULT eventid="1105" points="680" reactiontime="+78" swimtime="00:02:17.05" resultid="9648" heatid="14174" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="765" reactiontime="+82" swimtime="00:02:18.03" resultid="9649" heatid="14262" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="721" reactiontime="+70" swimtime="00:00:26.43" resultid="9650" heatid="14301" lane="1" entrytime="00:00:26.85" />
                <RESULT eventid="8630" points="809" reactiontime="+72" swimtime="00:00:57.87" resultid="9651" heatid="14360" lane="3" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="734" reactiontime="+79" swimtime="00:04:30.94" resultid="9652" heatid="14398" lane="3" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.07" />
                    <SPLIT distance="150" swimtime="00:01:41.14" />
                    <SPLIT distance="200" swimtime="00:02:16.28" />
                    <SPLIT distance="250" swimtime="00:02:51.28" />
                    <SPLIT distance="300" swimtime="00:03:24.97" />
                    <SPLIT distance="350" swimtime="00:03:57.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8892" name="Niezrzeszony Kraków">
          <ATHLETES>
            <ATHLETE birthdate="1938-04-28" firstname="Andrzej" gender="M" lastname="WIŚNIEWSKI" nation="POL" athleteid="8893">
              <RESULTS>
                <RESULT eventid="8179" points="337" swimtime="00:35:20.27" resultid="8894" heatid="14189" lane="7" entrytime="00:35:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                    <SPLIT distance="100" swimtime="00:02:03.47" />
                    <SPLIT distance="150" swimtime="00:03:12.03" />
                    <SPLIT distance="200" swimtime="00:04:20.61" />
                    <SPLIT distance="250" swimtime="00:05:30.06" />
                    <SPLIT distance="300" swimtime="00:06:39.86" />
                    <SPLIT distance="350" swimtime="00:07:49.51" />
                    <SPLIT distance="400" swimtime="00:09:00.03" />
                    <SPLIT distance="450" swimtime="00:10:10.98" />
                    <SPLIT distance="500" swimtime="00:11:21.55" />
                    <SPLIT distance="550" swimtime="00:12:33.85" />
                    <SPLIT distance="600" swimtime="00:13:44.33" />
                    <SPLIT distance="650" swimtime="00:14:55.02" />
                    <SPLIT distance="700" swimtime="00:16:06.26" />
                    <SPLIT distance="750" swimtime="00:17:17.45" />
                    <SPLIT distance="800" swimtime="00:18:29.48" />
                    <SPLIT distance="850" swimtime="00:19:40.80" />
                    <SPLIT distance="900" swimtime="00:20:52.94" />
                    <SPLIT distance="950" swimtime="00:22:05.68" />
                    <SPLIT distance="1000" swimtime="00:23:18.32" />
                    <SPLIT distance="1050" swimtime="00:24:30.15" />
                    <SPLIT distance="1100" swimtime="00:25:41.68" />
                    <SPLIT distance="1150" swimtime="00:26:53.72" />
                    <SPLIT distance="1200" swimtime="00:28:06.22" />
                    <SPLIT distance="1250" swimtime="00:29:18.00" />
                    <SPLIT distance="1300" swimtime="00:30:31.29" />
                    <SPLIT distance="1350" swimtime="00:31:45.11" />
                    <SPLIT distance="1400" swimtime="00:32:57.94" />
                    <SPLIT distance="1450" swimtime="00:34:10.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9370" name="Niezrzeszony Leszno">
          <ATHLETES>
            <ATHLETE birthdate="1985-06-12" firstname="Szymon" gender="M" lastname="Biedny" nation="POL" athleteid="9371">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1105" reactiontime="+66" status="DSQ" swimtime="00:02:30.00" resultid="9372" heatid="14173" lane="5" entrytime="00:02:23.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="150" swimtime="00:01:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="646" reactiontime="+100" swimtime="00:19:08.91" resultid="9373" heatid="14190" lane="4" entrytime="00:19:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:47.00" />
                    <SPLIT distance="200" swimtime="00:02:24.79" />
                    <SPLIT distance="250" swimtime="00:03:03.13" />
                    <SPLIT distance="300" swimtime="00:03:41.69" />
                    <SPLIT distance="350" swimtime="00:04:20.30" />
                    <SPLIT distance="400" swimtime="00:04:58.69" />
                    <SPLIT distance="450" swimtime="00:05:37.13" />
                    <SPLIT distance="500" swimtime="00:06:15.81" />
                    <SPLIT distance="550" swimtime="00:06:54.31" />
                    <SPLIT distance="600" swimtime="00:07:33.07" />
                    <SPLIT distance="650" swimtime="00:08:12.07" />
                    <SPLIT distance="700" swimtime="00:08:50.94" />
                    <SPLIT distance="750" swimtime="00:09:29.50" />
                    <SPLIT distance="800" swimtime="00:10:08.49" />
                    <SPLIT distance="850" swimtime="00:10:47.27" />
                    <SPLIT distance="900" swimtime="00:11:26.55" />
                    <SPLIT distance="950" swimtime="00:12:05.19" />
                    <SPLIT distance="1000" swimtime="00:12:44.09" />
                    <SPLIT distance="1050" swimtime="00:13:23.09" />
                    <SPLIT distance="1100" swimtime="00:14:01.95" />
                    <SPLIT distance="1150" swimtime="00:14:40.49" />
                    <SPLIT distance="1200" swimtime="00:15:19.81" />
                    <SPLIT distance="1250" swimtime="00:15:58.25" />
                    <SPLIT distance="1300" swimtime="00:16:36.97" />
                    <SPLIT distance="1350" swimtime="00:17:15.65" />
                    <SPLIT distance="1400" swimtime="00:17:55.33" />
                    <SPLIT distance="1450" swimtime="00:18:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="489" reactiontime="+89" swimtime="00:01:09.80" resultid="9374" heatid="14252" lane="2" entrytime="00:01:08.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="399" reactiontime="+89" swimtime="00:02:48.47" resultid="9375" heatid="14261" lane="6" entrytime="00:02:32.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="515" reactiontime="+94" swimtime="00:02:12.85" resultid="9376" heatid="14332" lane="2" entrytime="00:02:07.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="545" reactiontime="+119" swimtime="00:05:26.84" resultid="9377" heatid="14347" lane="4" entrytime="00:05:30.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:58.73" />
                    <SPLIT distance="200" swimtime="00:02:41.28" />
                    <SPLIT distance="250" swimtime="00:03:29.57" />
                    <SPLIT distance="300" swimtime="00:04:17.26" />
                    <SPLIT distance="350" swimtime="00:04:53.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="402" reactiontime="+83" swimtime="00:01:11.30" resultid="9378" heatid="14360" lane="8" entrytime="00:01:02.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="610" reactiontime="+80" swimtime="00:04:43.20" resultid="15629" heatid="14399" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:42.38" />
                    <SPLIT distance="200" swimtime="00:02:18.81" />
                    <SPLIT distance="250" swimtime="00:02:55.47" />
                    <SPLIT distance="300" swimtime="00:03:32.64" />
                    <SPLIT distance="350" swimtime="00:04:09.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9366" name="Niezrzeszony Nowy Targ">
          <ATHLETES>
            <ATHLETE birthdate="1992-08-04" firstname="Michał" gender="M" lastname="Starczowski" nation="POL" athleteid="9367">
              <RESULTS>
                <RESULT eventid="1075" points="626" reactiontime="+89" swimtime="00:00:26.70" resultid="9368" heatid="14156" lane="1" entrytime="00:00:26.90" />
                <RESULT eventid="8277" points="528" reactiontime="+84" swimtime="00:01:00.08" resultid="9369" heatid="14232" lane="4" entrytime="00:01:01.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8965" name="Niezrzeszony Olsztyn">
          <ATHLETES>
            <ATHLETE birthdate="1994-03-22" firstname="Sebastian" gender="M" lastname="Borowicz-Skoneczny " nation="POL" athleteid="8966">
              <RESULTS>
                <RESULT eventid="1075" points="629" reactiontime="+73" swimtime="00:00:26.77" resultid="8967" heatid="14156" lane="6" entrytime="00:00:26.63" />
                <RESULT eventid="8277" points="536" reactiontime="+78" swimtime="00:01:02.35" resultid="8968" heatid="14230" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="557" reactiontime="+72" swimtime="00:00:30.08" resultid="8969" heatid="14298" lane="7" entrytime="00:00:29.81" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8879" name="Niezrzeszony Sosnowiec">
          <ATHLETES>
            <ATHLETE birthdate="1941-11-11" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="8880">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="8881" heatid="14167" lane="8" entrytime="00:05:00.00" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="8882" heatid="14186" lane="7" entrytime="00:19:00.00" />
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="8883" heatid="14212" lane="7" entrytime="00:04:55.00" />
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="8884" heatid="14258" lane="8" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="8885" heatid="14324" lane="9" entrytime="00:03:55.00" />
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="8886" heatid="14344" lane="9" />
                <RESULT eventid="8662" status="DNS" swimtime="00:00:00.00" resultid="8887" heatid="14367" lane="8" entrytime="00:04:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8903" name="Niezrzeszony Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1989-02-17" firstname="Piotr" gender="M" lastname="Kister" nation="POL" athleteid="9451">
              <RESULTS>
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="9452" heatid="14215" lane="3" entrytime="00:03:01.00" />
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="9453" heatid="14261" lane="1" entrytime="00:02:45.00" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="9454" heatid="14281" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="9455" heatid="14296" lane="4" entrytime="00:00:30.80" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9456" heatid="14357" lane="6" entrytime="00:01:11.00" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="9457" heatid="14385" lane="4" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-07" firstname="Wieslaw" gender="M" lastname="Bar" nation="POL" athleteid="10822">
              <RESULTS>
                <RESULT eventid="1075" points="623" reactiontime="+89" swimtime="00:00:27.94" resultid="10823" heatid="14153" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="8179" points="583" reactiontime="+91" swimtime="00:19:42.93" resultid="10824" heatid="14190" lane="6" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:48.28" />
                    <SPLIT distance="200" swimtime="00:02:26.59" />
                    <SPLIT distance="250" swimtime="00:03:05.46" />
                    <SPLIT distance="300" swimtime="00:03:44.18" />
                    <SPLIT distance="350" swimtime="00:04:23.55" />
                    <SPLIT distance="400" swimtime="00:05:02.98" />
                    <SPLIT distance="450" swimtime="00:05:42.39" />
                    <SPLIT distance="500" swimtime="00:06:22.24" />
                    <SPLIT distance="550" swimtime="00:07:01.92" />
                    <SPLIT distance="600" swimtime="00:07:42.15" />
                    <SPLIT distance="650" swimtime="00:08:22.16" />
                    <SPLIT distance="700" swimtime="00:09:01.99" />
                    <SPLIT distance="750" swimtime="00:09:41.91" />
                    <SPLIT distance="800" swimtime="00:10:22.21" />
                    <SPLIT distance="850" swimtime="00:11:02.23" />
                    <SPLIT distance="900" swimtime="00:11:42.53" />
                    <SPLIT distance="950" swimtime="00:12:22.84" />
                    <SPLIT distance="1000" swimtime="00:13:02.92" />
                    <SPLIT distance="1050" swimtime="00:13:43.33" />
                    <SPLIT distance="1100" swimtime="00:14:23.80" />
                    <SPLIT distance="1150" swimtime="00:15:04.42" />
                    <SPLIT distance="1200" swimtime="00:15:44.60" />
                    <SPLIT distance="1250" swimtime="00:16:24.75" />
                    <SPLIT distance="1300" swimtime="00:17:05.25" />
                    <SPLIT distance="1350" swimtime="00:17:45.60" />
                    <SPLIT distance="1400" swimtime="00:18:25.96" />
                    <SPLIT distance="1450" swimtime="00:19:06.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="614" reactiontime="+80" swimtime="00:01:02.24" resultid="10825" heatid="14232" lane="9" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="577" reactiontime="+82" swimtime="00:01:12.15" resultid="10826" heatid="14251" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="8518" reactiontime="+73" status="DSQ" swimtime="00:02:15.11" resultid="10827" heatid="14330" lane="6" entrytime="00:02:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                    <SPLIT distance="150" swimtime="00:01:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="581" reactiontime="+100" swimtime="00:04:54.58" resultid="15636" heatid="14403" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="150" swimtime="00:01:43.38" />
                    <SPLIT distance="200" swimtime="00:02:21.39" />
                    <SPLIT distance="250" swimtime="00:02:59.14" />
                    <SPLIT distance="300" swimtime="00:03:38.23" />
                    <SPLIT distance="350" swimtime="00:04:17.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="8904">
              <RESULTS>
                <RESULT eventid="8245" points="417" reactiontime="+113" swimtime="00:03:26.98" resultid="8905" heatid="14214" lane="6" entrytime="00:03:18.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="253" reactiontime="+106" swimtime="00:03:39.46" resultid="8906" heatid="14259" lane="5" entrytime="00:03:33.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:42.69" />
                    <SPLIT distance="150" swimtime="00:02:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="397" reactiontime="+108" swimtime="00:01:34.63" resultid="8907" heatid="14278" lane="3" entrytime="00:01:31.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="8908" heatid="14345" lane="0" entrytime="00:07:25.22" />
                <RESULT eventid="8630" points="272" reactiontime="+99" swimtime="00:01:36.01" resultid="8909" heatid="14355" lane="7" entrytime="00:01:34.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="354" reactiontime="+104" swimtime="00:00:43.47" resultid="8910" heatid="14382" lane="5" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-13" firstname="Dmytro" gender="M" lastname="Bielskyi" nation="POL" athleteid="9005">
              <RESULTS>
                <RESULT eventid="8245" points="509" reactiontime="+86" swimtime="00:02:58.86" resultid="9006" heatid="14215" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:11.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="543" reactiontime="+85" swimtime="00:01:20.42" resultid="9007" heatid="14281" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="346" reactiontime="+95" swimtime="00:02:40.89" resultid="9008" heatid="14326" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:01:59.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11189" name="Niezrzeszony Wołomin">
          <ATHLETES>
            <ATHLETE birthdate="1992-07-23" firstname="Jakub" gender="M" lastname="Jeznach" nation="POL" athleteid="11190">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="11191" heatid="14168" lane="1" entrytime="00:03:50.00" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="11192" heatid="14225" lane="6" entrytime="00:01:35.00" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="11193" heatid="14291" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="11194" heatid="14354" lane="7" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9653" name="Niezrzeszony Wrocław">
          <ATHLETES>
            <ATHLETE birthdate="1998-04-26" firstname="Mateusz" gender="M" lastname="Pinkosz" nation="POL" athleteid="9654">
              <RESULTS>
                <RESULT eventid="1075" points="800" reactiontime="+66" swimtime="00:00:24.71" resultid="9655" heatid="14160" lane="6" entrytime="00:00:24.00" />
                <RESULT eventid="8179" points="742" reactiontime="+68" swimtime="00:17:38.96" resultid="9656" heatid="14189" lane="4" entrytime="00:15:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:37.40" />
                    <SPLIT distance="200" swimtime="00:02:11.90" />
                    <SPLIT distance="250" swimtime="00:02:46.88" />
                    <SPLIT distance="300" swimtime="00:03:21.72" />
                    <SPLIT distance="350" swimtime="00:03:56.52" />
                    <SPLIT distance="400" swimtime="00:04:31.63" />
                    <SPLIT distance="450" swimtime="00:05:06.66" />
                    <SPLIT distance="500" swimtime="00:05:42.13" />
                    <SPLIT distance="550" swimtime="00:06:17.49" />
                    <SPLIT distance="600" swimtime="00:06:52.20" />
                    <SPLIT distance="650" swimtime="00:07:27.36" />
                    <SPLIT distance="700" swimtime="00:08:02.83" />
                    <SPLIT distance="750" swimtime="00:08:38.23" />
                    <SPLIT distance="800" swimtime="00:09:13.90" />
                    <SPLIT distance="850" swimtime="00:09:49.42" />
                    <SPLIT distance="900" swimtime="00:10:25.33" />
                    <SPLIT distance="950" swimtime="00:11:01.30" />
                    <SPLIT distance="1000" swimtime="00:11:37.29" />
                    <SPLIT distance="1050" swimtime="00:12:13.36" />
                    <SPLIT distance="1100" swimtime="00:12:49.69" />
                    <SPLIT distance="1150" swimtime="00:13:25.93" />
                    <SPLIT distance="1200" swimtime="00:14:02.06" />
                    <SPLIT distance="1250" swimtime="00:14:38.47" />
                    <SPLIT distance="1300" swimtime="00:15:15.21" />
                    <SPLIT distance="1350" swimtime="00:15:52.02" />
                    <SPLIT distance="1400" swimtime="00:16:28.30" />
                    <SPLIT distance="1450" swimtime="00:17:04.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="817" reactiontime="+62" swimtime="00:00:54.19" resultid="9657" heatid="14237" lane="6" entrytime="00:00:51.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="735" reactiontime="+76" swimtime="00:02:01.92" resultid="9658" heatid="14333" lane="3" entrytime="00:01:57.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="100" swimtime="00:00:56.79" />
                    <SPLIT distance="150" swimtime="00:01:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="828" reactiontime="+62" swimtime="00:04:21.31" resultid="15635" heatid="14400" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:01:01.01" />
                    <SPLIT distance="150" swimtime="00:01:34.27" />
                    <SPLIT distance="200" swimtime="00:02:08.22" />
                    <SPLIT distance="250" swimtime="00:02:42.55" />
                    <SPLIT distance="300" swimtime="00:03:16.50" />
                    <SPLIT distance="350" swimtime="00:03:50.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9013" name="Niezrzeszony Łódź">
          <ATHLETES>
            <ATHLETE birthdate="1982-05-30" firstname="Łukasz" gender="M" lastname="Bogusiak" nation="POL" athleteid="9014">
              <RESULTS>
                <RESULT eventid="1075" points="205" reactiontime="+95" swimtime="00:00:38.98" resultid="9015" heatid="14147" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="8277" points="214" reactiontime="+83" swimtime="00:01:25.92" resultid="9016" heatid="14227" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="202" reactiontime="+86" swimtime="00:03:09.69" resultid="9017" heatid="14325" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:17.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="13277" name="Ocean’s 7 Inowrocław ">
          <ATHLETES>
            <ATHLETE birthdate="1982-02-27" firstname="Rafał" gender="M" lastname="Domeracki " nation="POL" athleteid="13278">
              <RESULTS>
                <RESULT eventid="8179" points="488" reactiontime="+100" swimtime="00:21:12.21" resultid="13279" heatid="14190" lane="7" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:01:59.87" />
                    <SPLIT distance="200" swimtime="00:02:42.11" />
                    <SPLIT distance="250" swimtime="00:03:24.53" />
                    <SPLIT distance="300" swimtime="00:04:06.98" />
                    <SPLIT distance="350" swimtime="00:04:49.45" />
                    <SPLIT distance="400" swimtime="00:05:31.83" />
                    <SPLIT distance="450" swimtime="00:06:14.72" />
                    <SPLIT distance="500" swimtime="00:06:57.87" />
                    <SPLIT distance="550" swimtime="00:07:40.66" />
                    <SPLIT distance="600" swimtime="00:08:23.54" />
                    <SPLIT distance="650" swimtime="00:09:06.35" />
                    <SPLIT distance="700" swimtime="00:09:49.39" />
                    <SPLIT distance="750" swimtime="00:10:32.51" />
                    <SPLIT distance="800" swimtime="00:11:15.00" />
                    <SPLIT distance="850" swimtime="00:11:57.58" />
                    <SPLIT distance="900" swimtime="00:12:40.28" />
                    <SPLIT distance="950" swimtime="00:13:23.37" />
                    <SPLIT distance="1000" swimtime="00:14:06.87" />
                    <SPLIT distance="1050" swimtime="00:14:50.42" />
                    <SPLIT distance="1100" swimtime="00:15:33.21" />
                    <SPLIT distance="1150" swimtime="00:16:16.41" />
                    <SPLIT distance="1200" swimtime="00:16:58.83" />
                    <SPLIT distance="1250" swimtime="00:17:41.74" />
                    <SPLIT distance="1300" swimtime="00:18:24.69" />
                    <SPLIT distance="1350" swimtime="00:19:07.51" />
                    <SPLIT distance="1400" swimtime="00:19:50.22" />
                    <SPLIT distance="1450" swimtime="00:20:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LAT" clubid="9959" name="PK CHAMPIONS Rīga">
          <ATHLETES>
            <ATHLETE birthdate="1974-05-17" firstname="Aiga" gender="F" lastname="Skabe" nation="LAT" athleteid="9968">
              <RESULTS>
                <RESULT eventid="1135" points="404" reactiontime="+106" swimtime="00:12:57.66" resultid="9969" heatid="14179" lane="2" entrytime="00:13:11.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:01:26.26" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                    <SPLIT distance="200" swimtime="00:03:03.73" />
                    <SPLIT distance="250" swimtime="00:03:52.97" />
                    <SPLIT distance="300" swimtime="00:04:42.31" />
                    <SPLIT distance="350" swimtime="00:05:32.38" />
                    <SPLIT distance="400" swimtime="00:06:22.47" />
                    <SPLIT distance="450" swimtime="00:07:12.26" />
                    <SPLIT distance="500" swimtime="00:08:02.15" />
                    <SPLIT distance="550" swimtime="00:08:52.07" />
                    <SPLIT distance="600" swimtime="00:09:42.21" />
                    <SPLIT distance="650" swimtime="00:10:32.26" />
                    <SPLIT distance="700" swimtime="00:11:22.15" />
                    <SPLIT distance="750" swimtime="00:12:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="484" reactiontime="+82" swimtime="00:03:31.51" resultid="9970" heatid="14210" lane="7" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                    <SPLIT distance="150" swimtime="00:02:35.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-02-07" firstname="Edgars" gender="M" lastname="Ozolins" nation="POL" athleteid="9960">
              <RESULTS>
                <RESULT eventid="8277" points="937" reactiontime="+91" swimtime="00:00:59.29" resultid="9961" heatid="14234" lane="0" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="954" reactiontime="+94" swimtime="00:02:13.08" resultid="9962" heatid="14330" lane="5" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.78" />
                    <SPLIT distance="150" swimtime="00:01:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="827" reactiontime="+85" swimtime="00:02:34.95" resultid="9963" heatid="14170" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:13.90" />
                    <SPLIT distance="150" swimtime="00:02:00.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-15" firstname="Andrejs" gender="M" lastname="Sibircevs" nation="LAT" athleteid="9964">
              <RESULTS>
                <RESULT eventid="1075" points="339" reactiontime="+80" swimtime="00:00:32.98" resultid="9965" heatid="14148" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="8277" points="337" reactiontime="+81" swimtime="00:01:13.87" resultid="9966" heatid="14227" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="309" reactiontime="+96" swimtime="00:02:44.86" resultid="9967" heatid="14326" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:01.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="8911" name="PK Zabreh">
          <ATHLETES>
            <ATHLETE birthdate="1973-09-19" firstname="Jiri" gender="M" lastname="Sip" nation="CZE" athleteid="8912">
              <RESULTS>
                <RESULT eventid="1075" points="710" reactiontime="+92" swimtime="00:00:26.75" resultid="8913" heatid="14155" lane="3" entrytime="00:00:27.10" />
                <RESULT eventid="1105" points="780" reactiontime="+96" swimtime="00:02:26.96" resultid="8914" heatid="14172" lane="4" entrytime="00:02:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="686" reactiontime="+86" swimtime="00:00:31.59" resultid="8915" heatid="14205" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="8277" points="735" reactiontime="+90" swimtime="00:00:58.63" resultid="8916" heatid="14234" lane="9" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="633" reactiontime="+89" swimtime="00:01:16.93" resultid="8917" heatid="14282" lane="9" entrytime="00:01:19.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="685" reactiontime="+91" swimtime="00:01:07.45" resultid="8918" heatid="14314" lane="0" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="750" reactiontime="+79" swimtime="00:02:29.96" resultid="8919" heatid="14370" lane="6" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-02" firstname="Jakub" gender="M" lastname="Smid" nation="CZE" athleteid="8920">
              <RESULTS>
                <RESULT eventid="1075" points="682" reactiontime="+89" swimtime="00:00:26.06" resultid="8921" heatid="14158" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1105" points="612" reactiontime="+77" swimtime="00:02:29.55" resultid="8922" heatid="14174" lane="9" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:06.56" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="695" reactiontime="+86" swimtime="00:00:57.18" resultid="8923" heatid="14236" lane="1" entrytime="00:00:56.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="684" reactiontime="+73" swimtime="00:01:03.79" resultid="8924" heatid="14254" lane="8" entrytime="00:01:04.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="723" reactiontime="+87" swimtime="00:01:08.76" resultid="8925" heatid="14283" lane="4" entrytime="00:01:08.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="664" reactiontime="+80" swimtime="00:00:28.38" resultid="8926" heatid="14299" lane="6" entrytime="00:00:28.53" />
                <RESULT eventid="8694" points="745" reactiontime="+76" swimtime="00:00:31.17" resultid="8927" heatid="14388" lane="5" entrytime="00:00:31.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-26" firstname="David" gender="M" lastname="Kochwasser" nation="CZE" athleteid="9114">
              <RESULTS>
                <RESULT eventid="1075" points="506" reactiontime="+77" swimtime="00:00:28.77" resultid="9115" heatid="14152" lane="4" entrytime="00:00:28.87" />
                <RESULT eventid="8277" points="498" reactiontime="+74" swimtime="00:01:03.88" resultid="9116" heatid="14230" lane="7" entrytime="00:01:05.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="498" reactiontime="+78" swimtime="00:01:17.86" resultid="9117" heatid="14281" lane="7" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="441" reactiontime="+83" swimtime="00:05:52.26" resultid="9118" heatid="14346" lane="8" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:06.11" />
                    <SPLIT distance="200" swimtime="00:02:53.49" />
                    <SPLIT distance="250" swimtime="00:03:41.74" />
                    <SPLIT distance="300" swimtime="00:04:30.98" />
                    <SPLIT distance="350" swimtime="00:05:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="8630" reactiontime="+93" status="DSQ" swimtime="00:01:12.60" resultid="9119" heatid="14357" lane="8" entrytime="00:01:14.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="548" reactiontime="+75" swimtime="00:00:34.53" resultid="9120" heatid="14386" lane="4" entrytime="00:00:35.25" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="11691" name="Pregel Kaliningrad">
          <CONTACT city="Kaliningrad" email="alkonter@gmail.com" name="Pregel" phone="+79062384111" street="Turgeneva 5-9" zip="236008" />
          <ATHLETES>
            <ATHLETE birthdate="1946-11-10" firstname="Vyacheslav" gender="M" lastname="Tikhonov" nation="RUS" athleteid="11734">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="11735" heatid="14146" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="11736" heatid="14201" lane="0" entrytime="00:00:45.50" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="11737" heatid="14226" lane="7" entrytime="00:01:24.50" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="11738" heatid="14292" lane="9" entrytime="00:00:44.50" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="11739" heatid="14381" lane="5" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-20" firstname="ALeksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="11753">
              <RESULTS>
                <RESULT eventid="1075" points="509" reactiontime="+95" swimtime="00:00:33.61" resultid="11754" heatid="14146" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="8213" points="365" reactiontime="+82" swimtime="00:00:44.46" resultid="11755" heatid="14201" lane="7" entrytime="00:00:43.50" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="11756" heatid="14277" lane="6" entrytime="00:01:43.50" />
                <RESULT eventid="8694" points="481" reactiontime="+90" swimtime="00:00:41.77" resultid="11757" heatid="14382" lane="1" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-06" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="11698">
              <RESULTS>
                <RESULT eventid="1058" points="631" swimtime="00:00:34.48" resultid="11699" heatid="14137" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="8196" points="582" reactiontime="+90" swimtime="00:00:43.22" resultid="11700" heatid="14195" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="8261" points="626" reactiontime="+95" swimtime="00:01:14.94" resultid="11701" heatid="14220" lane="4" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="608" swimtime="00:02:43.25" resultid="11702" heatid="14320" lane="7" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="628" swimtime="00:05:44.28" resultid="15637" heatid="14396" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-08-21" firstname="Grigorii" gender="M" lastname="Lopin" nation="RUS" athleteid="11764">
              <RESULTS>
                <RESULT eventid="1075" points="601" reactiontime="+91" swimtime="00:00:30.89" resultid="11765" heatid="14149" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1150" points="545" reactiontime="+110" swimtime="00:12:00.58" resultid="11766" heatid="14184" lane="0" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="200" swimtime="00:02:48.08" />
                    <SPLIT distance="250" swimtime="00:03:33.44" />
                    <SPLIT distance="300" swimtime="00:04:19.38" />
                    <SPLIT distance="350" swimtime="00:05:05.44" />
                    <SPLIT distance="400" swimtime="00:05:50.50" />
                    <SPLIT distance="450" swimtime="00:06:36.15" />
                    <SPLIT distance="500" swimtime="00:07:22.84" />
                    <SPLIT distance="550" swimtime="00:08:09.10" />
                    <SPLIT distance="600" swimtime="00:08:55.62" />
                    <SPLIT distance="650" swimtime="00:09:42.39" />
                    <SPLIT distance="700" swimtime="00:10:29.26" />
                    <SPLIT distance="750" swimtime="00:11:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="592" reactiontime="+103" swimtime="00:03:12.91" resultid="11767" heatid="14214" lane="3" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                    <SPLIT distance="150" swimtime="00:02:21.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="494" reactiontime="+99" swimtime="00:01:26.18" resultid="11768" heatid="14279" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="547" reactiontime="+93" swimtime="00:06:34.45" resultid="11769" heatid="14345" lane="5" entrytime="00:06:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:37.77" />
                    <SPLIT distance="150" swimtime="00:02:30.40" />
                    <SPLIT distance="200" swimtime="00:03:24.11" />
                    <SPLIT distance="250" swimtime="00:04:16.77" />
                    <SPLIT distance="300" swimtime="00:05:10.43" />
                    <SPLIT distance="350" swimtime="00:05:53.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="475" reactiontime="+90" swimtime="00:00:39.09" resultid="11770" heatid="14384" lane="9" entrytime="00:00:39.50" />
                <RESULT eventid="8742" points="552" reactiontime="+93" swimtime="00:05:45.64" resultid="11771" heatid="14401" lane="0" entrytime="00:05:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:20.53" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                    <SPLIT distance="200" swimtime="00:02:49.19" />
                    <SPLIT distance="250" swimtime="00:03:34.15" />
                    <SPLIT distance="300" swimtime="00:04:18.45" />
                    <SPLIT distance="350" swimtime="00:05:02.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-02-11" firstname="Nadezhda" gender="F" lastname="Davydova" nation="RUS" athleteid="11704">
              <RESULTS>
                <RESULT eventid="1090" points="550" reactiontime="+109" swimtime="00:03:09.50" resultid="11705" heatid="14163" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:02:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="561" reactiontime="+93" swimtime="00:01:26.86" resultid="11706" heatid="14240" lane="5" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="524" reactiontime="+99" swimtime="00:00:38.62" resultid="11707" heatid="14286" lane="4" entrytime="00:00:40.50" />
                <RESULT eventid="8502" points="518" reactiontime="+86" swimtime="00:02:47.84" resultid="11708" heatid="14319" lane="7" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="487" reactiontime="+98" swimtime="00:00:46.38" resultid="11709" heatid="14375" lane="1" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-04-17" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="11772">
              <RESULTS>
                <RESULT eventid="1075" points="572" reactiontime="+76" swimtime="00:00:30.60" resultid="11773" heatid="14149" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="1150" points="540" reactiontime="+69" swimtime="00:10:59.94" resultid="11774" heatid="14183" lane="8" entrytime="00:11:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                    <SPLIT distance="150" swimtime="00:02:00.34" />
                    <SPLIT distance="200" swimtime="00:02:42.51" />
                    <SPLIT distance="250" swimtime="00:03:24.65" />
                    <SPLIT distance="300" swimtime="00:04:07.29" />
                    <SPLIT distance="350" swimtime="00:04:50.09" />
                    <SPLIT distance="400" swimtime="00:05:32.62" />
                    <SPLIT distance="450" swimtime="00:06:14.53" />
                    <SPLIT distance="500" swimtime="00:06:56.48" />
                    <SPLIT distance="550" swimtime="00:07:38.17" />
                    <SPLIT distance="600" swimtime="00:08:19.98" />
                    <SPLIT distance="650" swimtime="00:09:01.55" />
                    <SPLIT distance="700" swimtime="00:09:42.29" />
                    <SPLIT distance="750" swimtime="00:10:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="571" reactiontime="+77" swimtime="00:01:08.02" resultid="11775" heatid="14229" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="616" reactiontime="+73" swimtime="00:01:16.54" resultid="11776" heatid="14249" lane="2" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="614" reactiontime="+63" swimtime="00:01:21.81" resultid="11777" heatid="14281" lane="9" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="592" reactiontime="+70" swimtime="00:02:28.31" resultid="11778" heatid="14328" lane="7" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="601" reactiontime="+66" swimtime="00:00:36.44" resultid="11779" heatid="14385" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="8742" points="557" reactiontime="+66" swimtime="00:05:16.53" resultid="11780" heatid="14401" lane="4" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                    <SPLIT distance="200" swimtime="00:02:39.50" />
                    <SPLIT distance="250" swimtime="00:03:19.39" />
                    <SPLIT distance="300" swimtime="00:03:59.05" />
                    <SPLIT distance="350" swimtime="00:04:38.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-06-27" firstname="Vladimir" gender="M" lastname="Getman" nation="RUS" athleteid="11745">
              <RESULTS>
                <RESULT eventid="1075" points="800" reactiontime="+77" swimtime="00:00:29.71" resultid="11746" heatid="14150" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1105" points="806" reactiontime="+96" swimtime="00:02:53.64" resultid="11747" heatid="14170" lane="0" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="150" swimtime="00:02:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="947" reactiontime="+80" swimtime="00:03:05.46" resultid="11748" heatid="14214" lane="5" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:18.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="861" reactiontime="+76" swimtime="00:01:17.67" resultid="11749" heatid="14249" lane="7" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="903" reactiontime="+87" swimtime="00:01:22.14" resultid="11750" heatid="14280" lane="4" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="813" reactiontime="+106" swimtime="00:06:34.49" resultid="11751" heatid="14346" lane="2" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                    <SPLIT distance="100" swimtime="00:01:33.81" />
                    <SPLIT distance="150" swimtime="00:02:29.18" />
                    <SPLIT distance="200" swimtime="00:03:23.70" />
                    <SPLIT distance="250" swimtime="00:04:13.88" />
                    <SPLIT distance="300" swimtime="00:05:06.13" />
                    <SPLIT distance="350" swimtime="00:05:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="836" reactiontime="+71" swimtime="00:00:37.03" resultid="11752" heatid="14385" lane="8" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-09-19" firstname="Sergei" gender="M" lastname="Mikhaylov" nation="RUS" athleteid="11758">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="11759" heatid="14145" lane="7" entrytime="00:00:39.50" />
                <RESULT eventid="8179" status="DNS" swimtime="00:00:00.00" resultid="11760" heatid="14192" lane="3" entrytime="00:26:59.00" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="11761" heatid="14225" lane="4" entrytime="00:01:28.50" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="11762" heatid="14324" lane="4" entrytime="00:03:12.00" />
                <RESULT eventid="8742" points="417" reactiontime="+81" swimtime="00:06:19.51" resultid="11763" heatid="14402" lane="8" entrytime="00:06:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:31.68" />
                    <SPLIT distance="150" swimtime="00:02:20.84" />
                    <SPLIT distance="200" swimtime="00:03:09.41" />
                    <SPLIT distance="250" swimtime="00:03:57.11" />
                    <SPLIT distance="300" swimtime="00:04:44.84" />
                    <SPLIT distance="350" swimtime="00:05:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-25" firstname="Elena" gender="F" lastname="Dautova" nation="RUS" athleteid="11710">
              <RESULTS>
                <RESULT eventid="1058" points="661" reactiontime="+86" swimtime="00:00:31.35" resultid="11711" heatid="14139" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="8196" points="552" reactiontime="+86" swimtime="00:00:37.58" resultid="11712" heatid="14196" lane="1" entrytime="00:00:38.50" />
                <RESULT eventid="8261" points="562" reactiontime="+78" swimtime="00:01:12.23" resultid="11713" heatid="14221" lane="4" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="531" reactiontime="+73" swimtime="00:01:26.41" resultid="11714" heatid="14306" lane="8" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="561" reactiontime="+84" swimtime="00:00:42.63" resultid="11715" heatid="14375" lane="6" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-05-10" firstname="Yuri" gender="M" lastname="Yakovenko" nation="RUS" athleteid="11740">
              <RESULTS>
                <RESULT eventid="1075" points="379" reactiontime="+118" swimtime="00:00:38.11" resultid="11741" heatid="14145" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="8245" points="454" reactiontime="+109" swimtime="00:03:56.97" resultid="11742" heatid="14213" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.51" />
                    <SPLIT distance="100" swimtime="00:01:51.63" />
                    <SPLIT distance="150" swimtime="00:02:55.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="423" reactiontime="+112" swimtime="00:01:45.76" resultid="11743" heatid="14277" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="469" reactiontime="+102" swimtime="00:00:44.88" resultid="11744" heatid="14381" lane="4" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-24" firstname="Vitalii" gender="M" lastname="Avdeev" nation="RUS" athleteid="11726">
              <RESULTS>
                <RESULT eventid="1105" points="393" reactiontime="+112" swimtime="00:03:40.56" resultid="11727" heatid="14168" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:53.96" />
                    <SPLIT distance="150" swimtime="00:02:55.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="719" reactiontime="+111" swimtime="00:24:34.22" resultid="11728" heatid="14191" lane="2" entrytime="00:26:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:16.20" />
                    <SPLIT distance="200" swimtime="00:03:05.29" />
                    <SPLIT distance="250" swimtime="00:03:54.15" />
                    <SPLIT distance="300" swimtime="00:04:43.51" />
                    <SPLIT distance="350" swimtime="00:05:33.61" />
                    <SPLIT distance="400" swimtime="00:06:22.79" />
                    <SPLIT distance="450" swimtime="00:07:11.78" />
                    <SPLIT distance="500" swimtime="00:08:00.70" />
                    <SPLIT distance="550" swimtime="00:08:49.99" />
                    <SPLIT distance="600" swimtime="00:09:39.33" />
                    <SPLIT distance="650" swimtime="00:10:27.60" />
                    <SPLIT distance="700" swimtime="00:11:17.54" />
                    <SPLIT distance="750" swimtime="00:12:06.97" />
                    <SPLIT distance="800" swimtime="00:12:57.08" />
                    <SPLIT distance="850" swimtime="00:13:46.99" />
                    <SPLIT distance="900" swimtime="00:14:36.46" />
                    <SPLIT distance="950" swimtime="00:15:25.18" />
                    <SPLIT distance="1000" swimtime="00:16:15.46" />
                    <SPLIT distance="1050" swimtime="00:17:05.75" />
                    <SPLIT distance="1100" swimtime="00:17:55.15" />
                    <SPLIT distance="1150" swimtime="00:18:44.52" />
                    <SPLIT distance="1200" swimtime="00:19:35.11" />
                    <SPLIT distance="1250" swimtime="00:20:25.69" />
                    <SPLIT distance="1300" swimtime="00:21:16.04" />
                    <SPLIT distance="1350" swimtime="00:22:05.99" />
                    <SPLIT distance="1400" swimtime="00:22:56.56" />
                    <SPLIT distance="1450" swimtime="00:23:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="447" reactiontime="+109" swimtime="00:01:36.62" resultid="11729" heatid="14246" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="421" reactiontime="+109" swimtime="00:03:43.22" resultid="11730" heatid="14259" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                    <SPLIT distance="100" swimtime="00:01:44.42" />
                    <SPLIT distance="150" swimtime="00:02:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="524" reactiontime="+121" swimtime="00:00:37.90" resultid="11731" heatid="14294" lane="3" entrytime="00:00:39.50" />
                <RESULT eventid="8518" points="514" reactiontime="+87" swimtime="00:02:58.17" resultid="11732" heatid="14325" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                    <SPLIT distance="150" swimtime="00:02:13.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="11733" heatid="14355" lane="8" entrytime="00:01:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-20" firstname="Sergei" gender="M" lastname="Karakchiev" nation="RUS" athleteid="11783">
              <RESULTS>
                <RESULT eventid="1075" points="773" reactiontime="+84" swimtime="00:00:27.68" resultid="11784" heatid="14153" lane="5" entrytime="00:00:28.00" />
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach." eventid="8213" reactiontime="+87" status="DSQ" swimtime="00:00:32.92" resultid="11785" heatid="14205" lane="9" entrytime="00:00:32.80" />
                <RESULT eventid="8309" points="862" reactiontime="+84" swimtime="00:01:08.44" resultid="11786" heatid="14252" lane="1" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="750" reactiontime="+101" swimtime="00:01:10.03" resultid="11787" heatid="14313" lane="5" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" status="DNS" swimtime="00:00:00.00" resultid="11788" heatid="14370" lane="0" entrytime="00:02:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-01" firstname="Elena" gender="F" lastname="Kolyadina" nation="RUS" athleteid="11692">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="11693" heatid="14137" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="8229" status="DNS" swimtime="00:00:00.00" resultid="11694" heatid="14210" lane="9" entrytime="00:03:37.00" />
                <RESULT eventid="8293" status="DNS" swimtime="00:00:00.00" resultid="11695" heatid="14240" lane="2" entrytime="00:01:31.50" />
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="11696" heatid="14272" lane="1" entrytime="00:01:37.50" />
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="11697" heatid="14375" lane="0" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-26" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="11781">
              <RESULTS>
                <RESULT eventid="8179" points="606" reactiontime="+90" swimtime="00:20:02.02" resultid="11782" heatid="14190" lane="5" entrytime="00:19:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:13.75" />
                    <SPLIT distance="150" swimtime="00:01:53.47" />
                    <SPLIT distance="200" swimtime="00:02:33.56" />
                    <SPLIT distance="250" swimtime="00:03:13.63" />
                    <SPLIT distance="300" swimtime="00:03:53.38" />
                    <SPLIT distance="350" swimtime="00:04:32.72" />
                    <SPLIT distance="400" swimtime="00:05:12.62" />
                    <SPLIT distance="450" swimtime="00:05:52.57" />
                    <SPLIT distance="500" swimtime="00:06:32.73" />
                    <SPLIT distance="550" swimtime="00:07:12.73" />
                    <SPLIT distance="600" swimtime="00:07:53.13" />
                    <SPLIT distance="650" swimtime="00:08:33.75" />
                    <SPLIT distance="700" swimtime="00:09:14.01" />
                    <SPLIT distance="750" swimtime="00:09:54.41" />
                    <SPLIT distance="800" swimtime="00:10:34.96" />
                    <SPLIT distance="850" swimtime="00:11:15.75" />
                    <SPLIT distance="900" swimtime="00:11:56.63" />
                    <SPLIT distance="950" swimtime="00:12:38.02" />
                    <SPLIT distance="1000" swimtime="00:13:18.50" />
                    <SPLIT distance="1050" swimtime="00:13:58.83" />
                    <SPLIT distance="1100" swimtime="00:14:40.21" />
                    <SPLIT distance="1150" swimtime="00:15:20.92" />
                    <SPLIT distance="1200" swimtime="00:16:01.03" />
                    <SPLIT distance="1250" swimtime="00:16:41.72" />
                    <SPLIT distance="1300" swimtime="00:17:22.70" />
                    <SPLIT distance="1350" swimtime="00:18:03.35" />
                    <SPLIT distance="1400" swimtime="00:18:44.22" />
                    <SPLIT distance="1450" swimtime="00:19:24.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-07-21" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="11721">
              <RESULTS>
                <RESULT eventid="1058" points="942" reactiontime="+85" swimtime="00:00:26.66" resultid="11722" heatid="14141" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="8196" points="792" reactiontime="+82" swimtime="00:00:32.81" resultid="11723" heatid="14197" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="8261" points="959" reactiontime="+85" swimtime="00:00:58.27" resultid="11724" heatid="14223" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="917" reactiontime="+84" swimtime="00:00:29.01" resultid="11725" heatid="14289" lane="3" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+84" swimtime="00:02:21.96" resultid="11795" heatid="14266" lane="0" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:10.50" />
                    <SPLIT distance="150" swimtime="00:01:48.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11783" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="11745" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="11726" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="11753" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" swimtime="00:02:07.57" resultid="11796" heatid="14337" lane="8" entrytime="00:02:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="150" swimtime="00:01:31.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11783" number="1" />
                    <RELAYPOSITION athleteid="11745" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="11753" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="11726" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT comment="S3 - Pływacy przepłynęli wyścig w kolejności niezgodnej ze zgłoszeniem." eventid="8357" reactiontime="+69" status="DSQ" swimtime="00:02:30.27" resultid="11793" heatid="14264" lane="9" entrytime="00:02:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:01:55.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11710" number="1" reactiontime="+69" status="DSQ" />
                    <RELAYPOSITION athleteid="11692" number="2" reactiontime="+59" status="DSQ" />
                    <RELAYPOSITION athleteid="11704" number="3" reactiontime="+54" status="DSQ" />
                    <RELAYPOSITION athleteid="11698" number="4" reactiontime="+43" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S3 - Pływacy przepłynęli wyścig w kolejności niezgodnej ze zgłoszeniem." eventid="8534" reactiontime="+90" status="DSQ" swimtime="00:02:06.14" resultid="11794" heatid="14335" lane="9" entrytime="00:02:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:31.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11698" number="1" reactiontime="+90" status="DSQ" />
                    <RELAYPOSITION athleteid="11692" number="2" reactiontime="+52" status="DSQ" />
                    <RELAYPOSITION athleteid="11721" number="3" reactiontime="+40" status="DSQ" />
                    <RELAYPOSITION athleteid="11704" number="4" reactiontime="+52" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S3 - Pływacy przepłynęli wyścig w kolejności niezgodnej ze zgłoszeniem." eventid="1120" reactiontime="+107" status="DSQ" swimtime="00:02:17.13" resultid="11789" heatid="14175" lane="5" entrytime="00:02:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                    <SPLIT distance="150" swimtime="00:01:40.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11753" number="1" reactiontime="+107" status="DSQ" />
                    <RELAYPOSITION athleteid="11704" number="2" reactiontime="+45" status="DSQ" />
                    <RELAYPOSITION athleteid="11692" number="3" reactiontime="+34" status="DSQ" />
                    <RELAYPOSITION athleteid="11726" number="4" reactiontime="+58" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+67" swimtime="00:02:23.60" resultid="11790" heatid="14392" lane="6" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:49.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11710" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="11745" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="11772" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="11704" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+79" swimtime="00:01:58.83" resultid="11792" heatid="14176" lane="7" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="150" swimtime="00:01:25.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11783" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="11745" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="11721" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="11698" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9486" name="RakTeam">
          <ATHLETES>
            <ATHLETE birthdate="1989-07-05" firstname="Maja " gender="F" lastname="Spychalska" nation="POL" athleteid="9487">
              <RESULTS>
                <RESULT eventid="1058" points="654" reactiontime="+82" swimtime="00:00:29.66" resultid="9488" heatid="14141" lane="9" entrytime="00:00:29.90" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="9489" heatid="14223" lane="9" entrytime="00:01:07.00" />
                <RESULT eventid="8404" points="642" reactiontime="+99" swimtime="00:01:21.86" resultid="9490" heatid="14273" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="661" reactiontime="+84" swimtime="00:00:36.25" resultid="9491" heatid="14377" lane="4" entrytime="00:00:36.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-15" firstname="Mateusz " gender="M" lastname="Rak" nation="POL" athleteid="9492">
              <RESULTS>
                <RESULT eventid="8179" status="DNS" swimtime="00:00:00.00" resultid="9493" heatid="14192" lane="4" entrytime="00:18:45.00" />
                <RESULT eventid="8213" points="737" reactiontime="+69" swimtime="00:00:27.73" resultid="9494" heatid="14207" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="8486" points="805" reactiontime="+77" swimtime="00:00:59.15" resultid="9495" heatid="14315" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="736" reactiontime="+69" swimtime="00:02:08.70" resultid="9496" heatid="14371" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8801" name="Rydułtowska AAS">
          <CONTACT name="MARIAN OTLIK" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="8809">
              <RESULTS>
                <RESULT eventid="1075" points="77" reactiontime="+99" swimtime="00:01:13.56" resultid="8810" heatid="14142" lane="3" />
                <RESULT eventid="8213" points="50" reactiontime="+121" swimtime="00:01:42.42" resultid="8811" heatid="14198" lane="5" />
                <RESULT eventid="8277" points="97" reactiontime="+106" swimtime="00:02:34.62" resultid="8812" heatid="14224" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="59" reactiontime="+189" swimtime="00:03:33.96" resultid="8813" heatid="14308" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="106" reactiontime="+139" swimtime="00:05:35.18" resultid="8814" heatid="14322" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.21" />
                    <SPLIT distance="100" swimtime="00:02:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="81" reactiontime="+81" swimtime="00:07:35.93" resultid="8815" heatid="14366" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="121" reactiontime="+121" swimtime="00:11:53.79" resultid="8816" heatid="14404" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.31" />
                    <SPLIT distance="100" swimtime="00:02:36.53" />
                    <SPLIT distance="150" swimtime="00:04:05.97" />
                    <SPLIT distance="200" swimtime="00:05:37.35" />
                    <SPLIT distance="250" swimtime="00:07:07.92" />
                    <SPLIT distance="300" swimtime="00:08:42.00" />
                    <SPLIT distance="350" swimtime="00:10:19.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="8834">
              <RESULTS>
                <RESULT comment="K13 - Pływak nie zwrócił stóp na zewnątrz w trakcie napędzającej części ruchu nóg." eventid="1105" reactiontime="+71" status="DSQ" swimtime="00:03:18.30" resultid="8835" heatid="14169" lane="9" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="150" swimtime="00:02:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="685" reactiontime="+106" swimtime="00:24:57.96" resultid="8836" heatid="14191" lane="3" entrytime="00:25:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:17.76" />
                    <SPLIT distance="200" swimtime="00:03:07.05" />
                    <SPLIT distance="250" swimtime="00:03:56.33" />
                    <SPLIT distance="300" swimtime="00:04:45.92" />
                    <SPLIT distance="350" swimtime="00:05:35.88" />
                    <SPLIT distance="400" swimtime="00:06:25.91" />
                    <SPLIT distance="450" swimtime="00:07:15.24" />
                    <SPLIT distance="500" swimtime="00:08:05.43" />
                    <SPLIT distance="550" swimtime="00:08:55.55" />
                    <SPLIT distance="600" swimtime="00:09:45.90" />
                    <SPLIT distance="650" swimtime="00:10:36.90" />
                    <SPLIT distance="700" swimtime="00:11:27.94" />
                    <SPLIT distance="750" swimtime="00:12:18.70" />
                    <SPLIT distance="800" swimtime="00:13:09.40" />
                    <SPLIT distance="850" swimtime="00:14:00.85" />
                    <SPLIT distance="900" swimtime="00:14:51.65" />
                    <SPLIT distance="950" swimtime="00:15:42.53" />
                    <SPLIT distance="1000" swimtime="00:16:33.39" />
                    <SPLIT distance="1050" swimtime="00:17:24.46" />
                    <SPLIT distance="1100" swimtime="00:18:14.97" />
                    <SPLIT distance="1150" swimtime="00:19:06.25" />
                    <SPLIT distance="1200" swimtime="00:19:56.42" />
                    <SPLIT distance="1250" swimtime="00:20:47.50" />
                    <SPLIT distance="1300" swimtime="00:21:37.57" />
                    <SPLIT distance="1350" swimtime="00:22:28.37" />
                    <SPLIT distance="1400" swimtime="00:23:18.90" />
                    <SPLIT distance="1450" swimtime="00:24:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="568" reactiontime="+94" swimtime="00:00:40.23" resultid="8837" heatid="14202" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="8341" points="347" reactiontime="+73" swimtime="00:03:58.19" resultid="8838" heatid="14259" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:47.62" />
                    <SPLIT distance="150" swimtime="00:02:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="505" reactiontime="+102" swimtime="00:00:38.37" resultid="8839" heatid="14293" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="8486" points="378" reactiontime="+187" swimtime="00:01:40.03" resultid="8840" heatid="14311" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="445" reactiontime="+76" swimtime="00:01:33.79" resultid="8841" heatid="14355" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="442" reactiontime="+97" swimtime="00:03:26.93" resultid="8842" heatid="14368" lane="7" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                    <SPLIT distance="100" swimtime="00:01:38.82" />
                    <SPLIT distance="150" swimtime="00:02:33.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="8826">
              <RESULTS>
                <RESULT eventid="1075" points="216" reactiontime="+96" swimtime="00:00:52.11" resultid="8827" heatid="14144" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1105" points="246" reactiontime="+113" swimtime="00:05:02.92" resultid="8828" heatid="14167" lane="2" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.17" />
                    <SPLIT distance="100" swimtime="00:02:25.24" />
                    <SPLIT distance="150" swimtime="00:03:47.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="218" reactiontime="+83" swimtime="00:01:02.95" resultid="8829" heatid="14199" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="8341" points="178" reactiontime="+109" swimtime="00:06:04.31" resultid="8830" heatid="14258" lane="2" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.22" />
                    <SPLIT distance="100" swimtime="00:02:50.84" />
                    <SPLIT distance="150" swimtime="00:04:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="260" reactiontime="+109" swimtime="00:10:45.71" resultid="8831" heatid="14344" lane="8" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.07" />
                    <SPLIT distance="100" swimtime="00:02:50.68" />
                    <SPLIT distance="150" swimtime="00:04:17.35" />
                    <SPLIT distance="200" swimtime="00:05:37.89" />
                    <SPLIT distance="250" swimtime="00:07:02.19" />
                    <SPLIT distance="300" swimtime="00:08:20.30" />
                    <SPLIT distance="350" swimtime="00:09:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="143" reactiontime="+102" swimtime="00:02:42.41" resultid="8832" heatid="14353" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="333" reactiontime="+83" swimtime="00:04:44.67" resultid="8833" heatid="14367" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.76" />
                    <SPLIT distance="100" swimtime="00:02:19.78" />
                    <SPLIT distance="150" swimtime="00:03:32.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="8843">
              <RESULTS>
                <RESULT eventid="1075" points="605" reactiontime="+66" swimtime="00:00:30.03" resultid="8844" heatid="14150" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1105" points="441" reactiontime="+87" swimtime="00:03:07.04" resultid="8845" heatid="14168" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:28.93" />
                    <SPLIT distance="150" swimtime="00:02:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="524" reactiontime="+74" swimtime="00:01:10.00" resultid="8846" heatid="14227" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="8341" points="322" reactiontime="+86" swimtime="00:03:22.70" resultid="8847" heatid="14259" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                    <SPLIT distance="150" swimtime="00:02:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="441" reactiontime="+86" swimtime="00:00:35.96" resultid="8848" heatid="14294" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="8582" points="388" reactiontime="+94" swimtime="00:07:02.71" resultid="8849" heatid="14343" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:32.46" />
                    <SPLIT distance="150" swimtime="00:02:31.60" />
                    <SPLIT distance="200" swimtime="00:03:33.47" />
                    <SPLIT distance="250" swimtime="00:04:31.64" />
                    <SPLIT distance="300" swimtime="00:05:31.30" />
                    <SPLIT distance="350" swimtime="00:06:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="371" reactiontime="+82" swimtime="00:01:26.66" resultid="8850" heatid="14355" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="388" reactiontime="+82" swimtime="00:00:42.15" resultid="8851" heatid="14382" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="8817">
              <RESULTS>
                <RESULT eventid="1075" points="195" reactiontime="+98" swimtime="00:00:49.93" resultid="8818" heatid="14142" lane="4" />
                <RESULT eventid="1105" points="257" reactiontime="+116" swimtime="00:04:39.26" resultid="8819" heatid="14167" lane="7" entrytime="00:04:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.05" />
                    <SPLIT distance="100" swimtime="00:02:13.71" />
                    <SPLIT distance="150" swimtime="00:03:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="232" reactiontime="+108" swimtime="00:05:01.49" resultid="8820" heatid="14212" lane="1" entrytime="00:04:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.83" />
                    <SPLIT distance="100" swimtime="00:02:24.75" />
                    <SPLIT distance="150" swimtime="00:03:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="212" reactiontime="+122" swimtime="00:02:11.46" resultid="8821" heatid="14245" lane="2" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="206" reactiontime="+110" swimtime="00:02:19.58" resultid="8822" heatid="14276" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="116" reactiontime="+111" swimtime="00:01:06.33" resultid="8823" heatid="14290" lane="3" />
                <RESULT eventid="8662" points="231" reactiontime="+110" swimtime="00:04:56.11" resultid="8824" heatid="14366" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.92" />
                    <SPLIT distance="100" swimtime="00:02:22.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="206" reactiontime="+95" swimtime="00:01:00.12" resultid="8825" heatid="14379" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-02" firstname="Maria" gender="F" lastname="Lippa" nation="POL" athleteid="8802">
              <RESULTS>
                <RESULT eventid="8196" points="110" reactiontime="+156" swimtime="00:01:27.15" resultid="8803" heatid="14193" lane="8" entrytime="00:01:22.00" />
                <RESULT eventid="8229" points="111" reactiontime="+122" swimtime="00:07:23.64" resultid="8804" heatid="14208" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.97" />
                    <SPLIT distance="100" swimtime="00:03:33.69" />
                    <SPLIT distance="150" swimtime="00:05:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="87" swimtime="00:03:38.33" resultid="8805" heatid="14269" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="112" swimtime="00:03:04.41" resultid="8806" heatid="14303" lane="4" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="137" reactiontime="+139" swimtime="00:06:23.70" resultid="8807" heatid="14362" lane="2" entrytime="00:06:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.15" />
                    <SPLIT distance="100" swimtime="00:03:10.06" />
                    <SPLIT distance="150" swimtime="00:04:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="91" reactiontime="+126" swimtime="00:01:35.74" resultid="8808" heatid="14372" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10857" name="Sikret Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@tlen.pl" internet="www.sikret-plywanie.pl" name="Joanna Zagała" phone="601427257" street="Kościuszki 35" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1950-10-13" firstname="Teresa" gender="F" lastname="Żylińska" nation="POL" athleteid="10883">
              <RESULTS>
                <RESULT eventid="1058" points="233" reactiontime="+124" swimtime="00:00:52.36" resultid="10884" heatid="14135" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="8196" points="262" reactiontime="+73" swimtime="00:01:02.56" resultid="10885" heatid="14193" lane="5" entrytime="00:00:57.00" />
                <RESULT eventid="8261" points="217" reactiontime="+101" swimtime="00:01:58.07" resultid="10886" heatid="14218" lane="6" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="264" reactiontime="+138" swimtime="00:02:16.46" resultid="10887" heatid="14304" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="10876">
              <RESULTS>
                <RESULT eventid="1075" points="441" reactiontime="+111" swimtime="00:00:35.26" resultid="10877" heatid="14146" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="8213" points="384" reactiontime="+91" swimtime="00:00:43.72" resultid="10878" heatid="14201" lane="3" entrytime="00:00:42.50" />
                <RESULT eventid="8277" points="375" reactiontime="+96" swimtime="00:01:22.98" resultid="10879" heatid="14227" lane="9" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="371" reactiontime="+76" swimtime="00:01:40.40" resultid="10880" heatid="14311" lane="8" entrytime="00:01:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="406" reactiontime="+99" swimtime="00:03:04.23" resultid="10881" heatid="14325" lane="1" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:15.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="390" reactiontime="+93" swimtime="00:06:43.64" resultid="10882" heatid="14402" lane="1" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:27.10" />
                    <SPLIT distance="150" swimtime="00:02:16.68" />
                    <SPLIT distance="200" swimtime="00:03:07.95" />
                    <SPLIT distance="250" swimtime="00:04:01.48" />
                    <SPLIT distance="300" swimtime="00:04:56.05" />
                    <SPLIT distance="350" swimtime="00:05:50.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="10858">
              <RESULTS>
                <RESULT eventid="1058" points="496" reactiontime="+87" swimtime="00:00:37.35" resultid="10859" heatid="14136" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1135" points="412" reactiontime="+89" swimtime="00:13:38.71" resultid="10860" heatid="14180" lane="6" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="150" swimtime="00:02:27.70" />
                    <SPLIT distance="200" swimtime="00:03:20.13" />
                    <SPLIT distance="350" swimtime="00:07:41.70" />
                    <SPLIT distance="500" swimtime="00:10:18.18" />
                    <SPLIT distance="550" swimtime="00:12:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="410" reactiontime="+93" swimtime="00:00:48.58" resultid="10861" heatid="14193" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="8261" points="445" reactiontime="+85" swimtime="00:01:23.96" resultid="10862" heatid="14219" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="417" reactiontime="+91" swimtime="00:01:51.97" resultid="10863" heatid="14270" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="410" reactiontime="+86" swimtime="00:03:06.11" resultid="10864" heatid="14318" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                    <SPLIT distance="150" swimtime="00:02:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="412" reactiontime="+81" swimtime="00:03:40.94" resultid="10865" heatid="14363" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="100" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:02:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="431" reactiontime="+89" swimtime="00:00:49.72" resultid="10866" heatid="14373" lane="2" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-04-20" firstname="Wojciech" gender="M" lastname="Kosiak" nation="POL" athleteid="10888">
              <RESULTS>
                <RESULT eventid="1075" points="413" reactiontime="+113" swimtime="00:00:42.01" resultid="10889" heatid="14145" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="8277" points="395" reactiontime="+143" swimtime="00:01:36.92" resultid="10890" heatid="14225" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="290" reactiontime="+111" swimtime="00:00:52.20" resultid="10891" heatid="14291" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="8518" points="349" reactiontime="+126" swimtime="00:03:45.69" resultid="10892" heatid="14324" lane="1" entrytime="00:03:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                    <SPLIT distance="100" swimtime="00:01:51.89" />
                    <SPLIT distance="150" swimtime="00:02:53.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="10867">
              <RESULTS>
                <RESULT eventid="1058" points="379" reactiontime="+84" swimtime="00:00:42.85" resultid="10868" heatid="14136" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1135" points="457" reactiontime="+96" swimtime="00:15:36.84" resultid="10869" heatid="14180" lane="7" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.48" />
                    <SPLIT distance="100" swimtime="00:01:45.91" />
                    <SPLIT distance="150" swimtime="00:02:46.90" />
                    <SPLIT distance="200" swimtime="00:03:47.15" />
                    <SPLIT distance="250" swimtime="00:04:46.80" />
                    <SPLIT distance="300" swimtime="00:05:46.43" />
                    <SPLIT distance="350" swimtime="00:06:46.51" />
                    <SPLIT distance="400" swimtime="00:07:46.19" />
                    <SPLIT distance="450" swimtime="00:08:46.10" />
                    <SPLIT distance="500" swimtime="00:09:45.31" />
                    <SPLIT distance="550" swimtime="00:10:44.47" />
                    <SPLIT distance="600" swimtime="00:11:43.95" />
                    <SPLIT distance="650" swimtime="00:12:44.23" />
                    <SPLIT distance="700" swimtime="00:13:43.93" />
                    <SPLIT distance="750" swimtime="00:14:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="427" reactiontime="+95" swimtime="00:04:08.74" resultid="10870" heatid="14208" lane="4" entrytime="00:04:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.76" />
                    <SPLIT distance="100" swimtime="00:02:01.67" />
                    <SPLIT distance="150" swimtime="00:03:05.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="334" reactiontime="+94" swimtime="00:04:52.81" resultid="10871" heatid="14256" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.82" />
                    <SPLIT distance="100" swimtime="00:02:16.87" />
                    <SPLIT distance="150" swimtime="00:03:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="426" reactiontime="+101" swimtime="00:01:54.12" resultid="10872" heatid="14271" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="357" reactiontime="+106" swimtime="00:08:57.17" resultid="10873" heatid="14340" lane="2" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.61" />
                    <SPLIT distance="100" swimtime="00:02:13.82" />
                    <SPLIT distance="150" swimtime="00:03:31.71" />
                    <SPLIT distance="200" swimtime="00:04:44.89" />
                    <SPLIT distance="250" swimtime="00:05:52.93" />
                    <SPLIT distance="300" swimtime="00:06:59.72" />
                    <SPLIT distance="350" swimtime="00:07:59.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="269" reactiontime="+88" swimtime="00:02:06.01" resultid="10874" heatid="14350" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="423" reactiontime="+84" swimtime="00:00:51.11" resultid="10875" heatid="14374" lane="0" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+83" swimtime="00:02:40.44" resultid="10893" heatid="14175" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10858" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="10876" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="10867" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="10888" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+82" swimtime="00:03:04.05" resultid="10894" heatid="14390" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:34.98" />
                    <SPLIT distance="150" swimtime="00:02:25.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10876" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="10867" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="10888" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="10858" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12066" name="SMT Szczecin">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1987-08-03" firstname="Edyta" gender="F" lastname="Adamiak" nation="POL" athleteid="12096">
              <RESULTS>
                <RESULT eventid="8261" points="213" reactiontime="+95" swimtime="00:01:36.13" resultid="12097" heatid="14218" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="226" reactiontime="+92" swimtime="00:01:46.39" resultid="12098" heatid="14238" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="230" reactiontime="+104" swimtime="00:03:25.33" resultid="12099" heatid="14316" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="273" reactiontime="+86" swimtime="00:00:48.27" resultid="12100" heatid="14372" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-20" firstname="Edyta" gender="F" lastname="BARNIK" nation="POL" athleteid="12109">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="12110" heatid="14136" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="8196" status="DNS" swimtime="00:00:00.00" resultid="12111" heatid="14195" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-09" firstname="Łukasz" gender="M" lastname="Rożek" nation="POL" athleteid="12087">
              <RESULTS>
                <RESULT eventid="1075" points="314" reactiontime="+82" swimtime="00:00:32.55" resultid="12088" heatid="14148" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1150" points="241" reactiontime="+82" swimtime="00:13:21.95" resultid="12089" heatid="14185" lane="9" entrytime="00:13:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:26.92" />
                    <SPLIT distance="150" swimtime="00:02:15.00" />
                    <SPLIT distance="200" swimtime="00:03:05.32" />
                    <SPLIT distance="250" swimtime="00:03:55.95" />
                    <SPLIT distance="300" swimtime="00:04:46.67" />
                    <SPLIT distance="350" swimtime="00:05:38.58" />
                    <SPLIT distance="400" swimtime="00:06:30.06" />
                    <SPLIT distance="450" swimtime="00:07:22.34" />
                    <SPLIT distance="500" swimtime="00:08:14.04" />
                    <SPLIT distance="550" swimtime="00:09:06.81" />
                    <SPLIT distance="600" swimtime="00:09:59.05" />
                    <SPLIT distance="650" swimtime="00:10:50.78" />
                    <SPLIT distance="700" swimtime="00:11:42.37" />
                    <SPLIT distance="750" swimtime="00:12:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="260" reactiontime="+93" swimtime="00:01:16.76" resultid="12090" heatid="14227" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="210" reactiontime="+84" swimtime="00:01:32.41" resultid="12091" heatid="14246" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="195" reactiontime="+95" swimtime="00:00:39.42" resultid="12092" heatid="14292" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="8518" points="236" reactiontime="+89" swimtime="00:02:52.27" resultid="12093" heatid="14325" lane="4" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:21.37" />
                    <SPLIT distance="150" swimtime="00:02:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="226" reactiontime="+83" swimtime="00:00:45.65" resultid="12094" heatid="14381" lane="7" entrytime="00:00:47.00" />
                <RESULT eventid="8742" points="262" reactiontime="+84" swimtime="00:06:15.24" resultid="12095" heatid="14404" lane="4" late="yes" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                    <SPLIT distance="200" swimtime="00:02:59.50" />
                    <SPLIT distance="250" swimtime="00:03:48.94" />
                    <SPLIT distance="300" swimtime="00:04:38.20" />
                    <SPLIT distance="350" swimtime="00:05:28.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="12074">
              <RESULTS>
                <RESULT eventid="1075" points="727" reactiontime="+86" swimtime="00:00:25.57" resultid="12075" heatid="14157" lane="0" entrytime="00:00:26.50" />
                <RESULT eventid="8277" points="753" reactiontime="+88" swimtime="00:00:56.52" resultid="12076" heatid="14233" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="629" reactiontime="+81" swimtime="00:01:06.27" resultid="12077" heatid="14253" lane="7" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="654" reactiontime="+79" swimtime="00:00:28.66" resultid="12078" heatid="14296" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="8630" points="623" reactiontime="+79" swimtime="00:01:04.60" resultid="12079" heatid="14358" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="569" reactiontime="+77" swimtime="00:00:34.83" resultid="12080" heatid="14384" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="12101">
              <RESULTS>
                <RESULT eventid="1075" points="518" reactiontime="+67" swimtime="00:00:29.58" resultid="12102" heatid="14153" lane="9" entrytime="00:00:28.80" />
                <RESULT eventid="8277" points="432" reactiontime="+71" swimtime="00:01:08.84" resultid="12103" heatid="14229" lane="6" entrytime="00:01:07.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="413" reactiontime="+68" swimtime="00:01:20.31" resultid="12104" heatid="14248" lane="8" entrytime="00:01:20.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="441" reactiontime="+78" swimtime="00:01:26.19" resultid="12105" heatid="14279" lane="2" entrytime="00:01:29.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="457" reactiontime="+68" swimtime="00:00:32.61" resultid="12106" heatid="14295" lane="8" entrytime="00:00:32.61" />
                <RESULT eventid="8630" points="406" reactiontime="+70" swimtime="00:01:16.44" resultid="12107" heatid="14355" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="451" reactiontime="+75" swimtime="00:00:38.45" resultid="12108" heatid="14385" lane="9" entrytime="00:00:37.61" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="12081">
              <RESULTS>
                <RESULT eventid="1090" points="607" reactiontime="+77" swimtime="00:02:43.03" resultid="12082" heatid="14165" lane="8" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:02:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="611" reactiontime="+76" swimtime="00:01:14.44" resultid="12083" heatid="14242" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="659" reactiontime="+85" swimtime="00:00:32.08" resultid="12084" heatid="14288" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="8470" points="710" reactiontime="+88" swimtime="00:01:12.15" resultid="12085" heatid="14307" lane="1" entrytime="00:01:13.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="580" reactiontime="+70" swimtime="00:01:14.49" resultid="12086" heatid="14352" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="12067">
              <RESULTS>
                <RESULT eventid="1165" points="574" reactiontime="+110" swimtime="00:22:09.46" resultid="12068" heatid="14187" lane="8" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:02.75" />
                    <SPLIT distance="200" swimtime="00:02:46.25" />
                    <SPLIT distance="250" swimtime="00:03:29.95" />
                    <SPLIT distance="300" swimtime="00:04:13.58" />
                    <SPLIT distance="350" swimtime="00:04:57.45" />
                    <SPLIT distance="400" swimtime="00:05:41.21" />
                    <SPLIT distance="450" swimtime="00:06:24.63" />
                    <SPLIT distance="500" swimtime="00:07:08.97" />
                    <SPLIT distance="550" swimtime="00:07:53.00" />
                    <SPLIT distance="600" swimtime="00:08:37.01" />
                    <SPLIT distance="650" swimtime="00:09:20.97" />
                    <SPLIT distance="700" swimtime="00:10:05.38" />
                    <SPLIT distance="750" swimtime="00:10:50.04" />
                    <SPLIT distance="800" swimtime="00:11:34.71" />
                    <SPLIT distance="850" swimtime="00:12:19.87" />
                    <SPLIT distance="900" swimtime="00:13:04.95" />
                    <SPLIT distance="950" swimtime="00:13:50.02" />
                    <SPLIT distance="1000" swimtime="00:14:35.58" />
                    <SPLIT distance="1050" swimtime="00:15:21.27" />
                    <SPLIT distance="1100" swimtime="00:16:06.49" />
                    <SPLIT distance="1150" swimtime="00:16:52.29" />
                    <SPLIT distance="1200" swimtime="00:17:38.12" />
                    <SPLIT distance="1250" swimtime="00:18:23.89" />
                    <SPLIT distance="1300" swimtime="00:19:09.40" />
                    <SPLIT distance="1350" swimtime="00:19:55.55" />
                    <SPLIT distance="1400" swimtime="00:20:41.06" />
                    <SPLIT distance="1450" swimtime="00:21:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="507" reactiontime="+109" swimtime="00:03:11.48" resultid="12069" heatid="14211" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:31.73" />
                    <SPLIT distance="150" swimtime="00:02:22.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="476" reactiontime="+99" swimtime="00:01:28.68" resultid="12070" heatid="14273" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="12071" heatid="14340" lane="1" />
                <RESULT eventid="8613" points="409" reactiontime="+95" swimtime="00:01:25.88" resultid="12072" heatid="14349" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="540" reactiontime="+89" swimtime="00:05:35.75" resultid="12073" heatid="14393" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.37" />
                    <SPLIT distance="200" swimtime="00:02:45.93" />
                    <SPLIT distance="250" swimtime="00:03:29.86" />
                    <SPLIT distance="300" swimtime="00:04:13.83" />
                    <SPLIT distance="350" swimtime="00:04:56.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="SMT SZCZECIN" number="1">
              <RESULTS>
                <RESULT eventid="8534" status="DNS" swimtime="00:00:00.00" resultid="12115" heatid="14335" lane="4" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12081" number="1" />
                    <RELAYPOSITION athleteid="12109" number="2" />
                    <RELAYPOSITION athleteid="12096" number="3" />
                    <RELAYPOSITION athleteid="12067" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT SZCZECIN" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+84" swimtime="00:01:56.44" resultid="12112" heatid="14177" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:00.91" />
                    <SPLIT distance="150" swimtime="00:01:31.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12101" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="12081" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="12067" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="12074" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+93" swimtime="00:02:25.53" resultid="12113" heatid="14392" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:01:54.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12074" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="12096" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="12067" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="12087" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" nation="POL" region="POM" clubid="10540" name="Sopot Masters">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1958-12-28" firstname="Dariusz" gender="M" lastname="Gorbaczow" nation="POL" athleteid="10541">
              <RESULTS>
                <RESULT eventid="1075" points="767" reactiontime="+86" swimtime="00:00:29.31" resultid="10542" heatid="14150" lane="6" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="8213" points="751" reactiontime="+89" swimtime="00:00:34.96" resultid="10543" heatid="14202" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="710" reactiontime="+87" swimtime="00:01:07.09" resultid="10544" heatid="14230" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="810" reactiontime="+83" swimtime="00:00:31.26" resultid="10545" heatid="14296" lane="8" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="10546" heatid="14327" lane="4" entrytime="00:02:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-28" firstname="Wojciech" gender="M" lastname="Kaczmarzyk" nation="POL" athleteid="10547">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="10548" heatid="14157" lane="5" entrytime="00:00:26.20" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="10549" heatid="14174" lane="6" entrytime="00:02:18.00" entrycourse="SCM" />
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="10550" heatid="14206" lane="0" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="10551" heatid="14252" lane="6" entrytime="00:01:08.00" entrycourse="SCM" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="10552" heatid="14301" lane="4" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="10553" heatid="14314" lane="3" entrytime="00:01:06.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-20" firstname="Piotr" gender="M" lastname="Suwara" nation="POL" athleteid="10554">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="10555" heatid="14150" lane="3" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1150" points="476" reactiontime="+94" swimtime="00:10:57.18" resultid="10556" heatid="14183" lane="9" entrytime="00:11:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                    <SPLIT distance="200" swimtime="00:02:39.13" />
                    <SPLIT distance="250" swimtime="00:03:21.59" />
                    <SPLIT distance="300" swimtime="00:04:04.01" />
                    <SPLIT distance="350" swimtime="00:04:46.48" />
                    <SPLIT distance="400" swimtime="00:05:28.74" />
                    <SPLIT distance="450" swimtime="00:06:11.05" />
                    <SPLIT distance="500" swimtime="00:06:54.07" />
                    <SPLIT distance="550" swimtime="00:07:36.33" />
                    <SPLIT distance="600" swimtime="00:08:18.41" />
                    <SPLIT distance="650" swimtime="00:08:59.65" />
                    <SPLIT distance="700" swimtime="00:09:40.65" />
                    <SPLIT distance="750" swimtime="00:10:20.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="421" reactiontime="+89" swimtime="00:00:34.78" resultid="10557" heatid="14202" lane="3" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="528" reactiontime="+94" swimtime="00:01:03.63" resultid="10558" heatid="14229" lane="4" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="435" reactiontime="+105" swimtime="00:01:14.48" resultid="10559" heatid="14311" lane="4" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="456" reactiontime="+96" swimtime="00:02:24.74" resultid="10560" heatid="14329" lane="1" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="150" swimtime="00:01:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="400" reactiontime="+103" swimtime="00:02:44.85" resultid="10561" heatid="14368" lane="3" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="466" reactiontime="+89" swimtime="00:05:12.45" resultid="10562" heatid="14401" lane="5" entrytime="00:05:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:54.82" />
                    <SPLIT distance="200" swimtime="00:02:35.53" />
                    <SPLIT distance="250" swimtime="00:03:16.13" />
                    <SPLIT distance="300" swimtime="00:03:56.47" />
                    <SPLIT distance="350" swimtime="00:04:35.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="12394" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" street="osiedle Stefana Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1982-07-01" firstname="Maciej" gender="M" lastname="Nowaczyk" nation="POL" athleteid="12416">
              <RESULTS>
                <RESULT eventid="8245" points="363" reactiontime="+107" swimtime="00:03:16.95" resultid="12417" heatid="14213" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                    <SPLIT distance="150" swimtime="00:02:24.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="340" reactiontime="+87" swimtime="00:01:13.63" resultid="12418" heatid="14227" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="381" reactiontime="+86" swimtime="00:01:28.28" resultid="12419" heatid="14279" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="12420" heatid="14311" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="8694" points="410" reactiontime="+78" swimtime="00:00:38.86" resultid="12421" heatid="14382" lane="2" entrytime="00:00:42.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-01" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="12403">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="12404" heatid="14137" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1135" points="458" reactiontime="+103" swimtime="00:12:19.48" resultid="12405" heatid="14179" lane="5" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:26.27" />
                    <SPLIT distance="150" swimtime="00:02:11.72" />
                    <SPLIT distance="200" swimtime="00:02:58.15" />
                    <SPLIT distance="250" swimtime="00:03:44.79" />
                    <SPLIT distance="300" swimtime="00:04:32.02" />
                    <SPLIT distance="350" swimtime="00:05:18.56" />
                    <SPLIT distance="400" swimtime="00:06:05.93" />
                    <SPLIT distance="450" swimtime="00:06:53.15" />
                    <SPLIT distance="500" swimtime="00:07:39.77" />
                    <SPLIT distance="550" swimtime="00:08:26.59" />
                    <SPLIT distance="600" swimtime="00:09:13.50" />
                    <SPLIT distance="650" swimtime="00:10:00.77" />
                    <SPLIT distance="700" swimtime="00:10:47.43" />
                    <SPLIT distance="750" swimtime="00:11:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="461" reactiontime="+103" swimtime="00:01:14.38" resultid="12406" heatid="14221" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="364" reactiontime="+110" swimtime="00:03:20.18" resultid="12407" heatid="14257" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                    <SPLIT distance="150" swimtime="00:02:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="446" reactiontime="+92" swimtime="00:00:36.89" resultid="12408" heatid="14288" lane="9" entrytime="00:00:37.30" />
                <RESULT eventid="8502" points="424" reactiontime="+119" swimtime="00:02:47.56" resultid="12409" heatid="14319" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:02:05.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="383" reactiontime="+95" swimtime="00:01:27.83" resultid="12410" heatid="14351" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" status="DNS" swimtime="00:00:00.00" resultid="12411" heatid="14394" lane="0" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-01" firstname="Sławomir" gender="M" lastname="Parysek" nation="POL" athleteid="12446">
              <RESULTS>
                <RESULT eventid="1075" points="530" reactiontime="+96" swimtime="00:00:29.35" resultid="12447" heatid="14152" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="12448" heatid="14184" lane="8" entrytime="00:12:00.00" />
                <RESULT eventid="8277" points="488" reactiontime="+96" swimtime="00:01:06.11" resultid="12449" heatid="14230" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="435" reactiontime="+95" swimtime="00:02:29.15" resultid="12450" heatid="14327" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="328" reactiontime="+84" swimtime="00:01:22.04" resultid="12451" heatid="14355" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="355" reactiontime="+84" swimtime="00:05:39.60" resultid="12452" heatid="14401" lane="1" entrytime="00:05:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                    <SPLIT distance="200" swimtime="00:02:46.20" />
                    <SPLIT distance="250" swimtime="00:03:31.35" />
                    <SPLIT distance="300" swimtime="00:04:16.14" />
                    <SPLIT distance="350" swimtime="00:05:01.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-07-01" firstname="Krzysztof" gender="M" lastname="Kapałczyński" nation="POL" athleteid="12395">
              <RESULTS>
                <RESULT eventid="1105" points="628" reactiontime="+82" swimtime="00:02:46.22" resultid="12396" heatid="14170" lane="6" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:02:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="620" reactiontime="+80" swimtime="00:03:01.38" resultid="12397" heatid="14216" lane="9" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="150" swimtime="00:02:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="488" reactiontime="+84" swimtime="00:02:56.48" resultid="12398" heatid="14260" lane="6" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="580" reactiontime="+89" swimtime="00:01:23.39" resultid="12399" heatid="14281" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="633" reactiontime="+83" swimtime="00:05:59.12" resultid="12400" heatid="14346" lane="3" entrytime="00:05:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                    <SPLIT distance="200" swimtime="00:02:53.94" />
                    <SPLIT distance="250" swimtime="00:03:45.68" />
                    <SPLIT distance="300" swimtime="00:04:37.07" />
                    <SPLIT distance="350" swimtime="00:05:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="512" reactiontime="+83" swimtime="00:01:17.84" resultid="12401" heatid="14357" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="491" reactiontime="+79" swimtime="00:00:38.97" resultid="12402" heatid="14384" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-07-01" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="12412">
              <RESULTS>
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="12413" heatid="14215" lane="2" entrytime="00:03:05.00" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="12414" heatid="14280" lane="6" entrytime="00:01:23.00" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="12415" heatid="14384" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-07-01" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="12437">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="12438" heatid="14164" lane="3" entrytime="00:03:00.00" />
                <RESULT eventid="1135" points="554" reactiontime="+100" swimtime="00:11:34.28" resultid="12439" heatid="14178" lane="0" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:00.17" />
                    <SPLIT distance="200" swimtime="00:02:43.56" />
                    <SPLIT distance="250" swimtime="00:03:27.35" />
                    <SPLIT distance="300" swimtime="00:04:10.93" />
                    <SPLIT distance="350" swimtime="00:04:54.79" />
                    <SPLIT distance="400" swimtime="00:05:38.90" />
                    <SPLIT distance="450" swimtime="00:06:23.24" />
                    <SPLIT distance="500" swimtime="00:07:07.73" />
                    <SPLIT distance="550" swimtime="00:07:51.90" />
                    <SPLIT distance="600" swimtime="00:08:36.62" />
                    <SPLIT distance="650" swimtime="00:09:22.30" />
                    <SPLIT distance="700" swimtime="00:10:07.23" />
                    <SPLIT distance="750" swimtime="00:10:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="617" reactiontime="+85" swimtime="00:00:35.66" resultid="12440" heatid="14197" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="8261" points="567" reactiontime="+97" swimtime="00:01:09.42" resultid="12441" heatid="14222" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="684" reactiontime="+95" swimtime="00:01:15.52" resultid="12442" heatid="14307" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="572" reactiontime="+117" swimtime="00:02:31.63" resultid="12443" heatid="14321" lane="0" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:52.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="660" reactiontime="+88" swimtime="00:02:42.63" resultid="12444" heatid="14365" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:20.59" />
                    <SPLIT distance="150" swimtime="00:02:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="588" reactiontime="+98" swimtime="00:05:26.41" resultid="12445" heatid="14394" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:01:58.62" />
                    <SPLIT distance="200" swimtime="00:02:40.52" />
                    <SPLIT distance="250" swimtime="00:03:21.90" />
                    <SPLIT distance="300" swimtime="00:04:03.88" />
                    <SPLIT distance="350" swimtime="00:04:45.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-07-01" firstname="Anna" gender="F" lastname="Rostkowska-Kaczmarek" nation="POL" athleteid="12431">
              <RESULTS>
                <RESULT eventid="1058" points="572" reactiontime="+90" swimtime="00:00:32.08" resultid="12432" heatid="14138" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1135" points="403" reactiontime="+97" swimtime="00:12:46.67" resultid="12433" heatid="14179" lane="1" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                    <SPLIT distance="150" swimtime="00:02:15.74" />
                    <SPLIT distance="200" swimtime="00:03:02.72" />
                    <SPLIT distance="250" swimtime="00:04:39.24" />
                    <SPLIT distance="300" swimtime="00:06:17.94" />
                    <SPLIT distance="350" swimtime="00:07:07.06" />
                    <SPLIT distance="400" swimtime="00:07:56.82" />
                    <SPLIT distance="450" swimtime="00:08:45.29" />
                    <SPLIT distance="500" swimtime="00:09:33.57" />
                    <SPLIT distance="550" swimtime="00:10:22.12" />
                    <SPLIT distance="600" swimtime="00:11:11.14" />
                    <SPLIT distance="650" swimtime="00:11:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="466" reactiontime="+92" swimtime="00:01:14.54" resultid="12434" heatid="14220" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="397" reactiontime="+98" swimtime="00:02:54.22" resultid="12435" heatid="14319" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="150" swimtime="00:02:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="412" reactiontime="+97" swimtime="00:06:06.88" resultid="12436" heatid="14395" lane="1" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                    <SPLIT distance="150" swimtime="00:02:14.02" />
                    <SPLIT distance="200" swimtime="00:03:00.63" />
                    <SPLIT distance="250" swimtime="00:03:48.15" />
                    <SPLIT distance="300" swimtime="00:04:34.77" />
                    <SPLIT distance="350" swimtime="00:05:22.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-01" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="12422">
              <RESULTS>
                <RESULT eventid="1075" points="833" reactiontime="+80" swimtime="00:00:27.00" resultid="12423" heatid="14155" lane="5" entrytime="00:00:27.10" />
                <RESULT eventid="1105" points="872" reactiontime="+91" swimtime="00:02:28.98" resultid="12424" heatid="14173" lane="1" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="935" reactiontime="+77" swimtime="00:00:57.70" resultid="12425" heatid="14235" lane="8" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="882" reactiontime="+84" swimtime="00:01:07.91" resultid="12426" heatid="14252" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="862" reactiontime="+86" swimtime="00:02:10.86" resultid="12427" heatid="14332" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="854" reactiontime="+79" swimtime="00:05:24.92" resultid="12428" heatid="14347" lane="5" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                    <SPLIT distance="200" swimtime="00:02:36.18" />
                    <SPLIT distance="250" swimtime="00:03:23.69" />
                    <SPLIT distance="300" swimtime="00:04:12.06" />
                    <SPLIT distance="350" swimtime="00:04:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="12429" heatid="14358" lane="7" entrytime="00:01:08.00" />
                <RESULT eventid="8742" points="781" reactiontime="+76" swimtime="00:04:42.77" resultid="12430" heatid="14399" lane="9" entrytime="00:04:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="150" swimtime="00:01:45.52" />
                    <SPLIT distance="200" swimtime="00:02:22.51" />
                    <SPLIT distance="250" swimtime="00:02:58.54" />
                    <SPLIT distance="300" swimtime="00:03:33.52" />
                    <SPLIT distance="350" swimtime="00:04:08.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+84" swimtime="00:02:18.20" resultid="12455" heatid="14266" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:47.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12395" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="12422" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="12446" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="12416" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+83" swimtime="00:02:06.35" resultid="12453" heatid="14176" lane="1" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:37.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12395" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="12403" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="12431" number="3" reactiontime="+84" />
                    <RELAYPOSITION athleteid="12422" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="8710" status="DNS" swimtime="00:00:00.00" resultid="12454" heatid="14391" lane="7" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12437" number="1" />
                    <RELAYPOSITION athleteid="12412" number="2" />
                    <RELAYPOSITION athleteid="12422" number="3" />
                    <RELAYPOSITION athleteid="12431" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="12043" name="Steef Wrocław">
          <CONTACT email="ste1@wp.pl" name="Skrzypek Stefan" phone="500388374" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="12052">
              <RESULTS>
                <RESULT eventid="8179" points="408" reactiontime="+110" swimtime="00:26:23.59" resultid="12053" heatid="14191" lane="6" entrytime="00:26:37.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:33.05" />
                    <SPLIT distance="150" swimtime="00:02:23.39" />
                    <SPLIT distance="200" swimtime="00:03:14.57" />
                    <SPLIT distance="250" swimtime="00:04:06.93" />
                    <SPLIT distance="300" swimtime="00:04:57.52" />
                    <SPLIT distance="350" swimtime="00:05:50.76" />
                    <SPLIT distance="400" swimtime="00:06:44.33" />
                    <SPLIT distance="450" swimtime="00:07:38.27" />
                    <SPLIT distance="500" swimtime="00:08:32.02" />
                    <SPLIT distance="550" swimtime="00:09:26.23" />
                    <SPLIT distance="600" swimtime="00:10:20.23" />
                    <SPLIT distance="650" swimtime="00:11:14.06" />
                    <SPLIT distance="700" swimtime="00:12:08.71" />
                    <SPLIT distance="750" swimtime="00:13:03.18" />
                    <SPLIT distance="800" swimtime="00:13:57.24" />
                    <SPLIT distance="850" swimtime="00:14:50.62" />
                    <SPLIT distance="900" swimtime="00:15:42.71" />
                    <SPLIT distance="950" swimtime="00:16:36.92" />
                    <SPLIT distance="1000" swimtime="00:17:30.41" />
                    <SPLIT distance="1050" swimtime="00:18:24.71" />
                    <SPLIT distance="1100" swimtime="00:19:19.08" />
                    <SPLIT distance="1150" swimtime="00:20:13.31" />
                    <SPLIT distance="1200" swimtime="00:21:08.55" />
                    <SPLIT distance="1250" swimtime="00:22:02.49" />
                    <SPLIT distance="1300" swimtime="00:22:56.36" />
                    <SPLIT distance="1350" swimtime="00:23:49.81" />
                    <SPLIT distance="1400" swimtime="00:24:42.57" />
                    <SPLIT distance="1450" swimtime="00:25:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="451" reactiontime="+104" swimtime="00:02:57.93" resultid="12054" heatid="14325" lane="7" entrytime="00:03:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:26.51" />
                    <SPLIT distance="150" swimtime="00:02:12.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="12044">
              <RESULTS>
                <RESULT eventid="1090" points="687" reactiontime="+101" swimtime="00:03:03.66" resultid="12045" heatid="14164" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:27.04" />
                    <SPLIT distance="150" swimtime="00:02:19.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="740" reactiontime="+105" swimtime="00:00:39.89" resultid="12046" heatid="14195" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="8293" points="671" reactiontime="+94" swimtime="00:01:25.80" resultid="12047" heatid="14241" lane="1" entrytime="00:01:25.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="790" reactiontime="+94" swimtime="00:01:24.49" resultid="12048" heatid="14306" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="843" reactiontime="+115" swimtime="00:06:31.41" resultid="12049" heatid="14341" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:02:23.14" />
                    <SPLIT distance="150" swimtime="00:03:10.77" />
                    <SPLIT distance="200" swimtime="00:04:06.67" />
                    <SPLIT distance="250" swimtime="00:05:02.38" />
                    <SPLIT distance="300" swimtime="00:05:48.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="723" reactiontime="+93" swimtime="00:03:03.24" resultid="12050" heatid="14365" lane="0" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:02:17.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="601" reactiontime="+97" swimtime="00:05:49.44" resultid="12051" heatid="14394" lane="5" entrytime="00:05:50.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:07.63" />
                    <SPLIT distance="200" swimtime="00:02:53.23" />
                    <SPLIT distance="250" swimtime="00:03:38.42" />
                    <SPLIT distance="300" swimtime="00:04:23.32" />
                    <SPLIT distance="350" swimtime="00:05:08.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9793" name="Swim Tri Rzeszów">
          <CONTACT city="RZESZÓW" email="KLUB@SWIMTRI.PL" name="SWIM TRI RZESZÓW" phone="797446677" street="POPIEŁUSZKI 26 C" zip="35-328" />
          <ATHLETES>
            <ATHLETE birthdate="1963-11-15" firstname="Mariusz" gender="M" lastname="Faff" nation="POL" athleteid="9801">
              <RESULTS>
                <RESULT eventid="1075" points="787" reactiontime="+98" swimtime="00:00:28.24" resultid="9802" heatid="14151" lane="4" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="602" reactiontime="+95" swimtime="00:02:52.22" resultid="9803" heatid="14171" lane="7" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="546" reactiontime="+105" swimtime="00:00:35.89" resultid="9804" heatid="14202" lane="5" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="733" reactiontime="+98" swimtime="00:01:04.34" resultid="9805" heatid="14231" lane="3" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="735" reactiontime="+87" swimtime="00:00:31.60" resultid="9806" heatid="14295" lane="7" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="8518" points="685" reactiontime="+154" swimtime="00:02:28.64" resultid="9807" heatid="14328" lane="0" entrytime="00:02:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:11.27" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-10-31" firstname="Tomasz" gender="M" lastname="Sarna" nation="POL" athleteid="9794">
              <RESULTS>
                <RESULT eventid="1075" points="660" reactiontime="+86" swimtime="00:00:27.28" resultid="9795" heatid="14156" lane="9" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="8179" points="602" reactiontime="+105" swimtime="00:19:40.31" resultid="9796" heatid="14190" lane="2" entrytime="00:20:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:46.31" />
                    <SPLIT distance="200" swimtime="00:02:24.92" />
                    <SPLIT distance="250" swimtime="00:03:04.01" />
                    <SPLIT distance="300" swimtime="00:03:43.09" />
                    <SPLIT distance="350" swimtime="00:04:22.17" />
                    <SPLIT distance="400" swimtime="00:05:02.08" />
                    <SPLIT distance="450" swimtime="00:05:42.41" />
                    <SPLIT distance="500" swimtime="00:06:22.30" />
                    <SPLIT distance="550" swimtime="00:07:02.24" />
                    <SPLIT distance="600" swimtime="00:07:42.38" />
                    <SPLIT distance="650" swimtime="00:08:22.50" />
                    <SPLIT distance="700" swimtime="00:09:02.36" />
                    <SPLIT distance="750" swimtime="00:09:42.68" />
                    <SPLIT distance="800" swimtime="00:10:22.73" />
                    <SPLIT distance="850" swimtime="00:11:03.30" />
                    <SPLIT distance="900" swimtime="00:11:43.75" />
                    <SPLIT distance="950" swimtime="00:12:24.40" />
                    <SPLIT distance="1000" swimtime="00:13:05.12" />
                    <SPLIT distance="1050" swimtime="00:13:45.73" />
                    <SPLIT distance="1100" swimtime="00:14:26.29" />
                    <SPLIT distance="1150" swimtime="00:15:07.06" />
                    <SPLIT distance="1200" swimtime="00:15:47.24" />
                    <SPLIT distance="1250" swimtime="00:16:27.64" />
                    <SPLIT distance="1300" swimtime="00:17:07.16" />
                    <SPLIT distance="1350" swimtime="00:17:47.11" />
                    <SPLIT distance="1400" swimtime="00:18:26.65" />
                    <SPLIT distance="1450" swimtime="00:19:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="630" reactiontime="+83" swimtime="00:01:00.71" resultid="9797" heatid="14233" lane="9" entrytime="00:01:01.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="615" reactiontime="+96" swimtime="00:01:10.34" resultid="9798" heatid="14254" lane="0" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="575" reactiontime="+92" swimtime="00:00:30.21" resultid="9799" heatid="14297" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="8518" points="575" reactiontime="+97" swimtime="00:02:15.85" resultid="9800" heatid="14331" lane="1" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:01:03.56" />
                    <SPLIT distance="150" swimtime="00:01:39.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9808" name="Team Karaś  Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1980-01-20" firstname="Ewa" gender="F" lastname="Łukasiuk" nation="POL" athleteid="9809">
              <RESULTS>
                <RESULT eventid="1058" points="544" reactiontime="+91" swimtime="00:00:32.62" resultid="9810" heatid="14139" lane="7" entrytime="00:00:32.59" />
                <RESULT eventid="8261" points="488" reactiontime="+86" swimtime="00:01:13.40" resultid="9811" heatid="14221" lane="0" entrytime="00:01:15.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="463" reactiontime="+74" swimtime="00:05:52.80" resultid="9812" heatid="14394" lane="2" entrytime="00:05:53.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:02:01.80" />
                    <SPLIT distance="200" swimtime="00:02:46.93" />
                    <SPLIT distance="250" swimtime="00:03:33.12" />
                    <SPLIT distance="300" swimtime="00:04:20.74" />
                    <SPLIT distance="350" swimtime="00:05:08.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="9940" name="Team Karaś Płońsk">
          <ATHLETES>
            <ATHLETE birthdate="1989-06-30" firstname="Alan" gender="M" lastname="Bistron" nation="POL" athleteid="9941">
              <RESULTS>
                <RESULT eventid="8245" status="DNS" swimtime="00:00:00.00" resultid="9942" heatid="14212" lane="9" />
                <RESULT eventid="8341" status="DNS" swimtime="00:00:00.00" resultid="9943" heatid="14258" lane="0" />
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="9944" heatid="14308" lane="3" />
                <RESULT eventid="8582" points="226" reactiontime="+100" swimtime="00:07:22.54" resultid="9945" heatid="14343" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:34.69" />
                    <SPLIT distance="150" swimtime="00:02:41.87" />
                    <SPLIT distance="200" swimtime="00:03:45.31" />
                    <SPLIT distance="250" swimtime="00:04:49.50" />
                    <SPLIT distance="300" swimtime="00:05:53.41" />
                    <SPLIT distance="350" swimtime="00:06:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" status="DNS" swimtime="00:00:00.00" resultid="9946" heatid="14366" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="11827" name="TKKF Koszalin Masters">
          <CONTACT email="rpieslak@wp.pl" name="Pieślak Roman" phone="600227112" />
          <ATHLETES>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="11883">
              <RESULTS>
                <RESULT eventid="1075" points="552" reactiontime="+89" swimtime="00:00:29.09" resultid="11884" heatid="14153" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="8277" points="545" reactiontime="+78" swimtime="00:01:04.78" resultid="11885" heatid="14231" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="445" reactiontime="+87" swimtime="00:01:18.68" resultid="11886" heatid="14250" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="499" reactiontime="+89" swimtime="00:00:33.32" resultid="11887" heatid="14295" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="8694" points="418" reactiontime="+88" swimtime="00:00:40.59" resultid="11888" heatid="14385" lane="0" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-14" firstname="Leszek" gender="M" lastname="Szwed" nation="POL" athleteid="11889">
              <RESULTS>
                <RESULT eventid="1075" points="187" reactiontime="+112" swimtime="00:00:44.38" resultid="11890" heatid="14144" lane="2" entrytime="00:00:43.63" />
                <RESULT eventid="8213" points="223" reactiontime="+102" swimtime="00:00:48.20" resultid="11891" heatid="14200" lane="5" entrytime="00:00:49.30" />
                <RESULT eventid="8277" points="180" reactiontime="+95" swimtime="00:01:39.79" resultid="11892" heatid="14225" lane="7" entrytime="00:01:39.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="182" reactiontime="+172" swimtime="00:01:52.19" resultid="11893" heatid="14310" lane="2" entrytime="00:01:48.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-28" firstname="Roman" gender="M" lastname="Pieślak" nation="POL" athleteid="11876">
              <RESULTS>
                <RESULT eventid="8245" points="503" reactiontime="+79" swimtime="00:02:56.68" resultid="11877" heatid="14215" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:08.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="508" reactiontime="+86" swimtime="00:01:04.42" resultid="11878" heatid="14230" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="533" reactiontime="+88" swimtime="00:01:18.92" resultid="11879" heatid="14280" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="431" reactiontime="+110" swimtime="00:02:27.47" resultid="11880" heatid="14328" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="547" reactiontime="+70" swimtime="00:00:35.29" resultid="11881" heatid="14384" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="8742" status="DNS" swimtime="00:00:00.00" resultid="11882" heatid="14401" lane="6" entrytime="00:05:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-25" firstname="Tomasz" gender="M" lastname="Szymanowski" nation="POL" athleteid="11894">
              <RESULTS>
                <RESULT eventid="1075" points="592" reactiontime="+78" swimtime="00:00:28.29" resultid="11895" heatid="14155" lane="7" entrytime="00:00:27.30" />
                <RESULT eventid="1150" points="430" reactiontime="+84" swimtime="00:11:17.47" resultid="11896" heatid="14183" lane="7" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:34.21" />
                    <SPLIT distance="250" swimtime="00:03:15.57" />
                    <SPLIT distance="300" swimtime="00:03:57.79" />
                    <SPLIT distance="350" swimtime="00:04:40.89" />
                    <SPLIT distance="400" swimtime="00:05:24.75" />
                    <SPLIT distance="450" swimtime="00:06:08.60" />
                    <SPLIT distance="500" swimtime="00:06:52.81" />
                    <SPLIT distance="550" swimtime="00:07:37.32" />
                    <SPLIT distance="600" swimtime="00:08:22.48" />
                    <SPLIT distance="650" swimtime="00:09:07.05" />
                    <SPLIT distance="700" swimtime="00:09:52.22" />
                    <SPLIT distance="750" swimtime="00:10:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="558" reactiontime="+86" swimtime="00:00:32.96" resultid="11897" heatid="14205" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="8277" points="580" reactiontime="+91" swimtime="00:01:02.41" resultid="11898" heatid="14233" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="525" reactiontime="+106" swimtime="00:01:13.17" resultid="11899" heatid="14313" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-29" firstname="Lidia" gender="F" lastname="Mikołajczyk" nation="POL" athleteid="11828">
              <RESULTS>
                <RESULT eventid="1090" points="583" reactiontime="+110" swimtime="00:02:51.13" resultid="11829" heatid="14164" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:19.28" />
                    <SPLIT distance="150" swimtime="00:02:09.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="488" reactiontime="+100" swimtime="00:03:13.95" resultid="11830" heatid="14211" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:02:22.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="570" reactiontime="+109" swimtime="00:01:18.17" resultid="11831" heatid="14242" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="471" reactiontime="+112" swimtime="00:01:28.96" resultid="11832" heatid="14273" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="11833" heatid="14342" lane="8" entrytime="00:06:15.00" />
                <RESULT eventid="8678" points="467" reactiontime="+100" swimtime="00:00:40.40" resultid="11834" heatid="14376" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="11853">
              <RESULTS>
                <RESULT eventid="1165" points="537" reactiontime="+103" swimtime="00:25:11.32" resultid="11854" heatid="14187" lane="9" entrytime="00:25:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                    <SPLIT distance="200" swimtime="00:03:13.28" />
                    <SPLIT distance="250" swimtime="00:04:04.11" />
                    <SPLIT distance="300" swimtime="00:04:54.81" />
                    <SPLIT distance="350" swimtime="00:05:45.39" />
                    <SPLIT distance="400" swimtime="00:06:36.03" />
                    <SPLIT distance="450" swimtime="00:07:26.59" />
                    <SPLIT distance="500" swimtime="00:08:17.59" />
                    <SPLIT distance="550" swimtime="00:09:08.71" />
                    <SPLIT distance="600" swimtime="00:09:59.24" />
                    <SPLIT distance="650" swimtime="00:10:49.80" />
                    <SPLIT distance="700" swimtime="00:11:40.31" />
                    <SPLIT distance="750" swimtime="00:12:31.24" />
                    <SPLIT distance="800" swimtime="00:13:21.80" />
                    <SPLIT distance="850" swimtime="00:14:12.38" />
                    <SPLIT distance="900" swimtime="00:15:03.32" />
                    <SPLIT distance="950" swimtime="00:15:53.51" />
                    <SPLIT distance="1000" swimtime="00:16:44.42" />
                    <SPLIT distance="1050" swimtime="00:17:34.92" />
                    <SPLIT distance="1100" swimtime="00:18:25.33" />
                    <SPLIT distance="1150" swimtime="00:19:16.50" />
                    <SPLIT distance="1200" swimtime="00:20:07.55" />
                    <SPLIT distance="1250" swimtime="00:20:58.98" />
                    <SPLIT distance="1300" swimtime="00:21:50.54" />
                    <SPLIT distance="1350" swimtime="00:22:41.34" />
                    <SPLIT distance="1400" swimtime="00:23:32.18" />
                    <SPLIT distance="1450" swimtime="00:24:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" status="DNS" swimtime="00:00:00.00" resultid="11855" heatid="14194" lane="7" entrytime="00:00:48.30" />
                <RESULT eventid="8293" points="440" reactiontime="+107" swimtime="00:01:38.76" resultid="11856" heatid="14239" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="471" reactiontime="+79" swimtime="00:01:40.36" resultid="11857" heatid="14305" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="573" reactiontime="+104" swimtime="00:07:25.12" resultid="11858" heatid="14340" lane="4" entrytime="00:07:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:48.58" />
                    <SPLIT distance="150" swimtime="00:02:45.17" />
                    <SPLIT distance="200" swimtime="00:03:39.47" />
                    <SPLIT distance="250" swimtime="00:04:42.92" />
                    <SPLIT distance="300" swimtime="00:05:46.85" />
                    <SPLIT distance="350" swimtime="00:06:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="455" reactiontime="+85" swimtime="00:03:33.79" resultid="11859" heatid="14364" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="150" swimtime="00:02:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="421" reactiontime="+106" swimtime="00:06:33.49" resultid="11860" heatid="14395" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="150" swimtime="00:02:21.27" />
                    <SPLIT distance="200" swimtime="00:03:11.72" />
                    <SPLIT distance="250" swimtime="00:04:02.28" />
                    <SPLIT distance="300" swimtime="00:04:53.32" />
                    <SPLIT distance="350" swimtime="00:05:44.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="11861">
              <RESULTS>
                <RESULT eventid="1105" points="475" reactiontime="+90" swimtime="00:02:43.89" resultid="11862" heatid="14171" lane="0" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:09.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="467" reactiontime="+94" swimtime="00:21:24.35" resultid="11863" heatid="14190" lane="1" entrytime="00:21:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                    <SPLIT distance="200" swimtime="00:02:43.60" />
                    <SPLIT distance="250" swimtime="00:03:26.36" />
                    <SPLIT distance="300" swimtime="00:04:08.98" />
                    <SPLIT distance="350" swimtime="00:04:51.70" />
                    <SPLIT distance="400" swimtime="00:05:34.24" />
                    <SPLIT distance="450" swimtime="00:06:16.42" />
                    <SPLIT distance="500" swimtime="00:06:58.73" />
                    <SPLIT distance="550" swimtime="00:07:40.93" />
                    <SPLIT distance="600" swimtime="00:08:23.30" />
                    <SPLIT distance="650" swimtime="00:09:05.93" />
                    <SPLIT distance="700" swimtime="00:09:49.11" />
                    <SPLIT distance="750" swimtime="00:10:32.38" />
                    <SPLIT distance="800" swimtime="00:11:15.92" />
                    <SPLIT distance="850" swimtime="00:11:59.63" />
                    <SPLIT distance="900" swimtime="00:12:43.55" />
                    <SPLIT distance="950" swimtime="00:13:27.16" />
                    <SPLIT distance="1000" swimtime="00:14:11.16" />
                    <SPLIT distance="1050" swimtime="00:14:55.64" />
                    <SPLIT distance="1100" swimtime="00:15:39.16" />
                    <SPLIT distance="1150" swimtime="00:16:23.50" />
                    <SPLIT distance="1200" swimtime="00:17:07.93" />
                    <SPLIT distance="1250" swimtime="00:17:52.01" />
                    <SPLIT distance="1300" swimtime="00:18:36.24" />
                    <SPLIT distance="1350" swimtime="00:19:19.88" />
                    <SPLIT distance="1400" swimtime="00:20:04.02" />
                    <SPLIT distance="1450" swimtime="00:20:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="556" reactiontime="+86" swimtime="00:00:33.01" resultid="11864" heatid="14204" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="8309" points="543" reactiontime="+76" swimtime="00:01:13.31" resultid="11865" heatid="14251" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="509" reactiontime="+128" swimtime="00:01:13.95" resultid="11866" heatid="14313" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="11867" heatid="14346" lane="4" entrytime="00:05:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-06" firstname="Joanna" gender="F" lastname="Stankiewicz-Majkowska" nation="POL" athleteid="11842">
              <RESULTS>
                <RESULT eventid="1090" points="353" reactiontime="+94" swimtime="00:03:32.30" resultid="11843" heatid="14163" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                    <SPLIT distance="100" swimtime="00:01:40.34" />
                    <SPLIT distance="150" swimtime="00:02:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="365" reactiontime="+84" swimtime="00:01:36.87" resultid="11844" heatid="14239" lane="5" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="370" reactiontime="+102" swimtime="00:07:30.43" resultid="11845" heatid="14341" lane="8" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:51.31" />
                    <SPLIT distance="150" swimtime="00:02:49.73" />
                    <SPLIT distance="200" swimtime="00:03:46.05" />
                    <SPLIT distance="250" swimtime="00:04:44.94" />
                    <SPLIT distance="300" swimtime="00:05:44.28" />
                    <SPLIT distance="350" swimtime="00:06:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="362" reactiontime="+81" swimtime="00:00:49.29" resultid="11846" heatid="14374" lane="6" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="11847">
              <RESULTS>
                <RESULT eventid="1058" points="521" reactiontime="+84" swimtime="00:00:33.76" resultid="11848" heatid="14138" lane="8" entrytime="00:00:34.70" />
                <RESULT eventid="8196" points="490" reactiontime="+75" swimtime="00:00:38.74" resultid="11849" heatid="14196" lane="9" entrytime="00:00:39.50" />
                <RESULT eventid="8261" points="465" reactiontime="+95" swimtime="00:01:16.67" resultid="11850" heatid="14220" lane="2" entrytime="00:01:18.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="456" reactiontime="+80" swimtime="00:01:28.24" resultid="11851" heatid="14306" lane="0" entrytime="00:01:27.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="519" reactiontime="+79" swimtime="00:03:05.83" resultid="11852" heatid="14364" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:30.79" />
                    <SPLIT distance="150" swimtime="00:02:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-28" firstname="Michał" gender="M" lastname="Pieślak" nation="POL" athleteid="11868">
              <RESULTS>
                <RESULT eventid="1075" points="588" reactiontime="+86" swimtime="00:00:28.36" resultid="11869" heatid="14154" lane="7" entrytime="00:00:27.80" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="11870" heatid="14183" lane="1" entrytime="00:11:00.00" />
                <RESULT eventid="8277" points="555" reactiontime="+86" swimtime="00:01:03.34" resultid="11871" heatid="14232" lane="8" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="11872" heatid="14280" lane="0" entrytime="00:01:25.00" />
                <RESULT eventid="8518" points="479" reactiontime="+79" swimtime="00:02:24.42" resultid="11873" heatid="14329" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="504" reactiontime="+79" swimtime="00:00:37.04" resultid="11874" heatid="14384" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="11835">
              <RESULTS>
                <RESULT eventid="1058" points="603" reactiontime="+86" swimtime="00:00:32.16" resultid="11836" heatid="14140" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="8261" points="529" reactiontime="+101" swimtime="00:01:13.44" resultid="11837" heatid="14222" lane="0" entrytime="00:01:13.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" status="DNS" swimtime="00:00:00.00" resultid="11838" heatid="14271" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="8502" points="501" reactiontime="+110" swimtime="00:02:42.75" resultid="11839" heatid="14320" lane="1" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:17.88" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="11840" heatid="14375" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="8726" points="481" reactiontime="+88" swimtime="00:05:53.45" resultid="11841" heatid="14394" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:07.63" />
                    <SPLIT distance="200" swimtime="00:02:53.36" />
                    <SPLIT distance="250" swimtime="00:03:38.97" />
                    <SPLIT distance="300" swimtime="00:04:24.40" />
                    <SPLIT distance="350" swimtime="00:05:10.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+80" swimtime="00:02:10.49" resultid="11903" heatid="14267" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:42.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11894" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="11876" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="11883" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="11868" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+90" swimtime="00:01:54.45" resultid="11905" heatid="14338" lane="1" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:00:58.19" />
                    <SPLIT distance="150" swimtime="00:01:26.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11868" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="11861" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="11883" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="11894" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="3">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8357" reactiontime="+82" status="DSQ" swimtime="00:02:32.36" resultid="11902" heatid="14264" lane="8" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:27.32" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11847" number="1" reactiontime="+82" status="DSQ" />
                    <RELAYPOSITION athleteid="11842" number="2" reactiontime="+42" status="DSQ" />
                    <RELAYPOSITION athleteid="11828" number="3" reactiontime="-7" status="DSQ" />
                    <RELAYPOSITION athleteid="11835" number="4" reactiontime="+11" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="8534" reactiontime="+104" swimtime="00:02:14.85" resultid="11904" heatid="14335" lane="1" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:43.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11828" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="11847" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="11853" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="11835" number="4" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+87" swimtime="00:01:59.31" resultid="11900" heatid="14176" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:00.41" />
                    <SPLIT distance="150" swimtime="00:01:30.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11835" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="11868" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="11828" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="11894" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+96" swimtime="00:02:15.33" resultid="11901" heatid="14176" lane="0" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11847" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="11883" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="11842" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="11861" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+72" swimtime="00:02:20.38" resultid="11906" heatid="14391" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11847" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="11828" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="11883" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="11868" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="505815" nation="POL" region="WIE" clubid="10666" name="TM Barracuda Kalisz">
          <CONTACT city="KALISZ" email="GALCZYNSKIWOJ@OP.PL" name="GAŁCZYŃSKI WOJCIECH" phone="790690666" state="WLKP" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1982-04-12" firstname="Karolina" gender="F" lastname="Radomska" nation="POL" athleteid="10689">
              <RESULTS>
                <RESULT eventid="8261" points="352" reactiontime="+90" swimtime="00:01:21.83" resultid="10690" heatid="14219" lane="4" entrytime="00:01:22.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="309" reactiontime="+105" swimtime="00:03:09.43" resultid="10691" heatid="14318" lane="6" entrytime="00:03:13.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:20.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="287" reactiontime="+93" swimtime="00:06:53.57" resultid="10692" heatid="14396" lane="7" entrytime="00:07:31.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:32.04" />
                    <SPLIT distance="150" swimtime="00:02:24.78" />
                    <SPLIT distance="200" swimtime="00:03:18.66" />
                    <SPLIT distance="250" swimtime="00:04:12.01" />
                    <SPLIT distance="300" swimtime="00:05:06.02" />
                    <SPLIT distance="350" swimtime="00:06:00.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-27" firstname="Małgorzata" gender="F" lastname="Rembowska-Świeboda" nation="POL" athleteid="10677">
              <RESULTS>
                <RESULT eventid="1058" points="711" reactiontime="+90" swimtime="00:00:31.93" resultid="10678" heatid="14139" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="8196" points="723" reactiontime="+81" swimtime="00:00:36.99" resultid="10679" heatid="14196" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="8293" points="713" reactiontime="+81" swimtime="00:01:20.20" resultid="10680" heatid="14242" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="623" reactiontime="+115" swimtime="00:00:36.47" resultid="10681" heatid="14288" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="8470" points="769" reactiontime="+76" swimtime="00:01:18.81" resultid="10682" heatid="14306" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-13" firstname="Agata" gender="F" lastname="Gałczyńska" nation="POL" athleteid="10667">
              <RESULTS>
                <RESULT eventid="8196" points="119" reactiontime="+93" swimtime="00:01:00.22" resultid="10668" heatid="14193" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="8404" points="152" reactiontime="+104" swimtime="00:02:12.33" resultid="10669" heatid="14270" lane="1" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="153" reactiontime="+87" swimtime="00:00:58.99" resultid="10670" heatid="14373" lane="0" entrytime="00:01:01.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-12" firstname="Wojciech" gender="M" lastname="Gałczyński" nation="POL" athleteid="10671">
              <RESULTS>
                <RESULT eventid="8213" points="561" reactiontime="+69" swimtime="00:00:32.13" resultid="10672" heatid="14205" lane="8" entrytime="00:00:32.45" />
                <RESULT eventid="8309" points="497" reactiontime="+79" swimtime="00:01:09.43" resultid="10673" heatid="14251" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="10674" heatid="14282" lane="6" entrytime="00:01:17.00" />
                <RESULT eventid="8486" points="543" reactiontime="+120" swimtime="00:01:10.54" resultid="10675" heatid="14313" lane="1" entrytime="00:01:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="577" reactiontime="+67" swimtime="00:00:33.40" resultid="10676" heatid="14388" lane="0" entrytime="00:00:33.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-30" firstname="Magdalena" gender="F" lastname="Kolera" nation="POL" athleteid="10683">
              <RESULTS>
                <RESULT eventid="8196" status="DNS" swimtime="00:00:00.00" resultid="10684" heatid="14195" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="8438" status="DNS" swimtime="00:00:00.00" resultid="10685" heatid="14285" lane="3" />
                <RESULT eventid="8470" status="DNS" swimtime="00:00:00.00" resultid="10686" heatid="14305" lane="2" entrytime="00:01:38.00" />
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="10687" heatid="14363" lane="4" entrytime="00:03:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="8357" status="DNS" swimtime="00:00:00.00" resultid="10693" heatid="14263" lane="5" entrytime="00:02:57.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10683" number="1" />
                    <RELAYPOSITION athleteid="10667" number="2" />
                    <RELAYPOSITION athleteid="10677" number="3" />
                    <RELAYPOSITION athleteid="10689" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="8534" status="DNS" swimtime="00:00:00.00" resultid="10694" heatid="14334" lane="5" entrytime="00:02:51.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10667" number="1" />
                    <RELAYPOSITION athleteid="10689" number="2" />
                    <RELAYPOSITION athleteid="10683" number="3" />
                    <RELAYPOSITION athleteid="10677" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="11797" name="Torpedos Marijampole">
          <CONTACT email="vilmantasenator@gmail.com" name="Vilmantas Krasauskas" phone="+370 687 46068" street="R. Jukneviciaus 78-10" street2="Marijampole" />
          <ATHLETES>
            <ATHLETE birthdate="1948-07-09" firstname="Antanas" gender="M" lastname="Guoga" nation="LTU" athleteid="11818">
              <RESULTS>
                <RESULT eventid="1105" points="410" reactiontime="+107" swimtime="00:03:59.21" resultid="11819" heatid="14167" lane="5" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.57" />
                    <SPLIT distance="100" swimtime="00:02:03.12" />
                    <SPLIT distance="150" swimtime="00:03:08.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8179" points="571" reactiontime="+109" swimtime="00:27:50.10" resultid="11820" heatid="14191" lane="8" entrytime="00:27:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                    <SPLIT distance="100" swimtime="00:01:40.96" />
                    <SPLIT distance="150" swimtime="00:02:35.53" />
                    <SPLIT distance="200" swimtime="00:03:30.87" />
                    <SPLIT distance="250" swimtime="00:04:26.68" />
                    <SPLIT distance="300" swimtime="00:05:21.98" />
                    <SPLIT distance="350" swimtime="00:06:17.43" />
                    <SPLIT distance="400" swimtime="00:07:13.27" />
                    <SPLIT distance="450" swimtime="00:08:09.67" />
                    <SPLIT distance="500" swimtime="00:09:05.76" />
                    <SPLIT distance="550" swimtime="00:10:02.26" />
                    <SPLIT distance="600" swimtime="00:10:59.53" />
                    <SPLIT distance="650" swimtime="00:11:56.43" />
                    <SPLIT distance="700" swimtime="00:12:52.40" />
                    <SPLIT distance="750" swimtime="00:13:48.45" />
                    <SPLIT distance="800" swimtime="00:14:44.21" />
                    <SPLIT distance="850" swimtime="00:15:40.19" />
                    <SPLIT distance="900" swimtime="00:16:37.09" />
                    <SPLIT distance="950" swimtime="00:17:33.95" />
                    <SPLIT distance="1000" swimtime="00:18:30.44" />
                    <SPLIT distance="1050" swimtime="00:19:26.61" />
                    <SPLIT distance="1100" swimtime="00:20:22.90" />
                    <SPLIT distance="1150" swimtime="00:21:19.14" />
                    <SPLIT distance="1200" swimtime="00:22:15.87" />
                    <SPLIT distance="1250" swimtime="00:23:12.05" />
                    <SPLIT distance="1300" swimtime="00:24:08.18" />
                    <SPLIT distance="1350" swimtime="00:25:03.44" />
                    <SPLIT distance="1400" swimtime="00:25:59.04" />
                    <SPLIT distance="1450" swimtime="00:26:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="377" reactiontime="+119" swimtime="00:04:16.26" resultid="11821" heatid="14212" lane="3" entrytime="00:04:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.02" />
                    <SPLIT distance="100" swimtime="00:02:02.16" />
                    <SPLIT distance="150" swimtime="00:03:10.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="303" reactiontime="+111" swimtime="00:04:50.33" resultid="11822" heatid="14259" lane="9" entrytime="00:04:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.10" />
                    <SPLIT distance="100" swimtime="00:02:20.26" />
                    <SPLIT distance="150" swimtime="00:03:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="447" reactiontime="+115" swimtime="00:03:16.96" resultid="11823" heatid="14324" lane="3" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="466" reactiontime="+114" swimtime="00:08:30.93" resultid="11824" heatid="14344" lane="5" entrytime="00:08:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.32" />
                    <SPLIT distance="100" swimtime="00:02:17.88" />
                    <SPLIT distance="150" swimtime="00:03:21.91" />
                    <SPLIT distance="200" swimtime="00:04:27.66" />
                    <SPLIT distance="250" swimtime="00:05:38.30" />
                    <SPLIT distance="300" swimtime="00:06:47.04" />
                    <SPLIT distance="350" swimtime="00:07:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="234" reactiontime="+112" swimtime="00:02:11.13" resultid="11825" heatid="14354" lane="2" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="521" reactiontime="+101" swimtime="00:06:55.88" resultid="11826" heatid="14403" lane="5" entrytime="00:06:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:37.33" />
                    <SPLIT distance="150" swimtime="00:02:30.00" />
                    <SPLIT distance="200" swimtime="00:03:23.50" />
                    <SPLIT distance="250" swimtime="00:04:16.99" />
                    <SPLIT distance="300" swimtime="00:05:10.77" />
                    <SPLIT distance="350" swimtime="00:06:04.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-07-31" firstname="Vilmantas" gender="M" lastname="Krasauskas" nation="LTU" athleteid="11804">
              <RESULTS>
                <RESULT eventid="1075" points="688" reactiontime="+87" swimtime="00:00:28.78" resultid="11805" heatid="14152" lane="3" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="8277" points="751" reactiontime="+88" swimtime="00:01:02.09" resultid="11806" heatid="14231" lane="5" entrytime="00:01:03.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="740" reactiontime="+83" swimtime="00:02:17.65" resultid="11807" heatid="14330" lane="8" entrytime="00:02:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:41.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="675" reactiontime="+86" swimtime="00:04:56.83" resultid="11808" heatid="14400" lane="9" entrytime="00:04:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:48.14" />
                    <SPLIT distance="200" swimtime="00:02:26.31" />
                    <SPLIT distance="250" swimtime="00:03:04.62" />
                    <SPLIT distance="300" swimtime="00:03:42.68" />
                    <SPLIT distance="350" swimtime="00:04:20.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-03-14" firstname="Stasys" gender="M" lastname="Grigas" nation="LTU" athleteid="11809">
              <RESULTS>
                <RESULT eventid="1075" points="230" reactiontime="+138" swimtime="00:00:51.02" resultid="11810" heatid="14143" lane="2" entrytime="00:00:51.00" entrycourse="SCM" />
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="11811" heatid="14186" lane="1" entrytime="00:23:40.00" entrycourse="SCM" />
                <RESULT eventid="8213" points="204" reactiontime="+122" swimtime="00:01:04.36" resultid="11812" heatid="14199" lane="3" entrytime="00:01:01.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="139" reactiontime="+130" swimtime="00:02:17.13" resultid="11813" heatid="14224" lane="4" entrytime="00:01:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="127" reactiontime="+121" swimtime="00:02:52.23" resultid="11814" heatid="14276" lane="8" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="182" reactiontime="+124" swimtime="00:02:27.11" resultid="11815" heatid="14309" lane="1" entrytime="00:02:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="213" reactiontime="+101" swimtime="00:05:30.44" resultid="11816" heatid="14366" lane="4" entrytime="00:05:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.13" />
                    <SPLIT distance="100" swimtime="00:02:45.58" />
                    <SPLIT distance="150" swimtime="00:04:10.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="268" reactiontime="+132" swimtime="00:01:00.74" resultid="11817" heatid="14380" lane="1" entrytime="00:01:03.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-04" firstname="Jurate" gender="F" lastname="Pranckeviciene" nation="LTU" athleteid="11798">
              <RESULTS>
                <RESULT eventid="1058" points="506" reactiontime="+88" swimtime="00:00:34.09" resultid="11799" heatid="14138" lane="3" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="8261" points="435" reactiontime="+89" swimtime="00:01:18.38" resultid="11800" heatid="14220" lane="3" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" status="DNS" swimtime="00:00:00.00" resultid="11801" heatid="14286" lane="3" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="11802" heatid="14341" lane="0" entrytime="00:07:30.00" entrycourse="SCM" />
                <RESULT eventid="8613" status="DNS" swimtime="00:00:00.00" resultid="11803" heatid="14350" lane="3" entrytime="00:01:43.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="10340" name="Toruń Multisport Team">
          <CONTACT email="g.arentewicz@onet.pl" name="Grzegorz Arentewicz" phone="535-763-476" />
          <ATHLETES>
            <ATHLETE birthdate="1981-02-04" firstname="Andrzej" gender="M" lastname="Marchewka" nation="POL" athleteid="10364">
              <RESULTS>
                <RESULT eventid="1075" points="671" reactiontime="+90" swimtime="00:00:26.26" resultid="10365" heatid="14146" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1105" points="582" reactiontime="+79" swimtime="00:02:32.42" resultid="10366" heatid="14171" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="599" reactiontime="+79" swimtime="00:00:30.91" resultid="10367" heatid="14204" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="8309" points="641" reactiontime="+92" swimtime="00:01:05.87" resultid="10368" heatid="14250" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="536" reactiontime="+153" swimtime="00:01:09.47" resultid="10369" heatid="14313" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="462" reactiontime="+80" swimtime="00:02:37.23" resultid="10370" heatid="14366" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:16.32" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="668" reactiontime="+78" swimtime="00:00:33.02" resultid="10371" heatid="14385" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-24" firstname="Anita" gender="F" lastname="Śliwa" nation="POL" athleteid="10416">
              <RESULTS>
                <RESULT eventid="1058" points="400" reactiontime="+99" swimtime="00:00:37.05" resultid="10417" heatid="14138" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1135" points="341" reactiontime="+102" swimtime="00:13:44.01" resultid="10418" heatid="14179" lane="7" entrytime="00:13:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:30.63" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                    <SPLIT distance="200" swimtime="00:03:12.58" />
                    <SPLIT distance="250" swimtime="00:04:04.46" />
                    <SPLIT distance="300" swimtime="00:04:56.19" />
                    <SPLIT distance="350" swimtime="00:05:49.02" />
                    <SPLIT distance="400" swimtime="00:06:41.79" />
                    <SPLIT distance="450" swimtime="00:07:34.83" />
                    <SPLIT distance="500" swimtime="00:08:27.68" />
                    <SPLIT distance="550" swimtime="00:09:20.55" />
                    <SPLIT distance="600" swimtime="00:10:14.10" />
                    <SPLIT distance="650" swimtime="00:11:07.76" />
                    <SPLIT distance="700" swimtime="00:12:01.25" />
                    <SPLIT distance="750" swimtime="00:12:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="358" reactiontime="+96" swimtime="00:00:43.40" resultid="10419" heatid="14195" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="8502" points="332" reactiontime="+144" swimtime="00:03:08.42" resultid="10420" heatid="14319" lane="0" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:27.36" />
                    <SPLIT distance="150" swimtime="00:02:18.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="412" reactiontime="+97" swimtime="00:03:26.57" resultid="10421" heatid="14364" lane="7" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:40.46" />
                    <SPLIT distance="150" swimtime="00:02:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" status="DNS" swimtime="00:00:00.00" resultid="10422" entrytime="00:07:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="10429">
              <RESULTS>
                <RESULT eventid="1075" points="74" reactiontime="+121" swimtime="00:01:19.11" resultid="10430" heatid="14143" lane="8" entrytime="00:01:05.10" />
                <RESULT eventid="8213" points="110" reactiontime="+106" swimtime="00:01:30.54" resultid="10431" heatid="14198" lane="4" entrytime="00:01:40.21" />
                <RESULT eventid="8406" status="DNS" swimtime="00:00:00.00" resultid="10432" heatid="14276" lane="9" entrytime="00:02:30.34" />
                <RESULT eventid="8694" points="60" reactiontime="+118" swimtime="00:01:51.35" resultid="10433" heatid="14379" lane="4" entrytime="00:01:25.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-12" firstname="Artur" gender="M" lastname="Kachniarz" nation="POL" athleteid="10359">
              <RESULTS>
                <RESULT eventid="1105" points="493" reactiontime="+98" swimtime="00:02:41.10" resultid="10360" heatid="14171" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:02:04.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="457" reactiontime="+97" swimtime="00:01:13.70" resultid="10361" heatid="14251" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="503" reactiontime="+79" swimtime="00:00:31.28" resultid="10362" heatid="14298" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="8630" points="416" reactiontime="+88" swimtime="00:01:13.94" resultid="10363" heatid="14357" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="10423">
              <RESULTS>
                <RESULT eventid="1075" points="432" reactiontime="+88" swimtime="00:00:30.42" resultid="10424" heatid="14149" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="8277" points="432" reactiontime="+88" swimtime="00:01:07.99" resultid="10425" heatid="14229" lane="3" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="447" reactiontime="+86" swimtime="00:00:32.53" resultid="10426" heatid="14295" lane="0" entrytime="00:00:32.78" />
                <RESULT eventid="8518" points="366" reactiontime="+98" swimtime="00:02:35.70" resultid="10427" heatid="14326" lane="5" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="368" reactiontime="+84" swimtime="00:01:16.99" resultid="10428" heatid="14356" lane="5" entrytime="00:01:17.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Edward" gender="M" lastname="Zientara" nation="POL" athleteid="12725" />
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="10377">
              <RESULTS>
                <RESULT eventid="1150" points="866" reactiontime="+81" swimtime="00:08:59.81" resultid="10378" heatid="14182" lane="4" entrytime="00:08:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:40.14" />
                    <SPLIT distance="200" swimtime="00:02:14.65" />
                    <SPLIT distance="250" swimtime="00:02:48.09" />
                    <SPLIT distance="300" swimtime="00:03:21.35" />
                    <SPLIT distance="350" swimtime="00:03:55.42" />
                    <SPLIT distance="400" swimtime="00:04:29.36" />
                    <SPLIT distance="450" swimtime="00:05:03.58" />
                    <SPLIT distance="500" swimtime="00:05:37.95" />
                    <SPLIT distance="550" swimtime="00:06:12.54" />
                    <SPLIT distance="600" swimtime="00:06:46.89" />
                    <SPLIT distance="650" swimtime="00:07:20.46" />
                    <SPLIT distance="700" swimtime="00:07:54.25" />
                    <SPLIT distance="750" swimtime="00:08:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="925" reactiontime="+79" swimtime="00:02:22.04" resultid="10379" heatid="14217" lane="4" entrytime="00:02:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                    <SPLIT distance="150" swimtime="00:01:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="827" reactiontime="+86" swimtime="00:01:06.07" resultid="10380" heatid="14284" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="854" reactiontime="+75" swimtime="00:04:44.13" resultid="10381" heatid="14348" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:45.37" />
                    <SPLIT distance="200" swimtime="00:02:23.84" />
                    <SPLIT distance="250" swimtime="00:03:01.95" />
                    <SPLIT distance="300" swimtime="00:03:40.67" />
                    <SPLIT distance="350" swimtime="00:04:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="742" reactiontime="+73" swimtime="00:00:59.55" resultid="10382" heatid="14360" lane="4" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8742" points="966" reactiontime="+71" swimtime="00:04:07.23" resultid="10383" heatid="14398" lane="4" entrytime="00:04:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="100" swimtime="00:00:58.86" />
                    <SPLIT distance="150" swimtime="00:01:29.93" />
                    <SPLIT distance="200" swimtime="00:02:01.87" />
                    <SPLIT distance="250" swimtime="00:02:33.80" />
                    <SPLIT distance="300" swimtime="00:03:05.77" />
                    <SPLIT distance="350" swimtime="00:03:37.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="10398">
              <RESULTS>
                <RESULT eventid="1058" points="680" reactiontime="+82" swimtime="00:00:29.72" resultid="10399" heatid="14141" lane="1" entrytime="00:00:29.34" />
                <RESULT eventid="1090" points="745" reactiontime="+68" swimtime="00:02:37.72" resultid="10400" heatid="14165" lane="7" entrytime="00:02:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:02:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="638" reactiontime="+79" swimtime="00:02:57.42" resultid="10401" heatid="14211" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="685" reactiontime="+77" swimtime="00:01:13.54" resultid="10402" heatid="14243" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="590" reactiontime="+71" swimtime="00:01:22.55" resultid="10403" heatid="14274" lane="9" entrytime="00:01:23.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="673" reactiontime="+87" swimtime="00:05:47.53" resultid="10404" heatid="14342" lane="7" entrytime="00:05:40.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                    <SPLIT distance="150" swimtime="00:02:06.17" />
                    <SPLIT distance="200" swimtime="00:02:51.81" />
                    <SPLIT distance="250" swimtime="00:03:39.34" />
                    <SPLIT distance="300" swimtime="00:04:27.99" />
                    <SPLIT distance="350" swimtime="00:05:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="617" reactiontime="+80" swimtime="00:01:14.90" resultid="10405" heatid="14352" lane="0" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="547" reactiontime="+76" swimtime="00:00:38.32" resultid="10406" heatid="14377" lane="9" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="10447">
              <RESULTS>
                <RESULT eventid="1075" points="181" reactiontime="+125" swimtime="00:00:48.72" resultid="10448" heatid="14143" lane="5" entrytime="00:00:48.20" />
                <RESULT eventid="1105" points="142" reactiontime="+123" swimtime="00:05:09.46" resultid="10449" heatid="14167" lane="6" entrytime="00:04:33.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.09" />
                    <SPLIT distance="100" swimtime="00:02:40.66" />
                    <SPLIT distance="150" swimtime="00:04:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="85" reactiontime="+116" swimtime="00:01:15.71" resultid="10450" heatid="14199" lane="1" entrytime="00:01:22.42" />
                <RESULT eventid="8341" points="96" reactiontime="+136" swimtime="00:06:04.88" resultid="10451" heatid="14258" lane="1" entrytime="00:05:48.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.88" />
                    <SPLIT distance="100" swimtime="00:03:02.68" />
                    <SPLIT distance="150" swimtime="00:04:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="81" reactiontime="+88" swimtime="00:02:46.65" resultid="10452" heatid="14309" lane="8" entrytime="00:02:36.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="193" reactiontime="+151" swimtime="00:10:36.60" resultid="10453" heatid="14344" lane="0" entrytime="00:10:40.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.45" />
                    <SPLIT distance="100" swimtime="00:04:32.32" />
                    <SPLIT distance="150" swimtime="00:06:08.04" />
                    <SPLIT distance="200" swimtime="00:07:47.65" />
                    <SPLIT distance="250" swimtime="00:09:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="74" reactiontime="+130" swimtime="00:02:50.32" resultid="10454" heatid="14353" lane="6" entrytime="00:02:31.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="166" reactiontime="+129" swimtime="00:09:17.76" resultid="10455" heatid="14404" lane="5" entrytime="00:08:58.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.66" />
                    <SPLIT distance="100" swimtime="00:02:17.66" />
                    <SPLIT distance="150" swimtime="00:03:34.04" />
                    <SPLIT distance="200" swimtime="00:04:48.52" />
                    <SPLIT distance="250" swimtime="00:06:01.56" />
                    <SPLIT distance="300" swimtime="00:07:12.29" />
                    <SPLIT distance="350" swimtime="00:08:16.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-14" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="10434">
              <RESULTS>
                <RESULT eventid="1075" points="379" reactiontime="+103" swimtime="00:00:43.24" resultid="10435" heatid="14144" lane="6" entrytime="00:00:42.23" />
                <RESULT eventid="8213" points="252" reactiontime="+79" swimtime="00:00:59.97" resultid="10436" heatid="14199" lane="7" entrytime="00:01:05.11" />
                <RESULT eventid="8277" points="318" reactiontime="+113" swimtime="00:01:44.17" resultid="10437" heatid="14225" lane="1" entrytime="00:01:42.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="218" reactiontime="+81" swimtime="00:02:18.42" resultid="10438" heatid="14309" lane="7" entrytime="00:02:12.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="276" swimtime="00:05:03.23" resultid="10439" heatid="14367" lane="0" entrytime="00:04:58.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.24" />
                    <SPLIT distance="100" swimtime="00:02:30.60" />
                    <SPLIT distance="150" swimtime="00:03:49.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="10407">
              <RESULTS>
                <RESULT eventid="1058" points="249" reactiontime="+133" swimtime="00:00:49.24" resultid="10408" heatid="14135" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1135" points="343" reactiontime="+130" swimtime="00:17:10.30" resultid="10409" heatid="14181" lane="5" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                    <SPLIT distance="100" swimtime="00:03:01.95" />
                    <SPLIT distance="150" swimtime="00:04:06.81" />
                    <SPLIT distance="200" swimtime="00:05:12.81" />
                    <SPLIT distance="250" swimtime="00:06:19.43" />
                    <SPLIT distance="300" swimtime="00:07:26.34" />
                    <SPLIT distance="350" swimtime="00:08:31.87" />
                    <SPLIT distance="400" swimtime="00:09:38.45" />
                    <SPLIT distance="450" swimtime="00:10:44.32" />
                    <SPLIT distance="500" swimtime="00:11:50.14" />
                    <SPLIT distance="550" swimtime="00:12:55.07" />
                    <SPLIT distance="600" swimtime="00:14:00.77" />
                    <SPLIT distance="650" swimtime="00:16:10.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="247" reactiontime="+107" swimtime="00:01:01.30" resultid="10410" heatid="14193" lane="7" entrytime="00:01:01.00" />
                <RESULT eventid="8261" points="242" reactiontime="+140" swimtime="00:01:54.58" resultid="10411" heatid="14218" lane="4" entrytime="00:01:54.00" />
                <RESULT eventid="8470" points="259" reactiontime="+92" swimtime="00:02:11.44" resultid="10412" heatid="14304" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="277" reactiontime="+145" swimtime="00:04:03.68" resultid="10413" heatid="14316" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="293" reactiontime="+93" swimtime="00:04:35.25" resultid="10414" heatid="14362" lane="4" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.21" />
                    <SPLIT distance="100" swimtime="00:03:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="268" reactiontime="+129" swimtime="00:09:02.71" resultid="10415" heatid="14396" lane="1" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.69" />
                    <SPLIT distance="100" swimtime="00:02:02.14" />
                    <SPLIT distance="150" swimtime="00:03:09.68" />
                    <SPLIT distance="200" swimtime="00:04:19.55" />
                    <SPLIT distance="250" swimtime="00:05:31.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="10384">
              <RESULTS>
                <RESULT eventid="1105" points="567" reactiontime="+87" swimtime="00:02:33.79" resultid="10385" heatid="14171" lane="5" entrytime="00:02:38.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="520" reactiontime="+83" swimtime="00:00:32.41" resultid="10386" heatid="14205" lane="1" entrytime="00:00:32.45" />
                <RESULT eventid="8309" points="513" reactiontime="+81" swimtime="00:01:10.93" resultid="10387" heatid="14251" lane="9" entrytime="00:01:12.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="509" reactiontime="+113" swimtime="00:01:10.66" resultid="10388" heatid="14313" lane="3" entrytime="00:01:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="558" reactiontime="+83" swimtime="00:05:31.49" resultid="10389" heatid="14347" lane="8" entrytime="00:05:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                    <SPLIT distance="200" swimtime="00:02:36.48" />
                    <SPLIT distance="250" swimtime="00:03:24.88" />
                    <SPLIT distance="300" swimtime="00:04:13.39" />
                    <SPLIT distance="350" swimtime="00:04:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="539" reactiontime="+77" swimtime="00:02:29.31" resultid="10390" heatid="14370" lane="4" entrytime="00:02:28.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:50.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-11" firstname="Kamil" gender="M" lastname="Kordowski" nation="POL" athleteid="10341">
              <RESULTS>
                <RESULT eventid="1075" points="652" reactiontime="+82" swimtime="00:00:26.45" resultid="10342" heatid="14154" lane="6" entrytime="00:00:27.63" />
                <RESULT eventid="8277" points="572" reactiontime="+77" swimtime="00:01:01.00" resultid="10343" heatid="14232" lane="6" entrytime="00:01:01.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="573" reactiontime="+83" swimtime="00:00:29.80" resultid="10344" heatid="14296" lane="5" entrytime="00:00:30.91" />
                <RESULT eventid="8630" points="396" reactiontime="+91" swimtime="00:01:13.96" resultid="10345" heatid="14356" lane="4" entrytime="00:01:17.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-24" firstname="Karolina" gender="F" lastname="Ścisłowicz" nation="POL" athleteid="10391">
              <RESULTS>
                <RESULT eventid="1090" points="329" reactiontime="+87" swimtime="00:03:27.09" resultid="10392" heatid="14164" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                    <SPLIT distance="100" swimtime="00:01:41.88" />
                    <SPLIT distance="150" swimtime="00:02:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit czasu" eventid="1165" reactiontime="+106" status="DSQ" swimtime="00:25:58.87" resultid="10393" heatid="14188" lane="4" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:33.33" />
                    <SPLIT distance="150" swimtime="00:02:24.72" />
                    <SPLIT distance="200" swimtime="00:03:17.45" />
                    <SPLIT distance="250" swimtime="00:04:09.53" />
                    <SPLIT distance="300" swimtime="00:05:01.78" />
                    <SPLIT distance="350" swimtime="00:05:54.00" />
                    <SPLIT distance="400" swimtime="00:06:47.51" />
                    <SPLIT distance="450" swimtime="00:07:40.25" />
                    <SPLIT distance="500" swimtime="00:08:33.00" />
                    <SPLIT distance="550" swimtime="00:09:27.01" />
                    <SPLIT distance="600" swimtime="00:10:19.25" />
                    <SPLIT distance="650" swimtime="00:11:11.53" />
                    <SPLIT distance="700" swimtime="00:12:04.96" />
                    <SPLIT distance="750" swimtime="00:12:57.48" />
                    <SPLIT distance="800" swimtime="00:13:50.53" />
                    <SPLIT distance="850" swimtime="00:14:43.88" />
                    <SPLIT distance="900" swimtime="00:15:37.01" />
                    <SPLIT distance="950" swimtime="00:16:29.64" />
                    <SPLIT distance="1000" swimtime="00:17:22.33" />
                    <SPLIT distance="1050" swimtime="00:18:15.45" />
                    <SPLIT distance="1100" swimtime="00:19:07.77" />
                    <SPLIT distance="1150" swimtime="00:20:00.80" />
                    <SPLIT distance="1200" swimtime="00:20:53.64" />
                    <SPLIT distance="1250" swimtime="00:21:45.92" />
                    <SPLIT distance="1300" swimtime="00:22:38.72" />
                    <SPLIT distance="1350" swimtime="00:23:29.95" />
                    <SPLIT distance="1400" swimtime="00:24:20.98" />
                    <SPLIT distance="1450" swimtime="00:25:11.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="322" reactiontime="+109" swimtime="00:03:42.72" resultid="10394" heatid="14210" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:46.21" />
                    <SPLIT distance="150" swimtime="00:02:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="326" reactiontime="+92" swimtime="00:01:34.13" resultid="10395" heatid="14239" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="247" reactiontime="+102" swimtime="00:00:44.92" resultid="10396" heatid="14286" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="8502" points="354" reactiontime="+112" swimtime="00:02:57.89" resultid="10397" heatid="14319" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-15" firstname="Artur" gender="M" lastname="Rybicki" nation="POL" athleteid="10372">
              <RESULTS>
                <RESULT eventid="1075" points="530" reactiontime="+77" swimtime="00:00:27.34" resultid="10373" heatid="14155" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="8454" points="393" reactiontime="+88" swimtime="00:00:31.20" resultid="10374" heatid="14295" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="8518" points="416" reactiontime="+75" swimtime="00:02:22.68" resultid="10375" heatid="14329" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:46.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="293" reactiontime="+72" swimtime="00:02:55.51" resultid="10376" heatid="14366" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                    <SPLIT distance="150" swimtime="00:02:12.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="10440">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="10441" heatid="14144" lane="9" entrytime="00:00:46.23" />
                <RESULT eventid="8213" points="254" reactiontime="+53" swimtime="00:00:54.74" resultid="10442" heatid="14200" lane="1" entrytime="00:00:52.32" />
                <RESULT eventid="8245" points="298" reactiontime="+108" swimtime="00:04:37.26" resultid="10443" heatid="14212" lane="6" entrytime="00:04:21.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.95" />
                    <SPLIT distance="100" swimtime="00:02:08.16" />
                    <SPLIT distance="150" swimtime="00:03:24.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="274" reactiontime="+100" swimtime="00:02:06.86" resultid="10444" heatid="14276" lane="2" entrytime="00:02:02.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="10445" heatid="14309" lane="2" entrytime="00:02:11.45" />
                <RESULT eventid="8694" points="316" reactiontime="+94" swimtime="00:00:52.13" resultid="10446" heatid="14380" lane="4" entrytime="00:00:51.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-16" firstname="Maciej" gender="M" lastname="Kujawa" nation="POL" athleteid="10346">
              <RESULTS>
                <RESULT eventid="1075" points="490" reactiontime="+98" swimtime="00:00:34.03" resultid="10347" heatid="14147" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="8309" points="531" reactiontime="+94" swimtime="00:01:27.49" resultid="10348" heatid="14247" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="482" reactiontime="+106" swimtime="00:01:34.16" resultid="10349" heatid="14279" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="509" reactiontime="+95" swimtime="00:00:41.00" resultid="10350" heatid="14383" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="10351">
              <RESULTS>
                <RESULT eventid="1075" points="581" reactiontime="+84" swimtime="00:00:33.05" resultid="10352" heatid="14148" lane="1" entrytime="00:00:32.80" />
                <RESULT eventid="1150" points="547" reactiontime="+91" swimtime="00:12:55.48" resultid="10353" heatid="14185" lane="7" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:01:29.58" />
                    <SPLIT distance="150" swimtime="00:02:18.89" />
                    <SPLIT distance="200" swimtime="00:03:08.00" />
                    <SPLIT distance="250" swimtime="00:03:57.28" />
                    <SPLIT distance="300" swimtime="00:04:47.23" />
                    <SPLIT distance="350" swimtime="00:05:37.68" />
                    <SPLIT distance="400" swimtime="00:06:26.80" />
                    <SPLIT distance="450" swimtime="00:07:15.98" />
                    <SPLIT distance="500" swimtime="00:08:04.85" />
                    <SPLIT distance="550" swimtime="00:08:54.37" />
                    <SPLIT distance="600" swimtime="00:09:43.41" />
                    <SPLIT distance="650" swimtime="00:10:33.22" />
                    <SPLIT distance="700" swimtime="00:11:20.75" />
                    <SPLIT distance="750" swimtime="00:12:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="547" reactiontime="+77" swimtime="00:01:14.68" resultid="10354" heatid="14228" lane="9" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="563" reactiontime="+76" swimtime="00:00:37.01" resultid="10355" heatid="14293" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="8518" points="557" reactiontime="+110" swimtime="00:02:53.42" resultid="10356" heatid="14326" lane="1" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="454" reactiontime="+79" swimtime="00:01:33.15" resultid="10357" heatid="14355" lane="3" entrytime="00:01:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="529" reactiontime="+80" swimtime="00:06:19.62" resultid="10358" heatid="14402" lane="2" entrytime="00:06:14.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:16.97" />
                    <SPLIT distance="200" swimtime="00:03:06.66" />
                    <SPLIT distance="250" swimtime="00:03:56.45" />
                    <SPLIT distance="300" swimtime="00:04:46.36" />
                    <SPLIT distance="350" swimtime="00:05:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+74" swimtime="00:01:58.03" resultid="10459" heatid="14268" lane="8" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:00.75" />
                    <SPLIT distance="150" swimtime="00:01:31.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10364" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="10377" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10359" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="10372" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+72" swimtime="00:02:17.73" resultid="10460" heatid="14266" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="150" swimtime="00:01:45.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10384" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="10346" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="10423" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="10351" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+67" swimtime="00:01:45.55" resultid="10461" heatid="14339" lane="9" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.59" />
                    <SPLIT distance="100" swimtime="00:00:53.70" />
                    <SPLIT distance="150" swimtime="00:01:19.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10377" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="10359" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="10364" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="10372" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="8550" swimtime="00:02:05.82" resultid="10462" heatid="14337" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:06.07" />
                    <SPLIT distance="150" swimtime="00:01:36.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10346" number="1" />
                    <RELAYPOSITION athleteid="10351" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="10423" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="10384" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+82" swimtime="00:04:41.05" resultid="12726" heatid="14265" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.21" />
                    <SPLIT distance="100" swimtime="00:02:50.27" />
                    <SPLIT distance="150" swimtime="00:03:58.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12725" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="10429" number="2" reactiontime="+102" />
                    <RELAYPOSITION athleteid="10447" number="3" reactiontime="+96" />
                    <RELAYPOSITION athleteid="10434" number="4" reactiontime="+96" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="10">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="8550" status="DSQ" swimtime="00:03:58.67" resultid="12727" heatid="14336" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.89" />
                    <SPLIT distance="100" swimtime="00:02:23.57" />
                    <SPLIT distance="150" swimtime="00:03:08.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10429" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="12725" number="2" reactiontime="-8" status="DSQ" />
                    <RELAYPOSITION athleteid="10434" number="3" reactiontime="+58" status="DSQ" />
                    <RELAYPOSITION athleteid="10447" number="4" reactiontime="+102" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+92" swimtime="00:02:52.50" resultid="10458" heatid="14263" lane="4" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:01:30.32" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10416" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="10391" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="10398" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="10407" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+105" swimtime="00:01:56.93" resultid="10456" heatid="14177" lane="0" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:32.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10391" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="10398" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="10372" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="10377" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+128" swimtime="00:02:32.51" resultid="10457" heatid="14175" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:01:58.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10407" number="1" reactiontime="+128" />
                    <RELAYPOSITION athleteid="10416" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="10351" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="10346" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+98" swimtime="00:02:11.67" resultid="10463" heatid="14392" lane="0" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:46.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10416" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="10377" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="10398" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="10364" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="10619" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="10620">
              <RESULTS>
                <RESULT eventid="1105" points="500" reactiontime="+105" swimtime="00:03:43.90" resultid="10621" heatid="14168" lane="7" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                    <SPLIT distance="100" swimtime="00:01:48.13" />
                    <SPLIT distance="150" swimtime="00:02:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="435" reactiontime="+79" swimtime="00:00:45.74" resultid="10622" heatid="14201" lane="9" entrytime="00:00:46.00" />
                <RESULT eventid="8309" points="480" reactiontime="+113" swimtime="00:01:40.12" resultid="10623" heatid="14246" lane="2" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="377" reactiontime="+76" swimtime="00:01:43.90" resultid="10624" heatid="14310" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="380" reactiontime="+108" swimtime="00:00:49.02" resultid="10625" heatid="14381" lane="8" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="10626">
              <RESULTS>
                <RESULT eventid="1150" points="381" reactiontime="+92" swimtime="00:14:34.18" resultid="10627" heatid="14186" lane="5" entrytime="00:15:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                    <SPLIT distance="100" swimtime="00:01:47.17" />
                    <SPLIT distance="150" swimtime="00:02:42.85" />
                    <SPLIT distance="200" swimtime="00:03:39.53" />
                    <SPLIT distance="250" swimtime="00:04:35.03" />
                    <SPLIT distance="300" swimtime="00:05:29.50" />
                    <SPLIT distance="350" swimtime="00:06:25.29" />
                    <SPLIT distance="400" swimtime="00:07:19.79" />
                    <SPLIT distance="450" swimtime="00:08:15.02" />
                    <SPLIT distance="500" swimtime="00:09:10.62" />
                    <SPLIT distance="550" swimtime="00:10:05.80" />
                    <SPLIT distance="600" swimtime="00:11:00.70" />
                    <SPLIT distance="650" swimtime="00:11:54.95" />
                    <SPLIT distance="700" swimtime="00:12:49.33" />
                    <SPLIT distance="750" swimtime="00:13:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="366" reactiontime="+97" swimtime="00:00:46.54" resultid="10628" heatid="14201" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="10629" heatid="14310" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="8662" points="354" reactiontime="+95" swimtime="00:03:42.78" resultid="10630" heatid="14368" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:51.29" />
                    <SPLIT distance="150" swimtime="00:02:48.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="376" reactiontime="+101" swimtime="00:07:05.46" resultid="10631" heatid="14403" lane="2" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="100" swimtime="00:01:44.28" />
                    <SPLIT distance="150" swimtime="00:02:39.32" />
                    <SPLIT distance="200" swimtime="00:03:33.37" />
                    <SPLIT distance="250" swimtime="00:04:26.83" />
                    <SPLIT distance="300" swimtime="00:05:19.90" />
                    <SPLIT distance="350" swimtime="00:06:12.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="10645">
              <RESULTS>
                <RESULT eventid="1058" points="430" reactiontime="+101" swimtime="00:00:42.71" resultid="10646" heatid="14136" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1165" points="587" reactiontime="+105" swimtime="00:28:53.79" resultid="10647" heatid="14188" lane="2" entrytime="00:32:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                    <SPLIT distance="100" swimtime="00:01:48.92" />
                    <SPLIT distance="150" swimtime="00:02:47.19" />
                    <SPLIT distance="200" swimtime="00:03:45.12" />
                    <SPLIT distance="250" swimtime="00:04:42.39" />
                    <SPLIT distance="300" swimtime="00:05:40.15" />
                    <SPLIT distance="350" swimtime="00:06:37.09" />
                    <SPLIT distance="400" swimtime="00:07:35.51" />
                    <SPLIT distance="450" swimtime="00:08:35.01" />
                    <SPLIT distance="500" swimtime="00:09:33.29" />
                    <SPLIT distance="550" swimtime="00:10:31.69" />
                    <SPLIT distance="600" swimtime="00:11:31.38" />
                    <SPLIT distance="650" swimtime="00:12:30.91" />
                    <SPLIT distance="700" swimtime="00:13:30.53" />
                    <SPLIT distance="750" swimtime="00:14:29.22" />
                    <SPLIT distance="800" swimtime="00:15:27.95" />
                    <SPLIT distance="850" swimtime="00:16:25.96" />
                    <SPLIT distance="900" swimtime="00:17:25.90" />
                    <SPLIT distance="950" swimtime="00:18:24.93" />
                    <SPLIT distance="1000" swimtime="00:19:24.17" />
                    <SPLIT distance="1050" swimtime="00:20:22.52" />
                    <SPLIT distance="1100" swimtime="00:21:21.81" />
                    <SPLIT distance="1150" swimtime="00:22:20.99" />
                    <SPLIT distance="1200" swimtime="00:23:19.43" />
                    <SPLIT distance="1250" swimtime="00:24:17.03" />
                    <SPLIT distance="1300" swimtime="00:25:16.84" />
                    <SPLIT distance="1350" swimtime="00:26:14.52" />
                    <SPLIT distance="1400" swimtime="00:27:11.15" />
                    <SPLIT distance="1450" swimtime="00:28:05.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="421" reactiontime="+86" swimtime="00:00:53.40" resultid="10648" heatid="14194" lane="9" entrytime="00:00:52.00" />
                <RESULT eventid="8261" points="419" reactiontime="+96" swimtime="00:01:34.83" resultid="10649" heatid="14219" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="356" reactiontime="+97" swimtime="00:00:51.44" resultid="10650" heatid="14286" lane="9" entrytime="00:00:55.00" />
                <RESULT eventid="8502" points="458" reactiontime="+115" swimtime="00:03:32.71" resultid="10651" heatid="14318" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                    <SPLIT distance="100" swimtime="00:01:45.82" />
                    <SPLIT distance="150" swimtime="00:02:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="453" reactiontime="+82" swimtime="00:04:05.32" resultid="10652" heatid="14363" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="100" swimtime="00:02:01.65" />
                    <SPLIT distance="150" swimtime="00:03:05.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="527" reactiontime="+103" swimtime="00:07:16.20" resultid="10653" heatid="14396" lane="3" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:43.75" />
                    <SPLIT distance="150" swimtime="00:02:40.18" />
                    <SPLIT distance="200" swimtime="00:03:37.12" />
                    <SPLIT distance="250" swimtime="00:04:33.94" />
                    <SPLIT distance="300" swimtime="00:05:30.09" />
                    <SPLIT distance="350" swimtime="00:06:24.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="10632">
              <RESULTS>
                <RESULT eventid="1105" points="550" reactiontime="+97" swimtime="00:03:10.84" resultid="10633" heatid="14169" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                    <SPLIT distance="150" swimtime="00:02:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="544" reactiontime="+111" swimtime="00:12:42.27" resultid="10634" heatid="14185" lane="3" entrytime="00:12:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:15.83" />
                    <SPLIT distance="200" swimtime="00:03:04.29" />
                    <SPLIT distance="250" swimtime="00:03:53.27" />
                    <SPLIT distance="300" swimtime="00:04:42.84" />
                    <SPLIT distance="350" swimtime="00:05:31.77" />
                    <SPLIT distance="400" swimtime="00:06:20.18" />
                    <SPLIT distance="450" swimtime="00:07:08.64" />
                    <SPLIT distance="500" swimtime="00:07:56.93" />
                    <SPLIT distance="550" swimtime="00:08:45.53" />
                    <SPLIT distance="600" swimtime="00:09:33.44" />
                    <SPLIT distance="650" swimtime="00:10:21.30" />
                    <SPLIT distance="700" swimtime="00:11:09.09" />
                    <SPLIT distance="750" swimtime="00:11:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="427" reactiontime="+92" swimtime="00:00:42.19" resultid="10635" heatid="14201" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="8309" points="589" reactiontime="+97" swimtime="00:01:24.53" resultid="10636" heatid="14247" lane="6" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="541" reactiontime="+107" swimtime="00:01:28.60" resultid="10637" heatid="14311" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="609" reactiontime="+109" swimtime="00:06:40.51" resultid="10638" heatid="14345" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.42" />
                    <SPLIT distance="100" swimtime="00:01:47.11" />
                    <SPLIT distance="150" swimtime="00:02:36.41" />
                    <SPLIT distance="200" swimtime="00:03:25.46" />
                    <SPLIT distance="250" swimtime="00:04:19.69" />
                    <SPLIT distance="300" swimtime="00:05:14.11" />
                    <SPLIT distance="350" swimtime="00:05:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="616" reactiontime="+89" swimtime="00:03:06.34" resultid="10639" heatid="14368" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                    <SPLIT distance="150" swimtime="00:02:19.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Joanna" gender="F" lastname="Bartosiewicz" nation="POL" athleteid="10654">
              <RESULTS>
                <RESULT eventid="8404" points="648" reactiontime="+93" swimtime="00:01:32.70" resultid="10655" heatid="14272" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="760" reactiontime="+116" swimtime="00:06:04.08" resultid="10656" heatid="14341" lane="2" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:02:12.14" />
                    <SPLIT distance="200" swimtime="00:03:01.10" />
                    <SPLIT distance="250" swimtime="00:03:50.30" />
                    <SPLIT distance="300" swimtime="00:04:41.43" />
                    <SPLIT distance="350" swimtime="00:05:23.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="687" reactiontime="+93" swimtime="00:01:20.17" resultid="10657" heatid="14351" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="680" reactiontime="+96" swimtime="00:00:41.48" resultid="10658" heatid="14374" lane="2" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="10640">
              <RESULTS>
                <RESULT eventid="1150" points="449" reactiontime="+93" swimtime="00:11:41.88" resultid="10641" heatid="14184" lane="5" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:18.88" />
                    <SPLIT distance="150" swimtime="00:02:02.05" />
                    <SPLIT distance="200" swimtime="00:02:46.02" />
                    <SPLIT distance="250" swimtime="00:03:29.73" />
                    <SPLIT distance="300" swimtime="00:04:13.66" />
                    <SPLIT distance="350" swimtime="00:04:57.58" />
                    <SPLIT distance="400" swimtime="00:05:41.70" />
                    <SPLIT distance="450" swimtime="00:06:26.41" />
                    <SPLIT distance="500" swimtime="00:07:11.47" />
                    <SPLIT distance="550" swimtime="00:07:56.45" />
                    <SPLIT distance="600" swimtime="00:08:41.56" />
                    <SPLIT distance="650" swimtime="00:09:26.77" />
                    <SPLIT distance="700" swimtime="00:10:12.59" />
                    <SPLIT distance="750" swimtime="00:10:58.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="500" reactiontime="+82" swimtime="00:03:14.94" resultid="10642" heatid="14214" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:24.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="574" reactiontime="+84" swimtime="00:01:23.66" resultid="10643" heatid="14280" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="604" reactiontime="+78" swimtime="00:00:36.38" resultid="10644" heatid="14385" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+87" swimtime="00:02:42.61" resultid="10659" heatid="14390" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10626" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="10640" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="10654" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="10645" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="WA" clubid="8971" name="UKS Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="PERL" phone="601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1990-05-19" firstname="Dawid" gender="M" lastname="Szulich" nation="POL" athleteid="8990">
              <RESULTS>
                <RESULT eventid="8406" points="964" reactiontime="+71" swimtime="00:01:02.79" resultid="8991" heatid="14284" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="987" reactiontime="+63" swimtime="00:00:28.38" resultid="8992" heatid="14389" lane="5" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-23" firstname="Krzysztof" gender="M" lastname="Żbikowski" nation="POL" athleteid="8984">
              <RESULTS>
                <RESULT eventid="1075" points="714" reactiontime="+76" swimtime="00:00:25.66" resultid="8985" heatid="14159" lane="5" entrytime="00:00:25.00" />
                <RESULT eventid="8245" points="761" reactiontime="+88" swimtime="00:02:30.10" resultid="8986" heatid="14217" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="714" reactiontime="+86" swimtime="00:01:02.91" resultid="8987" heatid="14254" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="818" reactiontime="+77" swimtime="00:01:06.00" resultid="8988" heatid="14284" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="821" reactiontime="+76" swimtime="00:00:30.18" resultid="8989" heatid="14389" lane="1" entrytime="00:00:29.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" athleteid="8972">
              <RESULTS>
                <RESULT eventid="1075" points="920" reactiontime="+70" swimtime="00:00:23.58" resultid="8973" heatid="14161" lane="8" entrytime="00:00:23.78" />
                <RESULT eventid="8277" points="832" reactiontime="+78" swimtime="00:00:53.85" resultid="8974" heatid="14237" lane="1" entrytime="00:00:54.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="822" reactiontime="+74" swimtime="00:01:05.89" resultid="8975" heatid="14284" lane="8" entrytime="00:01:06.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="813" reactiontime="+70" swimtime="00:00:26.52" resultid="8976" heatid="14301" lane="6" entrytime="00:00:26.29" />
                <RESULT eventid="8694" points="927" reactiontime="+70" swimtime="00:00:28.98" resultid="8977" heatid="14389" lane="7" entrytime="00:00:29.41" />
                <RESULT eventid="8742" status="DNS" swimtime="00:00:00.00" resultid="8978" heatid="14400" lane="8" entrytime="00:04:56.96" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-31" firstname="Joanna" gender="F" lastname="Żbikowska" nation="POL" athleteid="8979">
              <RESULTS>
                <RESULT eventid="1058" points="609" reactiontime="+80" swimtime="00:00:30.69" resultid="8980" heatid="14140" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="8293" points="582" reactiontime="+79" swimtime="00:01:15.66" resultid="8981" heatid="14242" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="639" reactiontime="+77" swimtime="00:01:22.09" resultid="8982" heatid="14273" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="709" reactiontime="+73" swimtime="00:00:36.82" resultid="8983" heatid="14377" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="10978" name="UKS Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="11001">
              <RESULTS>
                <RESULT eventid="1058" points="538" reactiontime="+94" swimtime="00:00:33.41" resultid="11002" heatid="14138" lane="4" entrytime="00:00:33.40" />
                <RESULT eventid="1090" points="541" reactiontime="+90" swimtime="00:03:00.13" resultid="11003" heatid="14164" lane="7" entrytime="00:03:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:25.94" />
                    <SPLIT distance="150" swimtime="00:02:18.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="549" reactiontime="+91" swimtime="00:03:22.82" resultid="11004" heatid="14210" lane="6" entrytime="00:03:22.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="528" reactiontime="+86" swimtime="00:01:24.28" resultid="11005" heatid="14240" lane="6" entrytime="00:01:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="533" reactiontime="+89" swimtime="00:01:33.30" resultid="11006" heatid="14272" lane="6" entrytime="00:01:34.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="505" reactiontime="+110" swimtime="00:06:39.60" resultid="11007" heatid="14341" lane="5" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:33.02" />
                    <SPLIT distance="150" swimtime="00:02:25.40" />
                    <SPLIT distance="200" swimtime="00:03:16.23" />
                    <SPLIT distance="250" swimtime="00:04:12.46" />
                    <SPLIT distance="300" swimtime="00:05:08.99" />
                    <SPLIT distance="350" swimtime="00:05:54.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="371" reactiontime="+91" swimtime="00:01:31.95" resultid="11008" heatid="14351" lane="0" entrytime="00:01:30.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="540" reactiontime="+86" swimtime="00:00:42.16" resultid="11009" heatid="14375" lane="4" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="11010">
              <RESULTS>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1105" reactiontime="+90" status="DSQ" swimtime="00:02:25.38" resultid="11011" heatid="14172" lane="0" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="765" reactiontime="+86" swimtime="00:02:41.41" resultid="11012" heatid="14216" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="744" reactiontime="+78" swimtime="00:01:12.90" resultid="11013" heatid="14282" lane="4" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="733" reactiontime="+91" swimtime="00:05:20.61" resultid="11014" heatid="14347" lane="0" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:54.27" />
                    <SPLIT distance="200" swimtime="00:02:36.54" />
                    <SPLIT distance="250" swimtime="00:03:19.55" />
                    <SPLIT distance="300" swimtime="00:04:04.43" />
                    <SPLIT distance="350" swimtime="00:04:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="763" reactiontime="+74" swimtime="00:00:33.23" resultid="11015" heatid="14387" lane="1" entrytime="00:00:34.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" athleteid="11016">
              <RESULTS>
                <RESULT eventid="1105" points="510" reactiontime="+86" swimtime="00:02:49.23" resultid="11017" heatid="14170" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                    <SPLIT distance="150" swimtime="00:02:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="418" reactiontime="+86" swimtime="00:02:56.04" resultid="11018" heatid="14260" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="150" swimtime="00:02:09.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="571" reactiontime="+90" swimtime="00:00:31.86" resultid="11019" heatid="14294" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="8630" points="467" reactiontime="+82" swimtime="00:01:15.75" resultid="11020" heatid="14357" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-14" firstname="Katarzyna" gender="F" lastname="Szwagiel" nation="POL" athleteid="11021">
              <RESULTS>
                <RESULT eventid="1090" points="600" reactiontime="+99" swimtime="00:02:53.96" resultid="11033" heatid="14164" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:02:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="562" reactiontime="+97" swimtime="00:11:36.66" resultid="11034" heatid="14178" lane="9" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:02:03.13" />
                    <SPLIT distance="200" swimtime="00:02:47.26" />
                    <SPLIT distance="250" swimtime="00:03:31.97" />
                    <SPLIT distance="300" swimtime="00:04:16.16" />
                    <SPLIT distance="350" swimtime="00:05:00.90" />
                    <SPLIT distance="400" swimtime="00:05:45.75" />
                    <SPLIT distance="450" swimtime="00:06:30.09" />
                    <SPLIT distance="500" swimtime="00:07:14.89" />
                    <SPLIT distance="550" swimtime="00:07:58.71" />
                    <SPLIT distance="600" swimtime="00:08:42.67" />
                    <SPLIT distance="650" swimtime="00:09:26.41" />
                    <SPLIT distance="700" swimtime="00:10:10.26" />
                    <SPLIT distance="750" swimtime="00:10:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="575" reactiontime="+102" swimtime="00:01:21.93" resultid="11035" heatid="14241" lane="0" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="575" reactiontime="+107" swimtime="00:02:35.51" resultid="11036" heatid="14320" lane="5" entrytime="00:02:39.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8566" points="556" reactiontime="+108" swimtime="00:06:26.88" resultid="11037" heatid="14342" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:31.90" />
                    <SPLIT distance="150" swimtime="00:02:22.85" />
                    <SPLIT distance="200" swimtime="00:03:13.66" />
                    <SPLIT distance="250" swimtime="00:04:07.20" />
                    <SPLIT distance="300" swimtime="00:05:00.77" />
                    <SPLIT distance="350" swimtime="00:05:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" status="DNS" swimtime="00:00:00.00" resultid="11038" heatid="14351" lane="9" entrytime="00:01:31.00" />
                <RESULT eventid="8726" points="550" reactiontime="+99" swimtime="00:05:38.00" resultid="11039" heatid="14394" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:01.73" />
                    <SPLIT distance="200" swimtime="00:02:44.72" />
                    <SPLIT distance="250" swimtime="00:03:28.01" />
                    <SPLIT distance="300" swimtime="00:04:11.95" />
                    <SPLIT distance="350" swimtime="00:04:56.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="10992">
              <RESULTS>
                <RESULT eventid="1075" points="515" reactiontime="+80" swimtime="00:00:29.63" resultid="10993" heatid="14151" lane="7" entrytime="00:00:29.80" />
                <RESULT eventid="1150" points="452" reactiontime="+89" swimtime="00:11:06.73" resultid="10994" heatid="14184" lane="4" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:02:37.14" />
                    <SPLIT distance="250" swimtime="00:03:19.04" />
                    <SPLIT distance="300" swimtime="00:04:01.16" />
                    <SPLIT distance="350" swimtime="00:04:43.60" />
                    <SPLIT distance="400" swimtime="00:05:26.12" />
                    <SPLIT distance="450" swimtime="00:06:08.90" />
                    <SPLIT distance="500" swimtime="00:06:51.31" />
                    <SPLIT distance="550" swimtime="00:07:33.69" />
                    <SPLIT distance="600" swimtime="00:08:16.50" />
                    <SPLIT distance="650" swimtime="00:08:59.85" />
                    <SPLIT distance="700" swimtime="00:09:43.39" />
                    <SPLIT distance="750" swimtime="00:10:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="489" reactiontime="+72" swimtime="00:01:06.09" resultid="10995" heatid="14230" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="342" reactiontime="+90" swimtime="00:03:00.23" resultid="10996" heatid="14260" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:26.61" />
                    <SPLIT distance="150" swimtime="00:02:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="451" reactiontime="+83" swimtime="00:02:27.30" resultid="10997" heatid="14328" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:11.38" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="388" reactiontime="+85" swimtime="00:06:11.49" resultid="10998" heatid="14346" lane="1" entrytime="00:06:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:15.21" />
                    <SPLIT distance="200" swimtime="00:03:01.79" />
                    <SPLIT distance="250" swimtime="00:03:56.92" />
                    <SPLIT distance="300" swimtime="00:04:51.39" />
                    <SPLIT distance="350" swimtime="00:05:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="399" reactiontime="+78" swimtime="00:02:57.15" resultid="10999" heatid="14369" lane="7" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:28.88" />
                    <SPLIT distance="150" swimtime="00:02:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="398" reactiontime="+74" swimtime="00:05:27.09" resultid="11000" heatid="14400" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:56.96" />
                    <SPLIT distance="200" swimtime="00:02:39.16" />
                    <SPLIT distance="250" swimtime="00:03:21.87" />
                    <SPLIT distance="300" swimtime="00:04:04.09" />
                    <SPLIT distance="350" swimtime="00:04:46.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="10987">
              <RESULTS>
                <RESULT eventid="1075" points="737" reactiontime="+81" swimtime="00:00:26.30" resultid="10988" heatid="14150" lane="9" entrytime="00:00:30.34" />
                <RESULT eventid="8277" points="715" reactiontime="+85" swimtime="00:00:58.21" resultid="10989" heatid="14231" lane="7" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="636" reactiontime="+87" swimtime="00:00:29.21" resultid="10990" heatid="14293" lane="5" entrytime="00:00:36.28" />
                <RESULT eventid="8518" points="652" reactiontime="+91" swimtime="00:02:10.30" resultid="10991" heatid="14330" lane="2" entrytime="00:02:16.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="150" swimtime="00:01:37.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="10979">
              <RESULTS>
                <RESULT eventid="1058" points="608" reactiontime="+75" swimtime="00:00:32.08" resultid="10980" heatid="14140" lane="8" entrytime="00:00:31.89" />
                <RESULT eventid="8261" points="557" reactiontime="+91" swimtime="00:01:12.20" resultid="10981" heatid="14222" lane="1" entrytime="00:01:11.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="545" reactiontime="+89" swimtime="00:01:23.40" resultid="10982" heatid="14241" lane="2" entrytime="00:01:22.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="485" reactiontime="+97" swimtime="00:00:38.00" resultid="10983" heatid="14288" lane="0" entrytime="00:00:37.11" />
                <RESULT eventid="8502" points="509" reactiontime="+108" swimtime="00:02:41.88" resultid="10984" heatid="14320" lane="2" entrytime="00:02:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:01.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="366" reactiontime="+86" swimtime="00:01:32.37" resultid="10985" heatid="14351" lane="6" entrytime="00:01:27.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="452" reactiontime="+83" swimtime="00:00:44.73" resultid="10986" heatid="14375" lane="3" entrytime="00:00:43.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+98" swimtime="00:02:08.32" resultid="11031" heatid="14267" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:42.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10992" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="11010" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="11016" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="10987" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+91" swimtime="00:01:53.68" resultid="11032" heatid="14338" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="100" swimtime="00:00:56.05" />
                    <SPLIT distance="150" swimtime="00:01:25.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10987" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="11016" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="10992" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="11010" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+88" swimtime="00:01:59.75" resultid="11029" heatid="14176" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:00:54.78" />
                    <SPLIT distance="150" swimtime="00:01:26.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11010" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="10987" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="10979" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="11001" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+75" swimtime="00:02:16.62" resultid="11030" heatid="14391" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="10979" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="11010" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="11016" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="11021" number="4" reactiontime="+79" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="10248" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska" street2="2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="10249">
              <RESULTS>
                <RESULT eventid="1105" points="338" reactiontime="+93" swimtime="00:04:14.94" resultid="10250" heatid="14168" lane="8" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                    <SPLIT distance="100" swimtime="00:02:02.49" />
                    <SPLIT distance="150" swimtime="00:03:16.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="321" reactiontime="+100" swimtime="00:16:44.46" resultid="10251" heatid="14186" lane="6" entrytime="00:16:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:51.63" />
                    <SPLIT distance="150" swimtime="00:02:52.75" />
                    <SPLIT distance="200" swimtime="00:03:56.92" />
                    <SPLIT distance="250" swimtime="00:05:01.48" />
                    <SPLIT distance="300" swimtime="00:06:05.70" />
                    <SPLIT distance="350" swimtime="00:07:09.54" />
                    <SPLIT distance="400" swimtime="00:08:12.86" />
                    <SPLIT distance="450" swimtime="00:09:17.80" />
                    <SPLIT distance="500" swimtime="00:10:22.13" />
                    <SPLIT distance="550" swimtime="00:11:26.16" />
                    <SPLIT distance="600" swimtime="00:12:29.78" />
                    <SPLIT distance="650" swimtime="00:13:34.14" />
                    <SPLIT distance="700" swimtime="00:14:38.36" />
                    <SPLIT distance="750" swimtime="00:15:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="285" reactiontime="+103" swimtime="00:04:41.44" resultid="10252" heatid="14212" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.61" />
                    <SPLIT distance="100" swimtime="00:02:16.47" />
                    <SPLIT distance="150" swimtime="00:03:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="333" reactiontime="+101" swimtime="00:04:41.38" resultid="10253" heatid="14258" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.93" />
                    <SPLIT distance="100" swimtime="00:02:14.03" />
                    <SPLIT distance="150" swimtime="00:03:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="161" reactiontime="+74" swimtime="00:00:59.38" resultid="10254" heatid="14291" lane="7" entrytime="00:00:54.00" />
                <RESULT eventid="8582" points="398" reactiontime="+94" swimtime="00:08:58.21" resultid="10255" heatid="14344" lane="7" entrytime="00:08:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.83" />
                    <SPLIT distance="100" swimtime="00:02:18.34" />
                    <SPLIT distance="150" swimtime="00:03:22.92" />
                    <SPLIT distance="200" swimtime="00:04:27.49" />
                    <SPLIT distance="250" swimtime="00:05:42.97" />
                    <SPLIT distance="300" swimtime="00:06:58.00" />
                    <SPLIT distance="350" swimtime="00:07:55.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="242" reactiontime="+90" swimtime="00:02:09.57" resultid="10256" heatid="14353" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17414" nation="POL" region="OL" clubid="9472" name="UKS Manta Warszawa Włochy">
          <CONTACT name="Barański" phone="510835478" />
          <ATHLETES>
            <ATHLETE birthdate="1993-09-09" firstname="Michał" gender="M" lastname="Bielawski" nation="POL" license="107414700127" athleteid="9473">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1075" points="956" reactiontime="+65" swimtime="00:00:23.18" resultid="9474" heatid="14161" lane="5" entrytime="00:00:23.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski" eventid="8277" points="935" reactiontime="+69" swimtime="00:00:49.68" resultid="9475" heatid="14237" lane="4" entrytime="00:00:49.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.93" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8518" points="1024" reactiontime="+69" swimtime="00:01:51.65" resultid="9476" heatid="14333" lane="4" entrytime="00:01:53.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                    <SPLIT distance="100" swimtime="00:00:53.61" />
                    <SPLIT distance="150" swimtime="00:01:22.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="879" reactiontime="+64" swimtime="00:00:56.29" resultid="9477" heatid="14360" lane="5" entrytime="00:00:59.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01305" nation="POL" region="LOD" clubid="10715" name="UKS Piątka Konstantynów Łódzki">
          <CONTACT name="Kotus Tomasz" />
          <ATHLETES>
            <ATHLETE birthdate="1981-01-14" firstname="Tomasz" gender="M" lastname="Kotus" nation="POL" athleteid="10721">
              <RESULTS>
                <RESULT eventid="1150" points="530" reactiontime="+102" swimtime="00:10:34.21" resultid="10722" heatid="14184" lane="1" entrytime="00:11:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:10.67" />
                    <SPLIT distance="150" swimtime="00:01:48.88" />
                    <SPLIT distance="200" swimtime="00:02:27.88" />
                    <SPLIT distance="250" swimtime="00:03:07.60" />
                    <SPLIT distance="300" swimtime="00:03:47.60" />
                    <SPLIT distance="350" swimtime="00:04:27.69" />
                    <SPLIT distance="400" swimtime="00:05:07.52" />
                    <SPLIT distance="450" swimtime="00:05:48.24" />
                    <SPLIT distance="500" swimtime="00:06:28.70" />
                    <SPLIT distance="550" swimtime="00:07:09.42" />
                    <SPLIT distance="600" swimtime="00:07:50.14" />
                    <SPLIT distance="650" swimtime="00:08:32.20" />
                    <SPLIT distance="700" swimtime="00:09:13.00" />
                    <SPLIT distance="750" swimtime="00:09:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="451" reactiontime="+97" swimtime="00:02:45.08" resultid="10723" heatid="14259" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="511" reactiontime="+84" swimtime="00:05:41.37" resultid="10724" heatid="14346" lane="9" entrytime="00:06:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                    <SPLIT distance="200" swimtime="00:02:45.94" />
                    <SPLIT distance="250" swimtime="00:03:36.55" />
                    <SPLIT distance="300" swimtime="00:04:26.91" />
                    <SPLIT distance="350" swimtime="00:05:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="10725" heatid="14357" lane="1" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-01" firstname="Krzysztof" gender="M" lastname="Staszak" nation="POL" athleteid="10716">
              <RESULTS>
                <RESULT comment="przekroczony limit czasu" eventid="8179" reactiontime="+96" status="DSQ" swimtime="00:20:46.57" resultid="10717" heatid="14190" lane="3" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.40" />
                    <SPLIT distance="100" swimtime="00:01:56.58" />
                    <SPLIT distance="150" swimtime="00:02:37.58" />
                    <SPLIT distance="200" swimtime="00:03:17.70" />
                    <SPLIT distance="250" swimtime="00:03:57.45" />
                    <SPLIT distance="300" swimtime="00:04:38.60" />
                    <SPLIT distance="350" swimtime="00:05:19.79" />
                    <SPLIT distance="400" swimtime="00:06:00.37" />
                    <SPLIT distance="450" swimtime="00:06:41.72" />
                    <SPLIT distance="500" swimtime="00:07:23.10" />
                    <SPLIT distance="550" swimtime="00:08:04.56" />
                    <SPLIT distance="600" swimtime="00:08:46.52" />
                    <SPLIT distance="650" swimtime="00:09:28.24" />
                    <SPLIT distance="700" swimtime="00:10:51.87" />
                    <SPLIT distance="750" swimtime="00:12:17.46" />
                    <SPLIT distance="800" swimtime="00:12:59.88" />
                    <SPLIT distance="850" swimtime="00:13:42.79" />
                    <SPLIT distance="900" swimtime="00:14:25.30" />
                    <SPLIT distance="950" swimtime="00:15:08.51" />
                    <SPLIT distance="1000" swimtime="00:17:16.31" />
                    <SPLIT distance="1050" swimtime="00:17:58.95" />
                    <SPLIT distance="1100" swimtime="00:18:41.20" />
                    <SPLIT distance="1150" swimtime="00:19:23.56" />
                    <SPLIT distance="1350" swimtime="00:20:05.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="540" reactiontime="+98" swimtime="00:01:00.20" resultid="10718" heatid="14231" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="469" reactiontime="+92" swimtime="00:02:17.03" resultid="10719" heatid="14330" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="374" reactiontime="+107" swimtime="00:02:41.86" resultid="10720" heatid="14369" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRPUL" nation="POL" region="LBL" clubid="9641" name="UKS Trójka Puławy">
          <CONTACT city="Puławy" name="Gogacz" street="Krańcowa" zip="24-100" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" license="500308700164" athleteid="9642">
              <RESULTS>
                <RESULT eventid="8179" points="579" reactiontime="+83" swimtime="00:19:55.74" resultid="9643" heatid="14189" lane="9" entrytime="00:19:29.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:51.20" />
                    <SPLIT distance="200" swimtime="00:02:30.65" />
                    <SPLIT distance="250" swimtime="00:03:10.01" />
                    <SPLIT distance="300" swimtime="00:03:49.67" />
                    <SPLIT distance="350" swimtime="00:04:28.97" />
                    <SPLIT distance="400" swimtime="00:05:08.61" />
                    <SPLIT distance="450" swimtime="00:05:48.47" />
                    <SPLIT distance="500" swimtime="00:06:28.69" />
                    <SPLIT distance="550" swimtime="00:07:08.50" />
                    <SPLIT distance="600" swimtime="00:07:48.05" />
                    <SPLIT distance="650" swimtime="00:08:27.04" />
                    <SPLIT distance="700" swimtime="00:09:06.65" />
                    <SPLIT distance="750" swimtime="00:09:46.16" />
                    <SPLIT distance="800" swimtime="00:10:25.78" />
                    <SPLIT distance="850" swimtime="00:11:05.94" />
                    <SPLIT distance="900" swimtime="00:11:46.20" />
                    <SPLIT distance="950" swimtime="00:12:26.52" />
                    <SPLIT distance="1000" swimtime="00:13:07.23" />
                    <SPLIT distance="1050" swimtime="00:13:47.83" />
                    <SPLIT distance="1100" swimtime="00:14:27.82" />
                    <SPLIT distance="1150" swimtime="00:15:08.71" />
                    <SPLIT distance="1200" swimtime="00:15:49.82" />
                    <SPLIT distance="1250" swimtime="00:16:30.33" />
                    <SPLIT distance="1300" swimtime="00:17:11.42" />
                    <SPLIT distance="1350" swimtime="00:17:52.30" />
                    <SPLIT distance="1400" swimtime="00:18:33.40" />
                    <SPLIT distance="1450" swimtime="00:19:14.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="582" reactiontime="+89" swimtime="00:02:30.92" resultid="9644" heatid="14261" lane="5" entrytime="00:02:30.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="9645" heatid="14347" lane="2" entrytime="00:05:38.19" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" nation="POL" region="MAZ" clubid="11907" name="UKS Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="11908">
              <RESULTS>
                <RESULT eventid="1150" points="540" reactiontime="+80" swimtime="00:11:00.12" resultid="11909" heatid="14183" lane="6" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                    <SPLIT distance="200" swimtime="00:02:39.94" />
                    <SPLIT distance="250" swimtime="00:03:22.59" />
                    <SPLIT distance="300" swimtime="00:04:05.00" />
                    <SPLIT distance="350" swimtime="00:04:47.37" />
                    <SPLIT distance="400" swimtime="00:05:29.42" />
                    <SPLIT distance="450" swimtime="00:06:10.82" />
                    <SPLIT distance="500" swimtime="00:06:52.52" />
                    <SPLIT distance="550" swimtime="00:07:34.54" />
                    <SPLIT distance="600" swimtime="00:08:15.96" />
                    <SPLIT distance="650" swimtime="00:08:57.63" />
                    <SPLIT distance="700" swimtime="00:09:39.21" />
                    <SPLIT distance="750" swimtime="00:10:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="600" reactiontime="+81" swimtime="00:03:03.38" resultid="11910" heatid="14215" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:27.86" />
                    <SPLIT distance="150" swimtime="00:02:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="11911" heatid="14250" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="8406" points="619" reactiontime="+86" swimtime="00:01:21.58" resultid="11912" heatid="14280" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="11913" heatid="14347" lane="1" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="KA" clubid="11195" name="UKS Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas" />
          <ATHLETES>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="11201">
              <RESULTS>
                <RESULT eventid="1075" points="710" reactiontime="+100" swimtime="00:00:30.08" resultid="11202" heatid="14151" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="8277" points="632" reactiontime="+97" swimtime="00:01:09.75" resultid="11203" heatid="14229" lane="9" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="570" reactiontime="+106" swimtime="00:03:12.59" resultid="11204" heatid="14260" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="702" reactiontime="+100" swimtime="00:00:32.79" resultid="11205" heatid="14295" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="8630" points="725" reactiontime="+96" swimtime="00:01:15.01" resultid="11206" heatid="14356" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="11207">
              <RESULTS>
                <RESULT eventid="1075" points="695" reactiontime="+91" swimtime="00:00:28.68" resultid="11208" heatid="14152" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1150" points="578" reactiontime="+116" swimtime="00:10:45.39" resultid="11209" heatid="14183" lane="0" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="150" swimtime="00:01:49.02" />
                    <SPLIT distance="200" swimtime="00:02:29.26" />
                    <SPLIT distance="250" swimtime="00:03:10.10" />
                    <SPLIT distance="300" swimtime="00:03:51.04" />
                    <SPLIT distance="350" swimtime="00:04:32.35" />
                    <SPLIT distance="400" swimtime="00:05:13.49" />
                    <SPLIT distance="450" swimtime="00:05:54.67" />
                    <SPLIT distance="500" swimtime="00:06:36.03" />
                    <SPLIT distance="550" swimtime="00:07:17.51" />
                    <SPLIT distance="600" swimtime="00:07:58.92" />
                    <SPLIT distance="650" swimtime="00:08:40.44" />
                    <SPLIT distance="700" swimtime="00:09:22.46" />
                    <SPLIT distance="750" swimtime="00:10:04.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="738" reactiontime="+94" swimtime="00:01:02.44" resultid="11210" heatid="14230" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="503" reactiontime="+92" swimtime="00:02:54.63" resultid="11211" heatid="14260" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:20.79" />
                    <SPLIT distance="150" swimtime="00:02:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="592" reactiontime="+108" swimtime="00:01:15.78" resultid="11212" heatid="14312" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="666" reactiontime="+91" swimtime="00:02:22.59" resultid="11213" heatid="14328" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="605" reactiontime="+97" swimtime="00:02:44.52" resultid="11214" heatid="14369" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:02.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="11196">
              <RESULTS>
                <RESULT eventid="1075" points="591" reactiontime="+92" swimtime="00:00:31.07" resultid="11197" heatid="14148" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="8245" points="768" reactiontime="+94" swimtime="00:02:56.90" resultid="11198" heatid="14215" lane="4" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:24.72" />
                    <SPLIT distance="150" swimtime="00:02:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="638" reactiontime="+81" swimtime="00:01:19.12" resultid="11199" heatid="14281" lane="4" entrytime="00:01:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="643" reactiontime="+79" swimtime="00:00:35.32" resultid="11200" heatid="14386" lane="3" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="11216">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="11217" heatid="14135" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1135" status="DNS" swimtime="00:00:00.00" resultid="11218" heatid="14181" lane="3" entrytime="00:24:00.00" />
                <RESULT eventid="8196" status="DNS" swimtime="00:00:00.00" resultid="11219" heatid="14193" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="8261" status="DNS" swimtime="00:00:00.00" resultid="11220" heatid="14218" lane="1" entrytime="00:02:40.00" />
                <RESULT eventid="8470" status="DNS" swimtime="00:00:00.00" resultid="11221" heatid="14304" lane="8" entrytime="00:02:40.00" />
                <RESULT eventid="8646" status="DNS" swimtime="00:00:00.00" resultid="11222" heatid="14362" lane="3" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="8895" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="8896">
              <RESULTS>
                <RESULT eventid="1075" points="580" reactiontime="+93" swimtime="00:00:28.62" resultid="8897" heatid="14151" lane="3" entrytime="00:00:29.30" />
                <RESULT eventid="8277" points="581" reactiontime="+81" swimtime="00:01:03.39" resultid="8898" heatid="14231" lane="8" entrytime="00:01:04.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="518" reactiontime="+78" swimtime="00:00:32.92" resultid="8899" heatid="14294" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="8518" points="463" reactiontime="+79" swimtime="00:02:28.24" resultid="8900" heatid="14328" lane="9" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="8901" heatid="14356" lane="0" entrytime="00:01:26.00" />
                <RESULT eventid="8742" points="408" reactiontime="+81" swimtime="00:05:31.49" resultid="8902" heatid="14404" lane="0" late="yes" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:55.11" />
                    <SPLIT distance="200" swimtime="00:02:38.52" />
                    <SPLIT distance="250" swimtime="00:03:22.60" />
                    <SPLIT distance="300" swimtime="00:04:07.56" />
                    <SPLIT distance="350" swimtime="00:04:52.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031/05" nation="POL" region="LOD" clubid="9830" name="UTW Masters Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="9925">
              <RESULTS>
                <RESULT eventid="1105" points="674" reactiontime="+88" swimtime="00:02:14.71" resultid="9926" heatid="14166" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                    <SPLIT distance="150" swimtime="00:01:41.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="9927" heatid="14244" lane="5" />
                <RESULT eventid="8518" points="690" reactiontime="+93" swimtime="00:02:00.49" resultid="9928" heatid="14322" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                    <SPLIT distance="150" swimtime="00:01:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="736" reactiontime="+78" swimtime="00:00:58.29" resultid="9929" heatid="14353" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-06" firstname="Robert" gender="M" lastname="Szalbierz" nation="POL" license="503105700056" athleteid="9844">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="9845" heatid="14152" lane="1" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="9846" heatid="14229" lane="2" entrytime="00:01:08.00" entrycourse="SCM" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="9847" heatid="14249" lane="1" entrytime="00:01:18.00" entrycourse="SCM" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="9848" heatid="14294" lane="6" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="9849" heatid="14327" lane="9" entrytime="00:02:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="9880">
              <RESULTS>
                <RESULT eventid="8245" points="367" reactiontime="+116" swimtime="00:03:46.24" resultid="9881" heatid="14213" lane="1" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.89" />
                    <SPLIT distance="100" swimtime="00:01:47.44" />
                    <SPLIT distance="150" swimtime="00:02:48.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="326" reactiontime="+135" swimtime="00:01:38.90" resultid="9882" heatid="14278" lane="1" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="366" reactiontime="+111" swimtime="00:00:42.62" resultid="9883" heatid="14383" lane="0" entrytime="00:00:41.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-25" firstname="Joanna" gender="F" lastname="Kańska-Papiernik" nation="POL" license="503105600" athleteid="9859">
              <RESULTS>
                <RESULT eventid="8196" points="549" reactiontime="+81" swimtime="00:00:37.29" resultid="9860" heatid="14197" lane="0" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="8293" points="602" reactiontime="+75" swimtime="00:01:20.67" resultid="9861" heatid="14242" lane="8" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="616" reactiontime="+88" swimtime="00:01:28.95" resultid="9862" heatid="14273" lane="2" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="597" reactiontime="+73" swimtime="00:01:20.68" resultid="9863" heatid="14306" lane="4" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="9864" heatid="14377" lane="1" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Woźniak" nation="POL" license="503105700039" athleteid="9873">
              <RESULTS>
                <RESULT eventid="8213" points="710" reactiontime="+61" swimtime="00:00:29.22" resultid="9874" heatid="14206" lane="4" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="9875" heatid="14253" lane="1" entrytime="00:01:07.00" entrycourse="SCM" />
                <RESULT eventid="8454" points="685" reactiontime="+77" swimtime="00:00:28.22" resultid="9876" heatid="14290" lane="4" />
                <RESULT eventid="8486" points="690" reactiontime="+70" swimtime="00:01:03.88" resultid="9877" heatid="14315" lane="0" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9878" heatid="14353" lane="1" />
                <RESULT eventid="8662" points="638" reactiontime="+63" swimtime="00:02:21.14" resultid="9879" heatid="14371" lane="7" entrytime="00:02:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-12" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="9919">
              <RESULTS>
                <RESULT eventid="1075" points="605" reactiontime="+92" swimtime="00:00:34.27" resultid="9920" heatid="14147" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="9921" heatid="14200" lane="4" entrytime="00:00:48.00" entrycourse="SCM" />
                <RESULT eventid="8277" points="563" reactiontime="+107" swimtime="00:01:22.14" resultid="9922" heatid="14226" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="476" reactiontime="+78" swimtime="00:00:41.42" resultid="9923" heatid="14293" lane="7" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="8630" points="387" reactiontime="+92" swimtime="00:01:50.82" resultid="9924" heatid="14354" lane="4" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-05-30" firstname="Adrianna" gender="F" lastname="Rzewuska" nation="POL" license="503105600" athleteid="9891">
              <RESULTS>
                <RESULT eventid="8196" points="708" reactiontime="+80" swimtime="00:00:32.85" resultid="9892" heatid="14197" lane="2" entrytime="00:00:32.50" entrycourse="SCM" />
                <RESULT eventid="8470" points="727" reactiontime="+90" swimtime="00:01:11.61" resultid="9893" heatid="14307" lane="2" entrytime="00:01:11.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="570" reactiontime="+74" swimtime="00:02:38.94" resultid="9894" heatid="14365" lane="6" entrytime="00:02:38.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8726" points="397" reactiontime="+72" swimtime="00:05:49.12" resultid="9895" heatid="14394" lane="4" entrytime="00:05:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="150" swimtime="00:02:01.21" />
                    <SPLIT distance="200" swimtime="00:02:46.17" />
                    <SPLIT distance="250" swimtime="00:03:32.33" />
                    <SPLIT distance="300" swimtime="00:04:18.77" />
                    <SPLIT distance="350" swimtime="00:05:04.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="9884">
              <RESULTS>
                <RESULT eventid="1150" points="675" reactiontime="+96" swimtime="00:11:49.35" resultid="9885" heatid="14185" lane="5" entrytime="00:12:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.15" />
                    <SPLIT distance="150" swimtime="00:02:04.03" />
                    <SPLIT distance="200" swimtime="00:02:48.95" />
                    <SPLIT distance="250" swimtime="00:03:34.22" />
                    <SPLIT distance="300" swimtime="00:04:19.39" />
                    <SPLIT distance="350" swimtime="00:05:04.69" />
                    <SPLIT distance="400" swimtime="00:05:50.65" />
                    <SPLIT distance="450" swimtime="00:06:36.65" />
                    <SPLIT distance="500" swimtime="00:07:21.57" />
                    <SPLIT distance="550" swimtime="00:08:07.27" />
                    <SPLIT distance="600" swimtime="00:08:52.34" />
                    <SPLIT distance="650" swimtime="00:09:37.08" />
                    <SPLIT distance="700" swimtime="00:10:21.47" />
                    <SPLIT distance="750" swimtime="00:11:06.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="637" reactiontime="+91" swimtime="00:00:36.94" resultid="9886" heatid="14203" lane="0" entrytime="00:00:36.50" entrycourse="SCM" />
                <RESULT eventid="8309" points="757" reactiontime="+81" swimtime="00:01:17.78" resultid="9887" heatid="14249" lane="9" entrytime="00:01:18.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="719" reactiontime="+95" swimtime="00:01:20.58" resultid="9888" heatid="14311" lane="5" entrytime="00:01:22.50" entrycourse="SCM" />
                <RESULT eventid="8582" status="DNS" swimtime="00:00:00.00" resultid="9889" heatid="14345" lane="4" entrytime="00:06:40.00" entrycourse="SCM" />
                <RESULT eventid="8662" points="641" reactiontime="+80" swimtime="00:03:03.90" resultid="9890" heatid="14369" lane="0" entrytime="00:03:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.78" />
                    <SPLIT distance="100" swimtime="00:02:17.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="9831">
              <RESULTS>
                <RESULT eventid="8213" points="506" reactiontime="+96" swimtime="00:00:43.51" resultid="9832" heatid="14201" lane="2" entrytime="00:00:43.50" entrycourse="SCM" />
                <RESULT eventid="8245" points="727" reactiontime="+111" swimtime="00:03:26.04" resultid="9833" heatid="14213" lane="3" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                    <SPLIT distance="150" swimtime="00:02:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="702" reactiontime="+105" swimtime="00:01:32.76" resultid="9834" heatid="14278" lane="6" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="493" reactiontime="+115" swimtime="00:01:35.00" resultid="9835" heatid="14311" lane="0" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="631" reactiontime="+98" swimtime="00:03:32.03" resultid="9836" heatid="14368" lane="1" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:42.71" />
                    <SPLIT distance="150" swimtime="00:02:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="593" reactiontime="+99" swimtime="00:00:42.27" resultid="9837" heatid="14383" lane="8" entrytime="00:00:40.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="9850">
              <RESULTS>
                <RESULT eventid="1075" points="312" reactiontime="+89" swimtime="00:00:39.57" resultid="9851" heatid="14145" lane="8" entrytime="00:00:39.76" entrycourse="SCM" />
                <RESULT eventid="1105" points="230" reactiontime="+83" swimtime="00:04:15.07" resultid="9852" heatid="14167" lane="3" entrytime="00:04:28.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                    <SPLIT distance="100" swimtime="00:02:03.51" />
                    <SPLIT distance="150" swimtime="00:03:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="218" reactiontime="+87" swimtime="00:01:57.67" resultid="9853" heatid="14246" lane="9" entrytime="00:01:54.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8341" points="136" reactiontime="+103" swimtime="00:05:09.93" resultid="9854" heatid="14258" lane="6" entrytime="00:05:07.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.52" />
                    <SPLIT distance="100" swimtime="00:02:23.49" />
                    <SPLIT distance="150" swimtime="00:03:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="196" reactiontime="+124" swimtime="00:02:04.18" resultid="9855" heatid="14309" lane="4" entrytime="00:02:06.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="226" reactiontime="+152" swimtime="00:09:16.97" resultid="9856" heatid="14344" lane="1" entrytime="00:09:04.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.29" />
                    <SPLIT distance="100" swimtime="00:02:21.55" />
                    <SPLIT distance="150" swimtime="00:03:33.68" />
                    <SPLIT distance="200" swimtime="00:04:45.53" />
                    <SPLIT distance="250" swimtime="00:06:07.11" />
                    <SPLIT distance="300" swimtime="00:07:27.59" />
                    <SPLIT distance="350" swimtime="00:08:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="113" reactiontime="+96" swimtime="00:02:19.22" resultid="9857" heatid="14354" lane="9" entrytime="00:02:10.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="209" reactiontime="+120" swimtime="00:04:26.93" resultid="9858" heatid="14367" lane="6" entrytime="00:04:30.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.38" />
                    <SPLIT distance="100" swimtime="00:02:11.18" />
                    <SPLIT distance="150" swimtime="00:03:21.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-05-25" firstname="Włodzimierz" gender="M" lastname="Łatecki" nation="POL" license="503105700032" athleteid="9838">
              <RESULTS>
                <RESULT eventid="1075" points="142" reactiontime="+104" swimtime="00:00:51.33" resultid="9839" heatid="14144" lane="5" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="8341" points="105" reactiontime="+100" swimtime="00:05:38.16" resultid="9840" heatid="14258" lane="3" entrytime="00:05:02.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.06" />
                    <SPLIT distance="100" swimtime="00:02:35.02" />
                    <SPLIT distance="150" swimtime="00:04:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="158" reactiontime="+120" swimtime="00:04:12.25" resultid="9841" heatid="14324" lane="0" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:03:05.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="108" reactiontime="+90" swimtime="00:05:32.40" resultid="9842" heatid="14367" lane="2" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:42.28" />
                    <SPLIT distance="150" swimtime="00:04:07.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="9865">
              <RESULTS>
                <RESULT eventid="1058" points="749" reactiontime="+93" swimtime="00:00:32.56" resultid="9866" heatid="14139" lane="3" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="8196" points="838" reactiontime="+77" swimtime="00:00:38.27" resultid="9867" heatid="14196" lane="8" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="8293" points="695" reactiontime="+92" swimtime="00:01:24.82" resultid="9868" heatid="14241" lane="4" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="829" reactiontime="+92" swimtime="00:00:34.85" resultid="9869" heatid="14288" lane="7" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="8470" points="750" reactiontime="+74" swimtime="00:01:25.98" resultid="9870" heatid="14306" lane="7" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8613" points="738" reactiontime="+99" swimtime="00:01:27.04" resultid="9871" heatid="14351" lane="5" entrytime="00:01:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="644" reactiontime="+96" swimtime="00:00:43.49" resultid="9872" heatid="14375" lane="7" entrytime="00:00:44.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="9910">
              <RESULTS>
                <RESULT eventid="1058" points="793" reactiontime="+93" swimtime="00:00:29.51" resultid="9911" heatid="14140" lane="4" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="8196" points="806" reactiontime="+91" swimtime="00:00:33.13" resultid="9912" heatid="14197" lane="1" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="8293" points="833" reactiontime="+95" swimtime="00:01:13.59" resultid="9913" heatid="14243" lane="1" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8470" points="833" reactiontime="+85" swimtime="00:01:14.37" resultid="9914" heatid="14307" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="830" reactiontime="+81" swimtime="00:02:43.59" resultid="9915" heatid="14365" lane="2" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:02:01.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="9901">
              <RESULTS>
                <RESULT eventid="1075" points="734" reactiontime="+82" swimtime="00:00:25.49" resultid="9902" heatid="14156" lane="2" entrytime="00:00:26.70" entrycourse="SCM" />
                <RESULT eventid="1105" points="669" reactiontime="+87" swimtime="00:02:25.56" resultid="9903" heatid="14172" lane="1" entrytime="00:02:35.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:07.76" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="732" reactiontime="+76" swimtime="00:00:57.06" resultid="9904" heatid="14234" lane="5" entrytime="00:00:58.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="680" reactiontime="+71" swimtime="00:01:04.59" resultid="9905" heatid="14253" lane="9" entrytime="00:01:07.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="741" reactiontime="+77" swimtime="00:01:10.72" resultid="9906" heatid="14283" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="9907" heatid="14298" lane="2" entrytime="00:00:29.55" entrycourse="SCM" />
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="9908" heatid="14357" lane="5" entrytime="00:01:10.20" entrycourse="SCM" />
                <RESULT eventid="8694" points="720" reactiontime="+69" swimtime="00:00:32.21" resultid="9909" heatid="14387" lane="4" entrytime="00:00:33.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" license="503105700049" athleteid="9916">
              <RESULTS>
                <RESULT eventid="1075" points="608" reactiontime="+84" swimtime="00:00:26.11" resultid="9917" heatid="14160" lane="0" entrytime="00:00:24.90" entrycourse="SCM" />
                <RESULT eventid="8454" points="564" reactiontime="+72" swimtime="00:00:27.68" resultid="9918" heatid="14301" lane="2" entrytime="00:00:26.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="9896">
              <RESULTS>
                <RESULT eventid="1090" points="827" reactiontime="+92" swimtime="00:02:39.85" resultid="9897" heatid="14165" lane="1" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="696" reactiontime="+91" swimtime="00:02:45.22" resultid="9898" heatid="14257" lane="6" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:00.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="836" reactiontime="+92" swimtime="00:00:31.86" resultid="9899" heatid="14289" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="8613" points="849" reactiontime="+83" swimtime="00:01:09.73" resultid="9900" heatid="14352" lane="6" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+68" swimtime="00:02:06.09" resultid="9932" heatid="14267" lane="2" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                    <SPLIT distance="100" swimtime="00:00:59.17" />
                    <SPLIT distance="150" swimtime="00:01:26.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9873" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="9925" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="9916" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="9850" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" swimtime="00:01:56.15" resultid="9933" heatid="14337" lane="4" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.04" />
                    <SPLIT distance="100" swimtime="00:01:04.17" />
                    <SPLIT distance="150" swimtime="00:01:29.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9873" number="1" />
                    <RELAYPOSITION athleteid="9850" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="9916" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="9925" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+96" swimtime="00:02:19.78" resultid="9934" heatid="14267" lane="6" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="150" swimtime="00:01:44.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9901" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="9831" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="9884" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="9919" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8550" reactiontime="+49" swimtime="00:02:09.81" resultid="9935" heatid="14337" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:44.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9919" number="1" reactiontime="+49" />
                    <RELAYPOSITION athleteid="9831" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="9884" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="9901" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+81" swimtime="00:02:18.60" resultid="9930" heatid="14264" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:36.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9910" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="9859" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="9896" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="9865" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8534" reactiontime="+95" swimtime="00:02:06.05" resultid="9931" heatid="14335" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:36.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9865" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="9859" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="9896" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="9910" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1120" reactiontime="+78" swimtime="00:01:53.72" resultid="9936" heatid="14177" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                    <SPLIT distance="100" swimtime="00:00:56.69" />
                    <SPLIT distance="150" swimtime="00:01:26.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9901" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="9896" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="9910" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="9916" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8710" reactiontime="+81" swimtime="00:02:01.66" resultid="9937" heatid="14392" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:35.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9910" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="9925" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="9896" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="9901" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="9938" heatid="14176" lane="9" entrytime="00:02:07.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9884" number="1" />
                    <RELAYPOSITION athleteid="9859" number="2" />
                    <RELAYPOSITION athleteid="9865" number="3" />
                    <RELAYPOSITION athleteid="9844" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="11224" name="Warsaw Masters Team">
          <CONTACT email="agnieszka.z.mazurkiewicz@gmail.com" name="Mazurkiewicz" phone="882185766" street="Agnieszka" />
          <ATHLETES>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="11336">
              <RESULTS>
                <RESULT eventid="1075" points="619" reactiontime="+75" swimtime="00:00:27.87" resultid="11337" heatid="14154" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1150" points="557" reactiontime="+81" swimtime="00:10:21.57" resultid="11338" heatid="14183" lane="5" entrytime="00:10:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                    <SPLIT distance="200" swimtime="00:02:31.11" />
                    <SPLIT distance="250" swimtime="00:03:10.39" />
                    <SPLIT distance="300" swimtime="00:03:49.72" />
                    <SPLIT distance="350" swimtime="00:04:29.17" />
                    <SPLIT distance="400" swimtime="00:05:08.57" />
                    <SPLIT distance="450" swimtime="00:05:47.62" />
                    <SPLIT distance="500" swimtime="00:06:27.33" />
                    <SPLIT distance="550" swimtime="00:07:07.19" />
                    <SPLIT distance="600" swimtime="00:07:47.18" />
                    <SPLIT distance="650" swimtime="00:08:26.93" />
                    <SPLIT distance="700" swimtime="00:09:06.66" />
                    <SPLIT distance="750" swimtime="00:09:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="513" reactiontime="+85" swimtime="00:00:33.91" resultid="11339" heatid="14203" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="8277" points="625" reactiontime="+87" swimtime="00:01:00.90" resultid="11340" heatid="14231" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="552" reactiontime="+78" swimtime="00:00:30.63" resultid="11341" heatid="14295" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="8518" points="585" reactiontime="+84" swimtime="00:02:15.12" resultid="11342" heatid="14330" lane="7" entrytime="00:02:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="535" reactiontime="+75" swimtime="00:04:56.29" resultid="11343" heatid="14400" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:49.15" />
                    <SPLIT distance="200" swimtime="00:02:27.31" />
                    <SPLIT distance="250" swimtime="00:03:05.37" />
                    <SPLIT distance="300" swimtime="00:03:43.27" />
                    <SPLIT distance="350" swimtime="00:04:21.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="11353">
              <RESULTS>
                <RESULT eventid="8245" points="702" reactiontime="+89" swimtime="00:02:38.08" resultid="11354" heatid="14216" lane="5" entrytime="00:02:43.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="638" reactiontime="+85" swimtime="00:01:11.22" resultid="11355" heatid="14283" lane="1" entrytime="00:01:13.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="380" reactiontime="+91" swimtime="00:00:31.57" resultid="11356" heatid="14296" lane="1" entrytime="00:00:31.13" />
                <RESULT eventid="8694" points="672" reactiontime="+76" swimtime="00:00:31.74" resultid="11357" heatid="14388" lane="6" entrytime="00:00:32.15" />
                <RESULT eventid="8742" points="497" reactiontime="+98" swimtime="00:05:03.24" resultid="11358" heatid="14400" lane="3" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:51.34" />
                    <SPLIT distance="200" swimtime="00:02:30.18" />
                    <SPLIT distance="250" swimtime="00:03:08.89" />
                    <SPLIT distance="300" swimtime="00:03:47.51" />
                    <SPLIT distance="350" swimtime="00:04:25.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="11281">
              <RESULTS>
                <RESULT eventid="1075" points="797" reactiontime="+73" swimtime="00:00:27.40" resultid="11282" heatid="14152" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1105" points="903" reactiontime="+79" swimtime="00:02:27.28" resultid="11283" heatid="14172" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:09.42" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="836" reactiontime="+85" swimtime="00:00:31.06" resultid="11284" heatid="14204" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="8309" points="891" reactiontime="+88" swimtime="00:01:07.70" resultid="11285" heatid="14251" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="766" reactiontime="+83" swimtime="00:00:29.92" resultid="11286" heatid="14298" lane="1" entrytime="00:00:29.99" />
                <RESULT eventid="8486" points="869" reactiontime="+89" swimtime="00:01:06.68" resultid="11287" heatid="14314" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="783" reactiontime="+78" swimtime="00:01:07.55" resultid="11288" heatid="14358" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="761" reactiontime="+91" swimtime="00:02:32.36" resultid="11289" heatid="14370" lane="9" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:54.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-28" firstname="Krzysztof" gender="M" lastname="Olszewski" nation="POL" athleteid="11320">
              <RESULTS>
                <RESULT eventid="1075" points="684" reactiontime="+81" swimtime="00:00:25.92" resultid="11321" heatid="14157" lane="3" entrytime="00:00:26.24" />
                <RESULT eventid="8213" points="583" reactiontime="+80" swimtime="00:00:29.98" resultid="11322" heatid="14206" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="8309" points="620" reactiontime="+78" swimtime="00:01:04.72" resultid="11323" heatid="14253" lane="6" entrytime="00:01:06.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="595" reactiontime="+86" swimtime="00:01:05.43" resultid="11324" heatid="14314" lane="5" entrytime="00:01:05.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="511" reactiontime="+77" swimtime="00:02:25.29" resultid="11325" heatid="14371" lane="9" entrytime="00:02:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="150" swimtime="00:01:47.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="11243">
              <RESULTS>
                <RESULT eventid="8293" points="1018" reactiontime="+75" swimtime="00:01:07.32" resultid="11244" heatid="14243" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski" eventid="8404" points="901" reactiontime="+80" swimtime="00:01:16.45" resultid="11245" heatid="14274" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="918" reactiontime="+74" swimtime="00:00:30.25" resultid="11246" heatid="14289" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="8678" points="927" reactiontime="+69" swimtime="00:00:34.75" resultid="11247" heatid="14378" lane="3" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="11256">
              <RESULTS>
                <RESULT eventid="1075" points="814" reactiontime="+91" swimtime="00:00:29.53" resultid="11257" heatid="14151" lane="1" entrytime="00:00:29.88" />
                <RESULT eventid="8213" points="847" reactiontime="+77" swimtime="00:00:35.21" resultid="11258" heatid="14202" lane="4" entrytime="00:00:36.95" />
                <RESULT eventid="8277" points="826" reactiontime="+103" swimtime="00:01:05.11" resultid="11259" heatid="14230" lane="2" entrytime="00:01:05.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="912" reactiontime="+80" swimtime="00:01:14.59" resultid="11260" heatid="14312" lane="7" entrytime="00:01:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="939" reactiontime="+96" swimtime="00:02:25.72" resultid="11261" heatid="14328" lane="6" entrytime="00:02:26.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="922" reactiontime="+70" swimtime="00:02:41.94" resultid="11262" heatid="14369" lane="6" entrytime="00:02:44.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:02:00.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-26" firstname="Ewa" gender="F" lastname="Galica" nation="POL" athleteid="13296">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="13297" heatid="14139" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="8261" points="532" reactiontime="+91" swimtime="00:01:10.89" resultid="13298" heatid="14222" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="511" reactiontime="+93" swimtime="00:00:35.26" resultid="13299" heatid="14287" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="8678" status="DNS" swimtime="00:00:00.00" resultid="13300" heatid="14374" lane="5" entrytime="00:00:45.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="11302">
              <RESULTS>
                <RESULT eventid="1075" points="809" reactiontime="+72" swimtime="00:00:24.68" resultid="11303" heatid="14160" lane="8" entrytime="00:00:24.89" />
                <RESULT eventid="8213" points="810" reactiontime="+83" swimtime="00:00:27.96" resultid="11304" heatid="14207" lane="2" entrytime="00:00:28.19" />
                <RESULT eventid="8309" points="768" reactiontime="+83" swimtime="00:01:02.01" resultid="11305" heatid="14255" lane="0" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="11306" heatid="14301" lane="8" entrytime="00:00:27.10" />
                <RESULT eventid="8486" status="DNS" swimtime="00:00:00.00" resultid="11307" heatid="14315" lane="1" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="11397">
              <RESULTS>
                <RESULT eventid="8277" points="719" reactiontime="+86" swimtime="00:00:54.22" resultid="11398" heatid="14224" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)., Z3" eventid="8309" reactiontime="+73" status="DSQ" swimtime="00:01:03.84" resultid="11399" heatid="14254" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="680" reactiontime="+76" swimtime="00:00:26.94" resultid="11400" heatid="14298" lane="3" entrytime="00:00:29.02" />
                <RESULT eventid="8518" points="788" reactiontime="+89" swimtime="00:02:01.81" resultid="11401" heatid="14322" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="100" swimtime="00:00:57.20" />
                    <SPLIT distance="150" swimtime="00:01:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="11402" heatid="14361" lane="7" entrytime="00:00:58.65" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="11403" heatid="14379" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-03" firstname="Karollina" gender="F" lastname="Kowalewska" nation="POL" athleteid="11349">
              <RESULTS>
                <RESULT eventid="8229" points="570" reactiontime="+88" swimtime="00:03:05.28" resultid="11350" heatid="14211" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:28.24" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="539" reactiontime="+98" swimtime="00:01:26.79" resultid="11351" heatid="14273" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="491" reactiontime="+84" swimtime="00:00:40.04" resultid="11352" heatid="14376" lane="4" entrytime="00:00:39.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="11330">
              <RESULTS>
                <RESULT eventid="8213" points="756" reactiontime="+66" swimtime="00:00:30.59" resultid="11331" heatid="14206" lane="9" entrytime="00:00:31.20" />
                <RESULT eventid="8309" points="653" reactiontime="+76" swimtime="00:01:09.21" resultid="11332" heatid="14252" lane="7" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="781" reactiontime="+81" swimtime="00:00:28.70" resultid="11333" heatid="14299" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="8518" points="627" reactiontime="+84" swimtime="00:02:14.01" resultid="11334" heatid="14331" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" status="DNS" swimtime="00:00:00.00" resultid="11335" heatid="14359" lane="7" entrytime="00:01:04.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="11372">
              <RESULTS>
                <RESULT eventid="1105" points="652" reactiontime="+96" swimtime="00:03:06.37" resultid="11373" heatid="14169" lane="5" entrytime="00:03:07.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                    <SPLIT distance="150" swimtime="00:02:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="864" reactiontime="+96" swimtime="00:03:11.19" resultid="11374" heatid="14215" lane="1" entrytime="00:03:07.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                    <SPLIT distance="150" swimtime="00:02:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="824" reactiontime="+77" swimtime="00:01:18.80" resultid="11375" heatid="14248" lane="6" entrytime="00:01:19.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="879" reactiontime="+89" swimtime="00:01:22.89" resultid="11376" heatid="14280" lane="5" entrytime="00:01:22.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="641" reactiontime="+91" swimtime="00:07:06.98" resultid="11377" heatid="14345" lane="8" entrytime="00:07:11.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                    <SPLIT distance="100" swimtime="00:01:47.16" />
                    <SPLIT distance="150" swimtime="00:03:41.88" />
                    <SPLIT distance="200" swimtime="00:04:35.62" />
                    <SPLIT distance="250" swimtime="00:05:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="825" reactiontime="+80" swimtime="00:00:37.19" resultid="11378" heatid="14386" lane="9" entrytime="00:00:36.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-02-17" firstname="Zbigniew" gender="M" lastname="Paluszak" nation="POL" athleteid="11270">
              <RESULTS>
                <RESULT eventid="8245" points="298" reactiontime="+86" swimtime="00:03:51.63" resultid="11271" heatid="14212" lane="4" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                    <SPLIT distance="100" swimtime="00:01:46.61" />
                    <SPLIT distance="150" swimtime="00:02:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G7 - Pływak znajdował się w pozycji na piersiach po opuszczaniu ściany nawrotowej., Z3" eventid="8309" reactiontime="+89" status="DSQ" swimtime="00:01:52.43" resultid="11272" heatid="14245" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="273" reactiontime="+96" swimtime="00:01:47.21" resultid="11273" heatid="14277" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="207" reactiontime="+93" swimtime="00:03:30.29" resultid="11274" heatid="14324" lane="7" entrytime="00:03:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:36.31" />
                    <SPLIT distance="150" swimtime="00:02:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="273" reactiontime="+90" swimtime="00:00:47.36" resultid="11275" heatid="14381" lane="0" entrytime="00:00:49.00" />
                <RESULT eventid="8742" points="184" reactiontime="+100" swimtime="00:07:37.93" resultid="11276" heatid="14403" lane="8" entrytime="00:07:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:41.99" />
                    <SPLIT distance="150" swimtime="00:02:41.92" />
                    <SPLIT distance="200" swimtime="00:03:40.57" />
                    <SPLIT distance="250" swimtime="00:04:39.14" />
                    <SPLIT distance="300" swimtime="00:05:40.63" />
                    <SPLIT distance="350" swimtime="00:06:39.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="11297">
              <RESULTS>
                <RESULT eventid="1165" points="427" reactiontime="+101" swimtime="00:32:07.40" resultid="11298" heatid="14188" lane="1" entrytime="00:34:09.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.78" />
                    <SPLIT distance="100" swimtime="00:02:05.43" />
                    <SPLIT distance="150" swimtime="00:03:11.15" />
                    <SPLIT distance="200" swimtime="00:04:16.47" />
                    <SPLIT distance="250" swimtime="00:05:21.78" />
                    <SPLIT distance="300" swimtime="00:06:26.53" />
                    <SPLIT distance="350" swimtime="00:07:30.57" />
                    <SPLIT distance="400" swimtime="00:08:35.04" />
                    <SPLIT distance="450" swimtime="00:09:39.55" />
                    <SPLIT distance="500" swimtime="00:10:43.86" />
                    <SPLIT distance="550" swimtime="00:11:48.37" />
                    <SPLIT distance="600" swimtime="00:12:52.19" />
                    <SPLIT distance="650" swimtime="00:13:56.64" />
                    <SPLIT distance="700" swimtime="00:15:01.61" />
                    <SPLIT distance="750" swimtime="00:16:05.56" />
                    <SPLIT distance="800" swimtime="00:17:10.37" />
                    <SPLIT distance="850" swimtime="00:18:15.06" />
                    <SPLIT distance="900" swimtime="00:19:20.10" />
                    <SPLIT distance="950" swimtime="00:20:23.91" />
                    <SPLIT distance="1000" swimtime="00:21:27.97" />
                    <SPLIT distance="1050" swimtime="00:22:33.10" />
                    <SPLIT distance="1100" swimtime="00:23:37.50" />
                    <SPLIT distance="1150" swimtime="00:24:41.54" />
                    <SPLIT distance="1200" swimtime="00:25:45.22" />
                    <SPLIT distance="1250" swimtime="00:26:48.89" />
                    <SPLIT distance="1300" swimtime="00:27:52.96" />
                    <SPLIT distance="1350" swimtime="00:28:56.49" />
                    <SPLIT distance="1400" swimtime="00:29:51.39" />
                    <SPLIT distance="1450" swimtime="00:31:06.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8261" points="200" swimtime="00:02:01.35" resultid="11299" heatid="14218" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" status="DNS" swimtime="00:00:00.00" resultid="11300" heatid="14317" lane="1" entrytime="00:04:15.00" />
                <RESULT eventid="8726" points="288" swimtime="00:08:53.39" resultid="11301" heatid="14396" lane="8" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.02" />
                    <SPLIT distance="100" swimtime="00:02:07.75" />
                    <SPLIT distance="150" swimtime="00:03:14.61" />
                    <SPLIT distance="200" swimtime="00:04:21.60" />
                    <SPLIT distance="250" swimtime="00:05:29.09" />
                    <SPLIT distance="300" swimtime="00:06:36.38" />
                    <SPLIT distance="350" swimtime="00:07:45.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-11" firstname="Bolek" gender="M" lastname="Szuter" nation="POL" athleteid="11386">
              <RESULTS>
                <RESULT eventid="1075" points="805" reactiontime="+83" swimtime="00:00:25.65" resultid="11387" heatid="14160" lane="1" entrytime="00:00:24.88" />
                <RESULT comment="Rekord Polski" eventid="8277" points="907" reactiontime="+76" swimtime="00:00:54.67" resultid="11388" heatid="14236" lane="6" entrytime="00:00:55.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="819" reactiontime="+77" swimtime="00:00:28.26" resultid="11389" heatid="14300" lane="7" entrytime="00:00:27.77" />
                <RESULT comment="Rekord Polski" eventid="8518" points="828" reactiontime="+83" swimtime="00:02:02.17" resultid="11390" heatid="14332" lane="6" entrytime="00:02:06.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="150" swimtime="00:01:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8630" points="726" reactiontime="+78" swimtime="00:01:05.42" resultid="11391" heatid="14358" lane="2" entrytime="00:01:07.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="11326">
              <RESULTS>
                <RESULT eventid="8213" points="628" reactiontime="+83" swimtime="00:00:30.93" resultid="11327" heatid="14206" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="8518" points="580" reactiontime="+84" swimtime="00:02:07.70" resultid="11328" heatid="14332" lane="1" entrytime="00:02:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                    <SPLIT distance="150" swimtime="00:01:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="616" reactiontime="+77" swimtime="00:04:42.32" resultid="11329" heatid="14399" lane="0" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:07.71" />
                    <SPLIT distance="150" swimtime="00:01:44.47" />
                    <SPLIT distance="200" swimtime="00:02:21.69" />
                    <SPLIT distance="250" swimtime="00:02:57.91" />
                    <SPLIT distance="300" swimtime="00:03:33.15" />
                    <SPLIT distance="350" swimtime="00:04:08.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-04-14" firstname="Wiesław" gender="M" lastname="Załuski" nation="POL" athleteid="11392">
              <RESULTS>
                <RESULT eventid="1075" points="740" reactiontime="+105" swimtime="00:00:30.48" resultid="11393" heatid="14149" lane="2" entrytime="00:00:30.55" />
                <RESULT eventid="8213" points="841" reactiontime="+62" swimtime="00:00:35.29" resultid="11394" heatid="14203" lane="8" entrytime="00:00:36.20" />
                <RESULT eventid="8309" points="854" reactiontime="+111" swimtime="00:01:17.87" resultid="11395" heatid="14248" lane="2" entrytime="00:01:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="750" reactiontime="+67" swimtime="00:01:19.62" resultid="11396" heatid="14312" lane="8" entrytime="00:01:20.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-18" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="11359">
              <RESULTS>
                <RESULT eventid="1058" points="517" reactiontime="+110" swimtime="00:00:41.54" resultid="11360" heatid="14136" lane="5" entrytime="00:00:39.41" />
                <RESULT eventid="8196" points="563" reactiontime="+87" swimtime="00:00:50.63" resultid="11361" heatid="14194" lane="1" entrytime="00:00:48.75" />
                <RESULT eventid="8470" points="471" reactiontime="+80" swimtime="00:01:54.49" resultid="11362" heatid="14305" lane="0" entrytime="00:01:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-10" firstname="Łukasz" gender="M" lastname="Rybiński" nation="POL" athleteid="11277">
              <RESULTS>
                <RESULT eventid="1075" points="506" reactiontime="+93" swimtime="00:00:29.80" resultid="11278" heatid="14149" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="8277" points="479" reactiontime="+94" swimtime="00:01:06.54" resultid="11279" heatid="14228" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="463" reactiontime="+97" swimtime="00:01:24.78" resultid="11280" heatid="14279" lane="6" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="11315">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="11316" heatid="14172" lane="9" entrytime="00:02:37.20" />
                <RESULT eventid="8277" status="DNS" swimtime="00:00:00.00" resultid="11317" heatid="14232" lane="1" entrytime="00:01:02.50" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="11318" heatid="14330" lane="3" entrytime="00:02:16.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="11344">
              <RESULTS>
                <RESULT eventid="1058" points="590" reactiontime="+78" swimtime="00:00:32.39" resultid="11345" heatid="14138" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="8229" points="520" reactiontime="+87" swimtime="00:03:26.49" resultid="11346" heatid="14209" lane="4" entrytime="00:03:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                    <SPLIT distance="150" swimtime="00:02:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="579" reactiontime="+84" swimtime="00:01:30.79" resultid="11347" heatid="14271" lane="4" entrytime="00:01:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="594" reactiontime="+86" swimtime="00:00:40.83" resultid="11348" heatid="14375" lane="8" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-10-11" firstname="Grzegorz" gender="M" lastname="Matyszewski" nation="POL" athleteid="11363">
              <RESULTS>
                <RESULT eventid="1075" points="399" reactiontime="+69" swimtime="00:00:32.42" resultid="11364" heatid="14148" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1105" points="359" reactiontime="+74" swimtime="00:03:10.31" resultid="11365" heatid="14169" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:32.56" />
                    <SPLIT distance="150" swimtime="00:02:22.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="455" reactiontime="+93" swimtime="00:03:11.92" resultid="11366" heatid="14215" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:20.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="368" reactiontime="+84" swimtime="00:01:23.80" resultid="11367" heatid="14247" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="455" reactiontime="+76" swimtime="00:01:25.87" resultid="11368" heatid="14280" lane="9" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="244" reactiontime="+89" swimtime="00:03:03.46" resultid="11369" heatid="14325" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:28.08" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="537" reactiontime="+71" swimtime="00:00:37.36" resultid="11370" heatid="14384" lane="0" entrytime="00:00:38.50" />
                <RESULT eventid="8742" points="224" reactiontime="+80" swimtime="00:06:44.65" resultid="11371" heatid="14403" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:30.98" />
                    <SPLIT distance="150" swimtime="00:02:20.30" />
                    <SPLIT distance="200" swimtime="00:03:11.11" />
                    <SPLIT distance="250" swimtime="00:04:02.39" />
                    <SPLIT distance="300" swimtime="00:04:56.28" />
                    <SPLIT distance="350" swimtime="00:05:50.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-07" firstname="Daniel" gender="M" lastname="Julian Aguilar" nation="POL" athleteid="11248">
              <RESULTS>
                <RESULT eventid="1075" points="666" reactiontime="+79" swimtime="00:00:26.33" resultid="11249" heatid="14156" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1105" points="585" reactiontime="+67" swimtime="00:02:32.22" resultid="11250" heatid="14173" lane="7" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" points="625" reactiontime="+69" swimtime="00:00:30.48" resultid="11251" heatid="14207" lane="9" entrytime="00:00:29.80" />
                <RESULT eventid="8277" points="714" reactiontime="+78" swimtime="00:00:57.53" resultid="11252" heatid="14234" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8518" points="599" reactiontime="+76" swimtime="00:02:12.21" resultid="11253" heatid="14331" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="559" reactiontime="+65" swimtime="00:02:27.52" resultid="11254" heatid="14371" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="585" reactiontime="+69" swimtime="00:04:49.73" resultid="11255" heatid="14399" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:44.61" />
                    <SPLIT distance="200" swimtime="00:02:21.71" />
                    <SPLIT distance="250" swimtime="00:02:58.66" />
                    <SPLIT distance="300" swimtime="00:03:35.87" />
                    <SPLIT distance="350" swimtime="00:04:13.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="11290">
              <RESULTS>
                <RESULT eventid="1075" points="309" reactiontime="+98" swimtime="00:00:38.57" resultid="11291" heatid="14145" lane="6" entrytime="00:00:39.10" />
                <RESULT eventid="1150" points="412" reactiontime="+116" swimtime="00:13:10.99" resultid="11292" heatid="14185" lane="0" entrytime="00:13:40.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:33.10" />
                    <SPLIT distance="150" swimtime="00:02:22.81" />
                    <SPLIT distance="200" swimtime="00:03:13.20" />
                    <SPLIT distance="250" swimtime="00:04:03.24" />
                    <SPLIT distance="300" swimtime="00:04:53.80" />
                    <SPLIT distance="350" swimtime="00:05:44.35" />
                    <SPLIT distance="400" swimtime="00:06:34.89" />
                    <SPLIT distance="450" swimtime="00:07:25.07" />
                    <SPLIT distance="500" swimtime="00:08:16.28" />
                    <SPLIT distance="550" swimtime="00:09:05.80" />
                    <SPLIT distance="600" swimtime="00:09:55.19" />
                    <SPLIT distance="650" swimtime="00:10:46.05" />
                    <SPLIT distance="700" swimtime="00:11:36.05" />
                    <SPLIT distance="750" swimtime="00:12:24.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8277" points="306" reactiontime="+117" swimtime="00:01:26.09" resultid="11293" heatid="14226" lane="0" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="208" reactiontime="+108" swimtime="00:00:48.10" resultid="11294" heatid="14291" lane="3" entrytime="00:00:46.76" />
                <RESULT eventid="8518" points="363" reactiontime="+112" swimtime="00:03:03.68" resultid="11295" heatid="14325" lane="8" entrytime="00:03:05.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8742" points="391" reactiontime="+102" swimtime="00:06:27.75" resultid="11296" heatid="14402" lane="9" entrytime="00:06:38.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.58" />
                    <SPLIT distance="100" swimtime="00:02:22.25" />
                    <SPLIT distance="200" swimtime="00:03:11.76" />
                    <SPLIT distance="250" swimtime="00:04:01.07" />
                    <SPLIT distance="300" swimtime="00:04:51.55" />
                    <SPLIT distance="350" swimtime="00:05:40.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="11379">
              <RESULTS>
                <RESULT eventid="1075" points="142" reactiontime="+114" swimtime="00:01:03.64" resultid="11380" heatid="14143" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="8213" points="201" reactiontime="+77" swimtime="00:01:14.22" resultid="11381" heatid="14199" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="8309" points="205" reactiontime="+130" swimtime="00:02:30.00" resultid="11382" heatid="14245" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="179" reactiontime="+127" swimtime="00:02:51.65" resultid="11383" heatid="14275" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="126" reactiontime="+103" swimtime="00:03:03.19" resultid="11384" heatid="14309" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="320" reactiontime="+122" swimtime="00:01:03.86" resultid="11385" heatid="14380" lane="9" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="11234">
              <RESULTS>
                <RESULT eventid="1075" points="492" reactiontime="+84" swimtime="00:00:29.13" resultid="11235" heatid="14153" lane="0" entrytime="00:00:28.57" />
                <RESULT eventid="1105" points="504" reactiontime="+93" swimtime="00:02:39.87" resultid="11236" heatid="14172" lane="8" entrytime="00:02:35.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:02:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8213" status="DNS" swimtime="00:00:00.00" resultid="11237" heatid="14203" lane="5" entrytime="00:00:34.77" />
                <RESULT eventid="8309" status="DNS" swimtime="00:00:00.00" resultid="11238" heatid="14251" lane="7" entrytime="00:01:11.15" />
                <RESULT eventid="8454" status="DNS" swimtime="00:00:00.00" resultid="11239" heatid="14297" lane="0" entrytime="00:00:30.53" />
                <RESULT eventid="8518" status="DNS" swimtime="00:00:00.00" resultid="11240" heatid="14330" lane="9" entrytime="00:02:18.50" />
                <RESULT eventid="8694" status="DNS" swimtime="00:00:00.00" resultid="11241" heatid="14386" lane="7" entrytime="00:00:35.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="11308">
              <RESULTS>
                <RESULT eventid="1090" points="504" reactiontime="+89" swimtime="00:02:59.64" resultid="11309" heatid="14162" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:24.70" />
                    <SPLIT distance="150" swimtime="00:02:17.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="564" reactiontime="+84" swimtime="00:11:30.30" resultid="11310" heatid="14178" lane="8" entrytime="00:11:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:00.78" />
                    <SPLIT distance="200" swimtime="00:02:44.03" />
                    <SPLIT distance="250" swimtime="00:03:27.14" />
                    <SPLIT distance="300" swimtime="00:04:10.59" />
                    <SPLIT distance="350" swimtime="00:04:53.90" />
                    <SPLIT distance="400" swimtime="00:05:37.77" />
                    <SPLIT distance="450" swimtime="00:06:21.83" />
                    <SPLIT distance="500" swimtime="00:07:06.24" />
                    <SPLIT distance="550" swimtime="00:07:50.99" />
                    <SPLIT distance="600" swimtime="00:08:35.03" />
                    <SPLIT distance="650" swimtime="00:09:19.30" />
                    <SPLIT distance="700" swimtime="00:10:04.12" />
                    <SPLIT distance="750" swimtime="00:10:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="484" reactiontime="+91" swimtime="00:01:22.52" resultid="11311" heatid="14242" lane="0" entrytime="00:01:20.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8325" points="330" reactiontime="+100" swimtime="00:03:26.89" resultid="11312" heatid="14256" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="519" reactiontime="+86" swimtime="00:00:35.06" resultid="11313" heatid="14288" lane="4" entrytime="00:00:33.90" />
                <RESULT eventid="8566" status="DNS" swimtime="00:00:00.00" resultid="11314" heatid="14342" lane="0" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-27" firstname="Wojciech" gender="M" lastname="Kossowski" nation="POL" athleteid="11263">
              <RESULTS>
                <RESULT eventid="1105" points="452" reactiontime="+120" swimtime="00:03:23.77" resultid="11264" heatid="14168" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:43.55" />
                    <SPLIT distance="150" swimtime="00:02:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8245" points="511" reactiontime="+126" swimtime="00:03:27.46" resultid="11265" heatid="14213" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:40.38" />
                    <SPLIT distance="150" swimtime="00:02:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8309" points="459" reactiontime="+130" swimtime="00:01:31.86" resultid="11266" heatid="14247" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="522" reactiontime="+123" swimtime="00:01:31.74" resultid="11267" heatid="14278" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8582" points="432" reactiontime="+129" swimtime="00:07:28.93" resultid="11268" heatid="14345" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                    <SPLIT distance="100" swimtime="00:01:47.55" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                    <SPLIT distance="200" swimtime="00:03:51.96" />
                    <SPLIT distance="250" swimtime="00:04:51.10" />
                    <SPLIT distance="300" swimtime="00:05:48.74" />
                    <SPLIT distance="350" swimtime="00:06:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="502" reactiontime="+112" swimtime="00:00:41.18" resultid="11269" heatid="14382" lane="7" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="11225">
              <RESULTS>
                <RESULT eventid="1090" points="425" reactiontime="+92" swimtime="00:03:19.61" resultid="11226" heatid="14163" lane="6" entrytime="00:03:20.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="150" swimtime="00:02:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="390" reactiontime="+102" swimtime="00:13:07.68" resultid="11227" heatid="14179" lane="0" entrytime="00:13:46.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:18.10" />
                    <SPLIT distance="200" swimtime="00:03:07.17" />
                    <SPLIT distance="250" swimtime="00:03:56.76" />
                    <SPLIT distance="300" swimtime="00:04:46.53" />
                    <SPLIT distance="350" swimtime="00:05:36.58" />
                    <SPLIT distance="400" swimtime="00:06:27.29" />
                    <SPLIT distance="450" swimtime="00:07:18.18" />
                    <SPLIT distance="500" swimtime="00:08:08.23" />
                    <SPLIT distance="550" swimtime="00:08:58.37" />
                    <SPLIT distance="600" swimtime="00:09:48.85" />
                    <SPLIT distance="650" swimtime="00:10:39.58" />
                    <SPLIT distance="700" swimtime="00:11:30.04" />
                    <SPLIT distance="750" swimtime="00:12:19.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="564" reactiontime="+106" swimtime="00:03:26.21" resultid="11228" heatid="14210" lane="0" entrytime="00:03:35.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8293" points="438" reactiontime="+94" swimtime="00:01:31.14" resultid="11229" heatid="14240" lane="1" entrytime="00:01:33.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="542" reactiontime="+91" swimtime="00:01:35.41" resultid="11230" heatid="14272" lane="7" entrytime="00:01:36.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="382" reactiontime="+110" swimtime="00:02:59.76" resultid="11231" heatid="14318" lane="4" entrytime="00:03:05.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:26.35" />
                    <SPLIT distance="150" swimtime="00:02:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="600" reactiontime="+86" swimtime="00:00:41.67" resultid="11232" heatid="14376" lane="9" entrytime="00:00:42.31" />
                <RESULT eventid="8726" points="408" reactiontime="+86" swimtime="00:06:22.65" resultid="11233" heatid="14395" lane="7" entrytime="00:06:17.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                    <SPLIT distance="150" swimtime="00:02:17.00" />
                    <SPLIT distance="200" swimtime="00:03:05.87" />
                    <SPLIT distance="250" swimtime="00:03:54.57" />
                    <SPLIT distance="300" swimtime="00:04:44.18" />
                    <SPLIT distance="350" swimtime="00:05:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+67" swimtime="00:01:57.78" resultid="11404" heatid="14267" lane="4" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:01.70" />
                    <SPLIT distance="150" swimtime="00:01:31.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11248" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="11353" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="11336" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="11320" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+84" swimtime="00:02:01.14" resultid="11405" heatid="14267" lane="5" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:33.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11302" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="11372" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="11386" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="11281" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski. Pierwsza zmiana" eventid="8550" reactiontime="+75" swimtime="00:01:42.00" resultid="11406" heatid="14339" lane="7" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.40" />
                    <SPLIT distance="100" swimtime="00:00:50.72" />
                    <SPLIT distance="150" swimtime="00:01:16.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11302" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="11326" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="11320" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="11248" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT comment="Rekord Polski, pierwsz zmiana" eventid="8550" reactiontime="+80" swimtime="00:01:48.39" resultid="11407" heatid="14338" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                    <SPLIT distance="100" swimtime="00:00:53.07" />
                    <SPLIT distance="150" swimtime="00:01:20.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11386" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="11281" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="11336" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="11330" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="9497" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="9513">
              <RESULTS>
                <RESULT eventid="8229" points="294" reactiontime="+123" swimtime="00:05:01.70" resultid="9514" heatid="14208" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.48" />
                    <SPLIT distance="100" swimtime="00:02:24.66" />
                    <SPLIT distance="150" swimtime="00:03:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="250" reactiontime="+101" swimtime="00:02:24.51" resultid="9515" heatid="14270" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="306" reactiontime="+100" swimtime="00:01:01.18" resultid="9516" heatid="14373" lane="7" entrytime="00:00:58.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="502611100004" athleteid="9538">
              <RESULTS>
                <RESULT eventid="8213" points="533" reactiontime="+73" swimtime="00:00:42.76" resultid="9539" heatid="14201" lane="6" entrytime="00:00:43.35" />
                <RESULT eventid="8486" points="440" reactiontime="+75" swimtime="00:01:38.64" resultid="9540" heatid="14311" lane="9" entrytime="00:01:39.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="573" reactiontime="+71" swimtime="00:03:38.95" resultid="9541" heatid="14368" lane="0" entrytime="00:03:41.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                    <SPLIT distance="100" swimtime="00:01:43.71" />
                    <SPLIT distance="150" swimtime="00:02:42.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-02-18" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" license="502611100006" athleteid="9498">
              <RESULTS>
                <RESULT eventid="1058" points="538" reactiontime="+75" swimtime="00:00:39.64" resultid="9499" heatid="14137" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="8196" points="859" reactiontime="+85" swimtime="00:00:42.11" resultid="9500" heatid="14195" lane="1" entrytime="00:00:42.50" />
                <RESULT eventid="8438" points="540" reactiontime="+89" swimtime="00:00:44.79" resultid="9501" heatid="14286" lane="6" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="102611600021" athleteid="9525">
              <RESULTS>
                <RESULT eventid="8213" points="383" reactiontime="+84" swimtime="00:00:40.41" resultid="9526" heatid="14202" lane="0" entrytime="00:00:40.24" />
                <RESULT eventid="8277" points="528" reactiontime="+98" swimtime="00:01:11.78" resultid="9527" heatid="14228" lane="0" entrytime="00:01:12.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="420" reactiontime="+93" swimtime="00:01:26.42" resultid="9528" heatid="14311" lane="3" entrytime="00:01:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="430" reactiontime="+80" swimtime="00:03:09.72" resultid="9529" heatid="14368" lane="6" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:31.14" />
                    <SPLIT distance="150" swimtime="00:02:20.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="102611600023" athleteid="9517">
              <RESULTS>
                <RESULT eventid="1058" points="751" reactiontime="+85" swimtime="00:00:38.03" resultid="9518" heatid="14137" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1090" points="709" reactiontime="+86" swimtime="00:03:55.81" resultid="9519" heatid="14162" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.95" />
                    <SPLIT distance="150" swimtime="00:03:07.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8196" points="753" reactiontime="+76" swimtime="00:00:47.96" resultid="9520" heatid="14194" lane="6" entrytime="00:00:47.61" />
                <RESULT eventid="8293" points="689" reactiontime="+95" swimtime="00:01:46.23" resultid="9521" heatid="14239" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="506" reactiontime="+82" swimtime="00:00:52.12" resultid="9522" heatid="14286" lane="8" entrytime="00:00:53.00" />
                <RESULT eventid="8502" points="686" swimtime="00:03:24.30" resultid="9523" heatid="14317" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8646" points="685" reactiontime="+70" swimtime="00:03:49.88" resultid="9524" heatid="14363" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.73" />
                    <SPLIT distance="100" swimtime="00:01:55.46" />
                    <SPLIT distance="150" swimtime="00:02:54.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-20" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="102611600015" athleteid="9530">
              <RESULTS>
                <RESULT eventid="1075" points="581" reactiontime="+74" swimtime="00:00:33.05" resultid="9531" heatid="14148" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="8309" points="438" reactiontime="+90" swimtime="00:01:37.25" resultid="9532" heatid="14247" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="515" reactiontime="+100" swimtime="00:00:38.12" resultid="9533" heatid="14293" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="102611600019" athleteid="9506">
              <RESULTS>
                <RESULT eventid="1135" points="579" reactiontime="+108" swimtime="00:16:42.05" resultid="9507" heatid="14180" lane="1" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.82" />
                    <SPLIT distance="100" swimtime="00:01:53.50" />
                    <SPLIT distance="150" swimtime="00:02:56.01" />
                    <SPLIT distance="200" swimtime="00:03:59.52" />
                    <SPLIT distance="250" swimtime="00:05:02.33" />
                    <SPLIT distance="300" swimtime="00:06:05.67" />
                    <SPLIT distance="350" swimtime="00:07:09.61" />
                    <SPLIT distance="400" swimtime="00:08:12.24" />
                    <SPLIT distance="450" swimtime="00:09:14.74" />
                    <SPLIT distance="500" swimtime="00:10:19.48" />
                    <SPLIT distance="550" swimtime="00:11:23.98" />
                    <SPLIT distance="600" swimtime="00:12:26.80" />
                    <SPLIT distance="650" swimtime="00:13:30.96" />
                    <SPLIT distance="700" swimtime="00:14:36.23" />
                    <SPLIT distance="750" swimtime="00:15:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="613" reactiontime="+111" swimtime="00:04:14.29" resultid="9508" heatid="14208" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.56" />
                    <SPLIT distance="100" swimtime="00:02:03.13" />
                    <SPLIT distance="150" swimtime="00:03:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="634" reactiontime="+104" swimtime="00:01:54.96" resultid="9509" heatid="14271" lane="8" entrytime="00:01:54.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8438" points="499" reactiontime="+113" swimtime="00:00:52.38" resultid="9510" heatid="14286" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="8613" points="699" reactiontime="+95" swimtime="00:02:00.51" resultid="9511" heatid="14350" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="585" reactiontime="+95" swimtime="00:00:56.37" resultid="9512" heatid="14373" lane="4" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="102611600024" athleteid="9549">
              <RESULTS>
                <RESULT eventid="1058" points="334" reactiontime="+95" swimtime="00:00:48.02" resultid="9550" heatid="14135" lane="6" entrytime="00:00:51.00" />
                <RESULT eventid="8196" points="420" reactiontime="+104" swimtime="00:00:55.80" resultid="9551" heatid="14193" lane="4" entrytime="00:00:56.00" />
                <RESULT eventid="8470" points="367" reactiontime="+103" swimtime="00:02:04.34" resultid="9552" heatid="14304" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:06.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="472" reactiontime="+103" swimtime="00:00:55.42" resultid="9553" heatid="14373" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="8293" points="333" reactiontime="+125" swimtime="00:02:00.27" resultid="13220" heatid="14239" lane="1" entrytime="00:01:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="102611600016" athleteid="9542">
              <RESULTS>
                <RESULT eventid="1135" points="818" reactiontime="+79" swimtime="00:10:15.54" resultid="9543" heatid="14178" lane="3" entrytime="00:10:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:13.48" />
                    <SPLIT distance="150" swimtime="00:01:52.03" />
                    <SPLIT distance="200" swimtime="00:02:30.53" />
                    <SPLIT distance="250" swimtime="00:03:09.24" />
                    <SPLIT distance="300" swimtime="00:03:47.90" />
                    <SPLIT distance="350" swimtime="00:04:26.72" />
                    <SPLIT distance="400" swimtime="00:05:05.84" />
                    <SPLIT distance="450" swimtime="00:05:44.67" />
                    <SPLIT distance="500" swimtime="00:06:23.52" />
                    <SPLIT distance="550" swimtime="00:07:02.46" />
                    <SPLIT distance="600" swimtime="00:07:41.52" />
                    <SPLIT distance="650" swimtime="00:08:20.79" />
                    <SPLIT distance="700" swimtime="00:08:59.76" />
                    <SPLIT distance="750" swimtime="00:09:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8229" points="822" reactiontime="+92" swimtime="00:03:01.85" resultid="9544" heatid="14211" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:13.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8404" points="849" reactiontime="+84" swimtime="00:01:22.15" resultid="9545" heatid="14274" lane="8" entrytime="00:01:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8502" points="743" reactiontime="+100" swimtime="00:02:24.00" resultid="9546" heatid="14321" lane="8" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:10.07" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8678" points="750" reactiontime="+81" swimtime="00:00:38.69" resultid="9547" heatid="14377" lane="0" entrytime="00:00:38.50" />
                <RESULT eventid="8726" points="829" reactiontime="+84" swimtime="00:05:02.07" resultid="9548" heatid="14393" lane="2" entrytime="00:04:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:30.17" />
                    <SPLIT distance="250" swimtime="00:03:08.72" />
                    <SPLIT distance="300" swimtime="00:03:47.35" />
                    <SPLIT distance="350" swimtime="00:04:25.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="102611600014" athleteid="9534">
              <RESULTS>
                <RESULT eventid="1075" points="309" reactiontime="+113" swimtime="00:00:42.89" resultid="9535" heatid="14145" lane="1" entrytime="00:00:39.50" />
                <RESULT eventid="8309" points="269" reactiontime="+94" swimtime="00:02:01.38" resultid="9536" heatid="14246" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8454" points="200" reactiontime="+106" swimtime="00:00:55.26" resultid="9537" heatid="14291" lane="5" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="102611600018" athleteid="9502">
              <RESULTS>
                <RESULT eventid="8245" points="646" reactiontime="+110" swimtime="00:03:46.12" resultid="9503" heatid="14213" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                    <SPLIT distance="100" swimtime="00:01:50.61" />
                    <SPLIT distance="150" swimtime="00:02:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8406" points="590" reactiontime="+86" swimtime="00:01:43.39" resultid="9504" heatid="14277" lane="7" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8694" points="573" reactiontime="+94" swimtime="00:00:47.18" resultid="9505" heatid="14381" lane="2" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="8373" reactiontime="+69" swimtime="00:02:54.68" resultid="9556" heatid="14266" lane="9" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:32.11" />
                    <SPLIT distance="150" swimtime="00:02:12.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9538" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="9502" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="9530" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="9534" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="8550" reactiontime="+110" swimtime="00:02:40.98" resultid="9558" heatid="14336" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:00.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9534" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="9538" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="9502" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="9530" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="8357" reactiontime="+87" swimtime="00:03:09.01" resultid="9555" heatid="14263" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                    <SPLIT distance="150" swimtime="00:02:30.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9498" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="9549" number="2" />
                    <RELAYPOSITION athleteid="9506" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="9517" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="8534" reactiontime="+126" swimtime="00:03:01.30" resultid="9557" heatid="14335" lane="0" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:40.51" />
                    <SPLIT distance="150" swimtime="00:02:21.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9549" number="1" reactiontime="+126" />
                    <RELAYPOSITION athleteid="9506" number="2" />
                    <RELAYPOSITION athleteid="9498" number="3" />
                    <RELAYPOSITION athleteid="9517" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1120" reactiontime="+89" status="DSQ" swimtime="00:02:36.33" resultid="9554" heatid="14175" lane="2" entrytime="00:02:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9517" number="1" reactiontime="+89" status="DSQ" />
                    <RELAYPOSITION athleteid="9498" number="2" reactiontime="-13" status="DSQ" />
                    <RELAYPOSITION athleteid="9534" number="3" reactiontime="+55" status="DSQ" />
                    <RELAYPOSITION athleteid="9530" number="4" reactiontime="+34" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="8710" reactiontime="+75" swimtime="00:03:03.65" resultid="9559" heatid="14390" lane="6" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:41.39" />
                    <SPLIT distance="150" swimtime="00:02:20.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9517" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="9549" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="9530" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="9534" number="4" reactiontime="+87" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="13221" name="WKS Śląsk Wrocław">
          <CONTACT email="marrot68@wp.pl" name="Rother Marek" phone="785209045" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="13222">
              <RESULTS>
                <RESULT eventid="8213" points="971" reactiontime="+74" swimtime="00:00:29.54" resultid="13223" heatid="14206" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="8309" points="941" reactiontime="+73" swimtime="00:01:06.47" resultid="13224" heatid="14252" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8486" points="923" reactiontime="+74" swimtime="00:01:05.35" resultid="13225" heatid="14314" lane="4" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="8662" points="970" reactiontime="+66" swimtime="00:02:20.53" resultid="13226" heatid="14371" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:43.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

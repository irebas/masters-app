<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Michał Derewecki" version="11.71436">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="Zimowe Otwarte Mistrzostwa Polski w Pływaniu w Kategoriach MASTERS POZNAŃ 2021" course="SCM" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-12-12" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Poznań" nation="POL" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <QUALIFY from="2020-03-01" until="2021-12-10" />
      <SESSIONS>
        <SESSION date="2021-12-11" daytime="09:00" endtime="12:44" number="1">
          <EVENTS>
            <EVENT eventid="1059" daytime="09:00" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2989" />
                    <RANKING order="2" place="2" resultid="5726" />
                    <RANKING order="3" place="3" resultid="5437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4359" />
                    <RANKING order="2" place="2" resultid="3428" />
                    <RANKING order="3" place="3" resultid="3878" />
                    <RANKING order="4" place="4" resultid="4896" />
                    <RANKING order="5" place="5" resultid="3345" />
                    <RANKING order="6" place="6" resultid="4343" />
                    <RANKING order="7" place="7" resultid="3003" />
                    <RANKING order="8" place="8" resultid="5077" />
                    <RANKING order="9" place="9" resultid="4746" />
                    <RANKING order="10" place="-1" resultid="3424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4802" />
                    <RANKING order="2" place="2" resultid="5072" />
                    <RANKING order="3" place="3" resultid="3680" />
                    <RANKING order="4" place="4" resultid="3530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5296" />
                    <RANKING order="2" place="2" resultid="3658" />
                    <RANKING order="3" place="3" resultid="3173" />
                    <RANKING order="4" place="4" resultid="3724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4569" />
                    <RANKING order="2" place="2" resultid="4737" />
                    <RANKING order="3" place="3" resultid="3151" />
                    <RANKING order="4" place="4" resultid="5503" />
                    <RANKING order="5" place="5" resultid="5371" />
                    <RANKING order="6" place="6" resultid="3578" />
                    <RANKING order="7" place="7" resultid="2954" />
                    <RANKING order="8" place="8" resultid="3448" />
                    <RANKING order="9" place="9" resultid="4575" />
                    <RANKING order="10" place="10" resultid="3563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3848" />
                    <RANKING order="2" place="2" resultid="3665" />
                    <RANKING order="3" place="3" resultid="3671" />
                    <RANKING order="4" place="4" resultid="3675" />
                    <RANKING order="5" place="5" resultid="4284" />
                    <RANKING order="6" place="6" resultid="4418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4602" />
                    <RANKING order="2" place="2" resultid="2967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4015" />
                    <RANKING order="2" place="2" resultid="4608" />
                    <RANKING order="3" place="3" resultid="5067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4055" />
                    <RANKING order="2" place="2" resultid="3259" />
                    <RANKING order="3" place="3" resultid="5168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4901" />
                    <RANKING order="2" place="2" resultid="4236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5184" />
                    <RANKING order="2" place="2" resultid="3454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="1073" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="1074" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="1075" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5766" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5767" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5768" daytime="09:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5769" daytime="09:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5770" daytime="09:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5771" daytime="09:08" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:10" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6054" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5651" />
                    <RANKING order="2" place="2" resultid="4882" />
                    <RANKING order="3" place="3" resultid="4823" />
                    <RANKING order="4" place="4" resultid="4366" />
                    <RANKING order="5" place="5" resultid="3639" />
                    <RANKING order="6" place="6" resultid="3475" />
                    <RANKING order="7" place="7" resultid="3948" />
                    <RANKING order="8" place="8" resultid="3023" />
                    <RANKING order="9" place="-1" resultid="3218" />
                    <RANKING order="10" place="-1" resultid="4249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6055" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2982" />
                    <RANKING order="2" place="2" resultid="4162" />
                    <RANKING order="3" place="3" resultid="3905" />
                    <RANKING order="4" place="4" resultid="4522" />
                    <RANKING order="5" place="5" resultid="5538" />
                    <RANKING order="6" place="6" resultid="3272" />
                    <RANKING order="7" place="7" resultid="3279" />
                    <RANKING order="8" place="8" resultid="3098" />
                    <RANKING order="9" place="9" resultid="2819" />
                    <RANKING order="10" place="10" resultid="5366" />
                    <RANKING order="11" place="11" resultid="3386" />
                    <RANKING order="12" place="-1" resultid="4131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6056" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4207" />
                    <RANKING order="2" place="2" resultid="5352" />
                    <RANKING order="3" place="3" resultid="3511" />
                    <RANKING order="4" place="4" resultid="4436" />
                    <RANKING order="5" place="5" resultid="2730" />
                    <RANKING order="6" place="6" resultid="4124" />
                    <RANKING order="7" place="7" resultid="3941" />
                    <RANKING order="8" place="8" resultid="3976" />
                    <RANKING order="9" place="8" resultid="5433" />
                    <RANKING order="10" place="10" resultid="3969" />
                    <RANKING order="11" place="-1" resultid="3310" />
                    <RANKING order="12" place="-1" resultid="3990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6057" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4533" />
                    <RANKING order="2" place="2" resultid="4906" />
                    <RANKING order="3" place="3" resultid="4749" />
                    <RANKING order="4" place="4" resultid="5414" />
                    <RANKING order="5" place="5" resultid="5205" />
                    <RANKING order="6" place="6" resultid="4181" />
                    <RANKING order="7" place="7" resultid="4188" />
                    <RANKING order="8" place="8" resultid="3962" />
                    <RANKING order="9" place="9" resultid="3983" />
                    <RANKING order="10" place="10" resultid="3129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6058" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4992" />
                    <RANKING order="2" place="2" resultid="5520" />
                    <RANKING order="3" place="3" resultid="3729" />
                    <RANKING order="4" place="4" resultid="4425" />
                    <RANKING order="5" place="5" resultid="3155" />
                    <RANKING order="6" place="6" resultid="3701" />
                    <RANKING order="7" place="7" resultid="4614" />
                    <RANKING order="8" place="8" resultid="4812" />
                    <RANKING order="9" place="9" resultid="3391" />
                    <RANKING order="10" place="10" resultid="2829" />
                    <RANKING order="11" place="11" resultid="4507" />
                    <RANKING order="12" place="12" resultid="3167" />
                    <RANKING order="13" place="13" resultid="3146" />
                    <RANKING order="14" place="14" resultid="2810" />
                    <RANKING order="15" place="15" resultid="5229" />
                    <RANKING order="16" place="16" resultid="5449" />
                    <RANKING order="17" place="17" resultid="3073" />
                    <RANKING order="18" place="18" resultid="4999" />
                    <RANKING order="19" place="19" resultid="5214" />
                    <RANKING order="20" place="20" resultid="3180" />
                    <RANKING order="21" place="-1" resultid="2756" />
                    <RANKING order="22" place="-1" resultid="2823" />
                    <RANKING order="23" place="-1" resultid="5515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6059" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4169" />
                    <RANKING order="2" place="2" resultid="2851" />
                    <RANKING order="3" place="3" resultid="5526" />
                    <RANKING order="4" place="4" resultid="3544" />
                    <RANKING order="5" place="5" resultid="4817" />
                    <RANKING order="6" place="6" resultid="2878" />
                    <RANKING order="7" place="7" resultid="4527" />
                    <RANKING order="8" place="8" resultid="4290" />
                    <RANKING order="9" place="9" resultid="5096" />
                    <RANKING order="10" place="10" resultid="4175" />
                    <RANKING order="11" place="11" resultid="3558" />
                    <RANKING order="12" place="12" resultid="4519" />
                    <RANKING order="13" place="13" resultid="5551" />
                    <RANKING order="14" place="14" resultid="4200" />
                    <RANKING order="15" place="-1" resultid="4009" />
                    <RANKING order="16" place="-1" resultid="3612" />
                    <RANKING order="17" place="-1" resultid="5005" />
                    <RANKING order="18" place="-1" resultid="5359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6060" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4069" />
                    <RANKING order="2" place="2" resultid="5235" />
                    <RANKING order="3" place="3" resultid="4383" />
                    <RANKING order="4" place="4" resultid="4971" />
                    <RANKING order="5" place="5" resultid="3488" />
                    <RANKING order="6" place="6" resultid="3381" />
                    <RANKING order="7" place="7" resultid="4194" />
                    <RANKING order="8" place="8" resultid="1664" />
                    <RANKING order="9" place="-1" resultid="4628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6061" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4807" />
                    <RANKING order="2" place="2" resultid="4582" />
                    <RANKING order="3" place="3" resultid="4041" />
                    <RANKING order="4" place="4" resultid="4788" />
                    <RANKING order="5" place="5" resultid="5461" />
                    <RANKING order="6" place="6" resultid="3894" />
                    <RANKING order="7" place="7" resultid="4431" />
                    <RANKING order="8" place="8" resultid="4244" />
                    <RANKING order="9" place="9" resultid="5426" />
                    <RANKING order="10" place="10" resultid="2779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6062" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3302" />
                    <RANKING order="2" place="2" resultid="4621" />
                    <RANKING order="3" place="3" resultid="3210" />
                    <RANKING order="4" place="4" resultid="4389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6063" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5729" />
                    <RANKING order="2" place="2" resultid="3236" />
                    <RANKING order="3" place="3" resultid="2764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6064" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5140" />
                    <RANKING order="2" place="2" resultid="5125" />
                    <RANKING order="3" place="3" resultid="4034" />
                    <RANKING order="4" place="4" resultid="1676" />
                    <RANKING order="5" place="-1" resultid="2749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6065" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6066" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6067" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6068" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6069" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5772" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5773" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5774" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5775" daytime="09:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5776" daytime="09:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5777" daytime="09:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5778" daytime="09:18" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5779" daytime="09:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5780" daytime="09:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5781" daytime="09:22" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5782" daytime="09:24" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5783" daytime="09:24" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="09:26" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6070" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4911" />
                    <RANKING order="2" place="2" resultid="5309" />
                    <RANKING order="3" place="3" resultid="5421" />
                    <RANKING order="4" place="4" resultid="2790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6071" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6072" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3366" />
                    <RANKING order="2" place="2" resultid="3839" />
                    <RANKING order="3" place="3" resultid="5325" />
                    <RANKING order="4" place="-1" resultid="5763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6073" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5012" />
                    <RANKING order="2" place="2" resultid="4874" />
                    <RANKING order="3" place="3" resultid="5429" />
                    <RANKING order="4" place="4" resultid="5084" />
                    <RANKING order="5" place="5" resultid="4098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6074" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5504" />
                    <RANKING order="2" place="2" resultid="4779" />
                    <RANKING order="3" place="3" resultid="5372" />
                    <RANKING order="4" place="4" resultid="3523" />
                    <RANKING order="5" place="5" resultid="4640" />
                    <RANKING order="6" place="6" resultid="5089" />
                    <RANKING order="7" place="7" resultid="4632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6075" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5175" />
                    <RANKING order="2" place="2" resultid="4922" />
                    <RANKING order="3" place="3" resultid="4636" />
                    <RANKING order="4" place="4" resultid="2874" />
                    <RANKING order="5" place="5" resultid="4419" />
                    <RANKING order="6" place="6" resultid="4441" />
                    <RANKING order="7" place="-1" resultid="4301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6076" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4256" />
                    <RANKING order="2" place="2" resultid="2858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6077" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6078" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3887" />
                    <RANKING order="2" place="2" resultid="3712" />
                    <RANKING order="3" place="3" resultid="5169" />
                    <RANKING order="4" place="4" resultid="4108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6079" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3232" />
                    <RANKING order="2" place="2" resultid="5400" />
                    <RANKING order="3" place="3" resultid="4853" />
                    <RANKING order="4" place="4" resultid="2913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6080" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5189" />
                    <RANKING order="2" place="2" resultid="4916" />
                    <RANKING order="3" place="3" resultid="2892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6081" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5135" />
                    <RANKING order="2" place="2" resultid="2899" />
                    <RANKING order="3" place="3" resultid="4091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6082" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6083" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6084" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6085" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5784" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5785" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5786" daytime="09:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5787" daytime="09:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5788" daytime="09:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="09:42" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6086" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4374" />
                    <RANKING order="2" place="2" resultid="3955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6087" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4984" />
                    <RANKING order="2" place="2" resultid="4659" />
                    <RANKING order="3" place="3" resultid="4841" />
                    <RANKING order="4" place="4" resultid="3112" />
                    <RANKING order="5" place="5" resultid="2996" />
                    <RANKING order="6" place="6" resultid="5292" />
                    <RANKING order="7" place="7" resultid="4497" />
                    <RANKING order="8" place="8" resultid="4927" />
                    <RANKING order="9" place="9" resultid="5346" />
                    <RANKING order="10" place="-1" resultid="4080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6088" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5019" />
                    <RANKING order="2" place="2" resultid="3567" />
                    <RANKING order="3" place="3" resultid="4125" />
                    <RANKING order="4" place="-1" resultid="4270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6089" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3040" />
                    <RANKING order="2" place="2" resultid="3357" />
                    <RANKING order="3" place="3" resultid="5240" />
                    <RANKING order="4" place="4" resultid="4182" />
                    <RANKING order="5" place="5" resultid="3322" />
                    <RANKING order="6" place="6" resultid="1656" />
                    <RANKING order="7" place="-1" resultid="3984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6090" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4426" />
                    <RANKING order="2" place="2" resultid="3392" />
                    <RANKING order="3" place="3" resultid="4683" />
                    <RANKING order="4" place="4" resultid="2824" />
                    <RANKING order="5" place="5" resultid="4218" />
                    <RANKING order="6" place="6" resultid="4308" />
                    <RANKING order="7" place="7" resultid="4838" />
                    <RANKING order="8" place="8" resultid="3185" />
                    <RANKING order="9" place="9" resultid="4677" />
                    <RANKING order="10" place="10" resultid="5103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6091" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3545" />
                    <RANKING order="2" place="2" resultid="4022" />
                    <RANKING order="3" place="3" resultid="3690" />
                    <RANKING order="4" place="4" resultid="4760" />
                    <RANKING order="5" place="5" resultid="3289" />
                    <RANKING order="6" place="6" resultid="4653" />
                    <RANKING order="7" place="7" resultid="4314" />
                    <RANKING order="8" place="-1" resultid="3268" />
                    <RANKING order="9" place="-1" resultid="4672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6092" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3551" />
                    <RANKING order="2" place="2" resultid="3503" />
                    <RANKING order="3" place="3" resultid="3285" />
                    <RANKING order="4" place="4" resultid="2927" />
                    <RANKING order="5" place="5" resultid="4195" />
                    <RANKING order="6" place="6" resultid="4263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6093" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5280" />
                    <RANKING order="2" place="2" resultid="5030" />
                    <RANKING order="3" place="3" resultid="5024" />
                    <RANKING order="4" place="4" resultid="4934" />
                    <RANKING order="5" place="5" resultid="4445" />
                    <RANKING order="6" place="6" resultid="4048" />
                    <RANKING order="7" place="-1" resultid="3617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6094" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5314" />
                    <RANKING order="2" place="2" resultid="5261" />
                    <RANKING order="3" place="3" resultid="4212" />
                    <RANKING order="4" place="4" resultid="3211" />
                    <RANKING order="5" place="5" resultid="4028" />
                    <RANKING order="6" place="6" resultid="4666" />
                    <RANKING order="7" place="7" resultid="4399" />
                    <RANKING order="8" place="8" resultid="4662" />
                    <RANKING order="9" place="9" resultid="2933" />
                    <RANKING order="10" place="10" resultid="3515" />
                    <RANKING order="11" place="-1" resultid="4404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6095" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3404" />
                    <RANKING order="2" place="2" resultid="4589" />
                    <RANKING order="3" place="3" resultid="5568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6096" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4646" />
                    <RANKING order="2" place="2" resultid="2920" />
                    <RANKING order="3" place="3" resultid="3015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6097" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3338" />
                    <RANKING order="2" place="2" resultid="3481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6098" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5130" />
                    <RANKING order="2" place="2" resultid="3460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6099" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6100" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3496" />
                    <RANKING order="2" place="2" resultid="2771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6101" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5789" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5790" daytime="09:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5791" daytime="09:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5792" daytime="09:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5793" daytime="09:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5794" daytime="09:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5795" daytime="09:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5796" daytime="10:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="10:02" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6102" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4938" />
                    <RANKING order="2" place="2" resultid="2815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6103" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3879" />
                    <RANKING order="2" place="2" resultid="3854" />
                    <RANKING order="3" place="3" resultid="3346" />
                    <RANKING order="4" place="4" resultid="4897" />
                    <RANKING order="5" place="5" resultid="4344" />
                    <RANKING order="6" place="6" resultid="3119" />
                    <RANKING order="7" place="-1" resultid="4747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6104" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3421" />
                    <RANKING order="2" place="2" resultid="4803" />
                    <RANKING order="3" place="3" resultid="5247" />
                    <RANKING order="4" place="4" resultid="3574" />
                    <RANKING order="5" place="5" resultid="3681" />
                    <RANKING order="6" place="6" resultid="3226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6105" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5013" />
                    <RANKING order="2" place="2" resultid="5297" />
                    <RANKING order="3" place="3" resultid="4875" />
                    <RANKING order="4" place="4" resultid="4103" />
                    <RANKING order="5" place="5" resultid="3659" />
                    <RANKING order="6" place="6" resultid="3174" />
                    <RANKING order="7" place="7" resultid="4099" />
                    <RANKING order="8" place="-1" resultid="3644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6106" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4570" />
                    <RANKING order="2" place="2" resultid="3898" />
                    <RANKING order="3" place="3" resultid="4738" />
                    <RANKING order="4" place="4" resultid="2948" />
                    <RANKING order="5" place="5" resultid="5318" />
                    <RANKING order="6" place="6" resultid="3579" />
                    <RANKING order="7" place="7" resultid="2955" />
                    <RANKING order="8" place="8" resultid="4641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6107" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4690" />
                    <RANKING order="2" place="2" resultid="4764" />
                    <RANKING order="3" place="3" resultid="4062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6108" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6109" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4016" />
                    <RANKING order="2" place="2" resultid="4609" />
                    <RANKING order="3" place="3" resultid="4859" />
                    <RANKING order="4" place="4" resultid="2959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6110" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5161" />
                    <RANKING order="2" place="2" resultid="3260" />
                    <RANKING order="3" place="3" resultid="4319" />
                    <RANKING order="4" place="4" resultid="3888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6111" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4902" />
                    <RANKING order="2" place="2" resultid="4237" />
                    <RANKING order="3" place="3" resultid="2906" />
                    <RANKING order="4" place="4" resultid="2914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6112" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5185" />
                    <RANKING order="2" place="2" resultid="3455" />
                    <RANKING order="3" place="3" resultid="5151" />
                    <RANKING order="4" place="4" resultid="5190" />
                    <RANKING order="5" place="5" resultid="2893" />
                    <RANKING order="6" place="6" resultid="4917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6113" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2900" />
                    <RANKING order="2" place="2" resultid="4092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6114" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6115" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6116" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6117" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5797" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5798" daytime="10:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5799" daytime="10:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5800" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5801" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5802" daytime="10:12" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="10:14" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6118" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4883" />
                    <RANKING order="2" place="2" resultid="3441" />
                    <RANKING order="3" place="3" resultid="5652" />
                    <RANKING order="4" place="4" resultid="3949" />
                    <RANKING order="5" place="5" resultid="2737" />
                    <RANKING order="6" place="6" resultid="3476" />
                    <RANKING order="7" place="7" resultid="3219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6119" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5531" />
                    <RANKING order="2" place="2" resultid="3906" />
                    <RANKING order="3" place="3" resultid="3273" />
                    <RANKING order="4" place="-1" resultid="5722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6120" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5120" />
                    <RANKING order="2" place="2" resultid="2972" />
                    <RANKING order="3" place="3" resultid="3942" />
                    <RANKING order="4" place="4" resultid="4075" />
                    <RANKING order="5" place="5" resultid="4772" />
                    <RANKING order="6" place="6" resultid="3977" />
                    <RANKING order="7" place="7" resultid="3318" />
                    <RANKING order="8" place="8" resultid="3970" />
                    <RANKING order="9" place="-1" resultid="3991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6121" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3398" />
                    <RANKING order="2" place="2" resultid="2978" />
                    <RANKING order="3" place="3" resultid="3686" />
                    <RANKING order="4" place="4" resultid="5209" />
                    <RANKING order="5" place="-1" resultid="3314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6122" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4993" />
                    <RANKING order="2" place="2" resultid="3730" />
                    <RANKING order="3" place="3" resultid="3156" />
                    <RANKING order="4" place="4" resultid="4469" />
                    <RANKING order="5" place="5" resultid="4615" />
                    <RANKING order="6" place="6" resultid="3047" />
                    <RANKING order="7" place="7" resultid="4223" />
                    <RANKING order="8" place="8" resultid="5043" />
                    <RANKING order="9" place="9" resultid="2811" />
                    <RANKING order="10" place="10" resultid="4678" />
                    <RANKING order="11" place="11" resultid="5225" />
                    <RANKING order="12" place="12" resultid="5450" />
                    <RANKING order="13" place="13" resultid="3147" />
                    <RANKING order="14" place="14" resultid="4978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6123" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4528" />
                    <RANKING order="2" place="2" resultid="5527" />
                    <RANKING order="3" place="3" resultid="4450" />
                    <RANKING order="4" place="4" resultid="4326" />
                    <RANKING order="5" place="5" resultid="5097" />
                    <RANKING order="6" place="6" resultid="4330" />
                    <RANKING order="7" place="7" resultid="3537" />
                    <RANKING order="8" place="8" resultid="4846" />
                    <RANKING order="9" place="9" resultid="5386" />
                    <RANKING order="10" place="10" resultid="4201" />
                    <RANKING order="11" place="-1" resultid="3613" />
                    <RANKING order="12" place="-1" resultid="4768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6124" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3627" />
                    <RANKING order="2" place="2" resultid="2928" />
                    <RANKING order="3" place="3" resultid="3011" />
                    <RANKING order="4" place="4" resultid="4948" />
                    <RANKING order="5" place="5" resultid="3695" />
                    <RANKING order="6" place="6" resultid="4547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6125" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4808" />
                    <RANKING order="2" place="2" resultid="3376" />
                    <RANKING order="3" place="3" resultid="4457" />
                    <RANKING order="4" place="4" resultid="4042" />
                    <RANKING order="5" place="5" resultid="4789" />
                    <RANKING order="6" place="6" resultid="5462" />
                    <RANKING order="7" place="7" resultid="2844" />
                    <RANKING order="8" place="8" resultid="3090" />
                    <RANKING order="9" place="9" resultid="5457" />
                    <RANKING order="10" place="10" resultid="3134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6126" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                    <RANKING order="2" place="2" resultid="4351" />
                    <RANKING order="3" place="3" resultid="4869" />
                    <RANKING order="4" place="4" resultid="5218" />
                    <RANKING order="5" place="5" resultid="5036" />
                    <RANKING order="6" place="6" resultid="4410" />
                    <RANKING order="7" place="7" resultid="4667" />
                    <RANKING order="8" place="8" resultid="4405" />
                    <RANKING order="9" place="-1" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6127" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5730" />
                    <RANKING order="2" place="2" resultid="5144" />
                    <RANKING order="3" place="3" resultid="4942" />
                    <RANKING order="4" place="4" resultid="4511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6128" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4552" />
                    <RANKING order="2" place="2" resultid="4647" />
                    <RANKING order="3" place="3" resultid="5126" />
                    <RANKING order="4" place="4" resultid="2940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6129" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6130" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3461" />
                    <RANKING order="2" place="2" resultid="3061" />
                    <RANKING order="3" place="3" resultid="5743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6131" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6132" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6133" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5803" daytime="10:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5804" daytime="10:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5805" daytime="10:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5806" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5807" daytime="10:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5808" daytime="10:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5809" daytime="10:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5810" daytime="10:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5811" daytime="10:28" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1161" daytime="10:30" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6134" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2990" />
                    <RANKING order="2" place="2" resultid="5422" />
                    <RANKING order="3" place="3" resultid="5310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6135" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4360" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="3429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6136" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3351" />
                    <RANKING order="2" place="2" resultid="5341" />
                    <RANKING order="3" place="3" resultid="5509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6137" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3929" />
                    <RANKING order="2" place="2" resultid="5757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6138" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3899" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="3160" />
                    <RANKING order="4" place="4" resultid="5758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6139" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4923" />
                    <RANKING order="2" place="2" resultid="4285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6140" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4603" />
                    <RANKING order="2" place="2" resultid="2859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6141" agemax="59" agemin="55" name="Kategoria G" />
                <AGEGROUP agegroupid="6142" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4320" />
                    <RANKING order="2" place="2" resultid="4109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6143" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="6144" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="6145" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6146" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6147" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6148" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6149" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5812" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5813" daytime="10:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5814" daytime="10:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1178" daytime="10:42" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6150" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                    <RANKING order="2" place="2" resultid="3294" />
                    <RANKING order="3" place="3" resultid="3203" />
                    <RANKING order="4" place="4" resultid="3956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6151" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4163" />
                    <RANKING order="2" place="2" resultid="2997" />
                    <RANKING order="3" place="3" resultid="3099" />
                    <RANKING order="4" place="4" resultid="3280" />
                    <RANKING order="5" place="-1" resultid="4474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6152" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5353" />
                    <RANKING order="2" place="2" resultid="3568" />
                    <RANKING order="3" place="3" resultid="5434" />
                    <RANKING order="4" place="4" resultid="3844" />
                    <RANKING order="5" place="5" resultid="3240" />
                    <RANKING order="6" place="6" resultid="5393" />
                    <RANKING order="7" place="-1" resultid="5064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6153" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="5720" />
                    <RANKING order="3" place="3" resultid="3963" />
                    <RANKING order="4" place="4" resultid="3871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6154" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2802" />
                    <RANKING order="2" place="2" resultid="3048" />
                    <RANKING order="3" place="3" resultid="4684" />
                    <RANKING order="4" place="4" resultid="5044" />
                    <RANKING order="5" place="5" resultid="3186" />
                    <RANKING order="6" place="6" resultid="3181" />
                    <RANKING order="7" place="-1" resultid="2757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6155" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2852" />
                    <RANKING order="2" place="2" resultid="4889" />
                    <RANKING order="3" place="3" resultid="4023" />
                    <RANKING order="4" place="4" resultid="4291" />
                    <RANKING order="5" place="5" resultid="3559" />
                    <RANKING order="6" place="-1" resultid="5006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6156" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="5254" />
                    <RANKING order="3" place="3" resultid="5236" />
                    <RANKING order="4" place="4" resultid="2882" />
                    <RANKING order="5" place="5" resultid="4972" />
                    <RANKING order="6" place="6" resultid="1665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6157" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3377" />
                    <RANKING order="2" place="2" resultid="5281" />
                    <RANKING order="3" place="3" resultid="4583" />
                    <RANKING order="4" place="4" resultid="2866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6158" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4352" />
                    <RANKING order="2" place="2" resultid="2785" />
                    <RANKING order="3" place="3" resultid="4213" />
                    <RANKING order="4" place="4" resultid="4694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6159" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3405" />
                    <RANKING order="2" place="2" resultid="4943" />
                    <RANKING order="3" place="3" resultid="4698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6160" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5750" />
                    <RANKING order="2" place="2" resultid="3054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6161" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6162" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6163" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6164" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6165" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5815" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5816" daytime="10:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5817" daytime="10:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5818" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5819" daytime="11:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5820" daytime="11:06" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="11:10" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6166" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3648" />
                    <RANKING order="2" place="2" resultid="3437" />
                    <RANKING order="3" place="3" resultid="5764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6167" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5081" />
                    <RANKING order="2" place="2" resultid="4556" />
                    <RANKING order="3" place="3" resultid="2796" />
                    <RANKING order="4" place="4" resultid="3004" />
                    <RANKING order="5" place="5" resultid="3120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6168" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5074" />
                    <RANKING order="2" place="2" resultid="3531" />
                    <RANKING order="3" place="3" resultid="5248" />
                    <RANKING order="4" place="4" resultid="4335" />
                    <RANKING order="5" place="5" resultid="5342" />
                    <RANKING order="6" place="6" resultid="3227" />
                    <RANKING order="7" place="7" resultid="3840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6169" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3930" />
                    <RANKING order="2" place="2" resultid="4705" />
                    <RANKING order="3" place="3" resultid="3126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6170" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3142" />
                    <RANKING order="2" place="2" resultid="5319" />
                    <RANKING order="3" place="3" resultid="2949" />
                    <RANKING order="4" place="4" resultid="3161" />
                    <RANKING order="5" place="5" resultid="4576" />
                    <RANKING order="6" place="6" resultid="5090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6171" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5176" />
                    <RANKING order="2" place="2" resultid="3849" />
                    <RANKING order="3" place="3" resultid="4302" />
                    <RANKING order="4" place="4" resultid="3666" />
                    <RANKING order="5" place="5" resultid="4063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6172" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6173" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3244" />
                    <RANKING order="2" place="2" resultid="4480" />
                    <RANKING order="3" place="3" resultid="5069" />
                    <RANKING order="4" place="-1" resultid="2960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6174" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4056" />
                    <RANKING order="2" place="2" resultid="5162" />
                    <RANKING order="3" place="3" resultid="4593" />
                    <RANKING order="4" place="4" resultid="3859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6175" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3067" />
                    <RANKING order="2" place="2" resultid="2907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6176" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6177" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6178" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6179" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6180" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6181" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5821" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5822" daytime="11:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5823" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5824" daytime="11:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5825" daytime="11:28" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="11:32" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6182" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3295" />
                    <RANKING order="2" place="2" resultid="4378" />
                    <RANKING order="3" place="3" resultid="4367" />
                    <RANKING order="4" place="4" resultid="4824" />
                    <RANKING order="5" place="-1" resultid="2738" />
                    <RANKING order="6" place="-1" resultid="4250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6183" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5532" />
                    <RANKING order="2" place="2" resultid="2983" />
                    <RANKING order="3" place="3" resultid="4561" />
                    <RANKING order="4" place="4" resultid="4928" />
                    <RANKING order="5" place="5" resultid="5367" />
                    <RANKING order="6" place="6" resultid="5380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6184" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5721" />
                    <RANKING order="2" place="2" resultid="3264" />
                    <RANKING order="3" place="3" resultid="5394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6185" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5050" />
                    <RANKING order="2" place="2" resultid="4534" />
                    <RANKING order="3" place="3" resultid="3041" />
                    <RANKING order="4" place="4" resultid="3399" />
                    <RANKING order="5" place="5" resultid="4189" />
                    <RANKING order="6" place="6" resultid="3029" />
                    <RANKING order="7" place="7" resultid="4276" />
                    <RANKING order="8" place="8" resultid="3872" />
                    <RANKING order="9" place="9" resultid="1657" />
                    <RANKING order="10" place="-1" resultid="4907" />
                    <RANKING order="11" place="-1" resultid="4955" />
                    <RANKING order="12" place="-1" resultid="5466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6186" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2803" />
                    <RANKING order="2" place="2" resultid="4224" />
                    <RANKING order="3" place="3" resultid="4486" />
                    <RANKING order="4" place="4" resultid="5451" />
                    <RANKING order="5" place="5" resultid="4979" />
                    <RANKING order="6" place="6" resultid="5000" />
                    <RANKING order="7" place="7" resultid="3074" />
                    <RANKING order="8" place="8" resultid="5560" />
                    <RANKING order="9" place="9" resultid="5104" />
                    <RANKING order="10" place="-1" resultid="4309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6187" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4170" />
                    <RANKING order="2" place="2" resultid="4795" />
                    <RANKING order="3" place="3" resultid="4451" />
                    <RANKING order="4" place="4" resultid="5442" />
                    <RANKING order="5" place="5" resultid="4176" />
                    <RANKING order="6" place="6" resultid="3538" />
                    <RANKING order="7" place="7" resultid="4847" />
                    <RANKING order="8" place="8" resultid="4654" />
                    <RANKING order="9" place="9" resultid="5387" />
                    <RANKING order="10" place="-1" resultid="3653" />
                    <RANKING order="11" place="-1" resultid="3691" />
                    <RANKING order="12" place="-1" resultid="4331" />
                    <RANKING order="13" place="-1" resultid="5114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6188" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5255" />
                    <RANKING order="2" place="2" resultid="3504" />
                    <RANKING order="3" place="3" resultid="3628" />
                    <RANKING order="4" place="4" resultid="3489" />
                    <RANKING order="5" place="5" resultid="4949" />
                    <RANKING order="6" place="6" resultid="3696" />
                    <RANKING order="7" place="7" resultid="3382" />
                    <RANKING order="8" place="8" resultid="4264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6189" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2725" />
                    <RANKING order="2" place="2" resultid="4458" />
                    <RANKING order="3" place="3" resultid="5025" />
                    <RANKING order="4" place="4" resultid="4049" />
                    <RANKING order="5" place="5" resultid="2845" />
                    <RANKING order="6" place="6" resultid="3091" />
                    <RANKING order="7" place="7" resultid="4432" />
                    <RANKING order="8" place="8" resultid="2867" />
                    <RANKING order="9" place="9" resultid="3135" />
                    <RANKING order="10" place="10" resultid="2780" />
                    <RANKING order="11" place="-1" resultid="3618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6190" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4622" />
                    <RANKING order="2" place="2" resultid="4715" />
                    <RANKING order="3" place="3" resultid="5037" />
                    <RANKING order="4" place="4" resultid="4390" />
                    <RANKING order="5" place="5" resultid="3361" />
                    <RANKING order="6" place="6" resultid="2934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6191" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5145" />
                    <RANKING order="2" place="2" resultid="3035" />
                    <RANKING order="3" place="3" resultid="4512" />
                    <RANKING order="4" place="4" resultid="2765" />
                    <RANKING order="5" place="5" resultid="4699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6192" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4710" />
                    <RANKING order="2" place="2" resultid="4035" />
                    <RANKING order="3" place="3" resultid="2750" />
                    <RANKING order="4" place="4" resultid="2921" />
                    <RANKING order="5" place="5" resultid="5751" />
                    <RANKING order="6" place="6" resultid="2941" />
                    <RANKING order="7" place="7" resultid="1677" />
                    <RANKING order="8" place="8" resultid="3016" />
                    <RANKING order="9" place="-1" resultid="3055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6193" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4463" />
                    <RANKING order="2" place="2" resultid="3482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6194" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5156" />
                    <RANKING order="2" place="2" resultid="4085" />
                    <RANKING order="3" place="3" resultid="5744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6195" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6196" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6197" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5826" daytime="11:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5827" daytime="11:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5828" daytime="11:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5829" daytime="11:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5830" daytime="11:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5831" daytime="11:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5832" daytime="12:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5833" daytime="12:04" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5834" daytime="12:06" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5835" daytime="12:10" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1229" daytime="12:14" gender="X" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1230" agemax="-1" agemin="-1" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="1231" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL" />
                <AGEGROUP agegroupid="1232" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3734" />
                    <RANKING order="2" place="2" resultid="3911" />
                    <RANKING order="3" place="3" resultid="3735" />
                    <RANKING order="4" place="-1" resultid="3584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4728" />
                    <RANKING order="2" place="2" resultid="3191" />
                    <RANKING order="3" place="3" resultid="3716" />
                    <RANKING order="4" place="4" resultid="3585" />
                    <RANKING order="5" place="5" resultid="5330" />
                    <RANKING order="6" place="6" resultid="3910" />
                    <RANKING order="7" place="7" resultid="4489" />
                    <RANKING order="8" place="-1" resultid="3717" />
                    <RANKING order="9" place="-1" resultid="5566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="5329" />
                    <RANKING order="3" place="3" resultid="3909" />
                    <RANKING order="4" place="4" resultid="3718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4118" />
                    <RANKING order="2" place="2" resultid="4727" />
                    <RANKING order="3" place="3" resultid="4962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="-1" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5194" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5836" daytime="12:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5837" daytime="12:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5838" daytime="12:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-12-11" daytime="15:10" endtime="18:45" number="2">
          <EVENTS>
            <EVENT eventid="1247" daytime="15:10" gender="F" number="12" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6198" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2991" />
                    <RANKING order="2" place="2" resultid="3649" />
                    <RANKING order="3" place="3" resultid="3433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6199" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="2797" />
                    <RANKING order="3" place="3" resultid="4361" />
                    <RANKING order="4" place="4" resultid="3880" />
                    <RANKING order="5" place="5" resultid="3121" />
                    <RANKING order="6" place="6" resultid="4557" />
                    <RANKING order="7" place="7" resultid="3005" />
                    <RANKING order="8" place="8" resultid="5078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6200" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4804" />
                    <RANKING order="2" place="2" resultid="5073" />
                    <RANKING order="3" place="3" resultid="3532" />
                    <RANKING order="4" place="4" resultid="4336" />
                    <RANKING order="5" place="5" resultid="5249" />
                    <RANKING order="6" place="6" resultid="5343" />
                    <RANKING order="7" place="-1" resultid="5640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6201" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3175" />
                    <RANKING order="2" place="2" resultid="3127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6202" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4739" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="2950" />
                    <RANKING order="4" place="4" resultid="3580" />
                    <RANKING order="5" place="5" resultid="2956" />
                    <RANKING order="6" place="6" resultid="5320" />
                    <RANKING order="7" place="7" resultid="5091" />
                    <RANKING order="8" place="8" resultid="4633" />
                    <RANKING order="9" place="-1" resultid="4780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6203" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5177" />
                    <RANKING order="2" place="2" resultid="4303" />
                    <RANKING order="3" place="3" resultid="3667" />
                    <RANKING order="4" place="4" resultid="3672" />
                    <RANKING order="5" place="5" resultid="4064" />
                    <RANKING order="6" place="6" resultid="4420" />
                    <RANKING order="7" place="7" resultid="3868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6204" agemax="54" agemin="50" name="Kategoria F" />
                <AGEGROUP agegroupid="6205" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3245" />
                    <RANKING order="2" place="2" resultid="4860" />
                    <RANKING order="3" place="3" resultid="4481" />
                    <RANKING order="4" place="4" resultid="5068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6206" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4057" />
                    <RANKING order="2" place="2" resultid="4594" />
                    <RANKING order="3" place="3" resultid="3860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6207" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4238" />
                    <RANKING order="2" place="2" resultid="2908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6208" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5152" />
                    <RANKING order="2" place="2" resultid="3373" />
                    <RANKING order="3" place="3" resultid="2894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6209" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2901" />
                    <RANKING order="2" place="2" resultid="4093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6210" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6211" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6212" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6213" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5839" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5840" daytime="15:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5841" daytime="15:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5842" daytime="15:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5843" daytime="15:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5844" daytime="15:24" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1265" daytime="15:26" gender="M" number="13" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6214" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4368" />
                    <RANKING order="2" place="2" resultid="4825" />
                    <RANKING order="3" place="3" resultid="4379" />
                    <RANKING order="4" place="4" resultid="3641" />
                    <RANKING order="5" place="5" resultid="2739" />
                    <RANKING order="6" place="6" resultid="3950" />
                    <RANKING order="7" place="7" resultid="3024" />
                    <RANKING order="8" place="8" resultid="3204" />
                    <RANKING order="9" place="-1" resultid="4251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6215" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4523" />
                    <RANKING order="2" place="2" resultid="3907" />
                    <RANKING order="3" place="3" resultid="5539" />
                    <RANKING order="4" place="4" resultid="5663" />
                    <RANKING order="5" place="5" resultid="2984" />
                    <RANKING order="6" place="6" resultid="4132" />
                    <RANKING order="7" place="7" resultid="4565" />
                    <RANKING order="8" place="8" resultid="4562" />
                    <RANKING order="9" place="9" resultid="4929" />
                    <RANKING order="10" place="10" resultid="2820" />
                    <RANKING order="11" place="11" resultid="5347" />
                    <RANKING order="12" place="12" resultid="4081" />
                    <RANKING order="13" place="13" resultid="5381" />
                    <RANKING order="14" place="14" resultid="3387" />
                    <RANKING order="15" place="-1" resultid="4475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6216" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4208" />
                    <RANKING order="2" place="2" resultid="4437" />
                    <RANKING order="3" place="3" resultid="4501" />
                    <RANKING order="4" place="4" resultid="2973" />
                    <RANKING order="5" place="5" resultid="5435" />
                    <RANKING order="6" place="6" resultid="2731" />
                    <RANKING order="7" place="7" resultid="3943" />
                    <RANKING order="8" place="8" resultid="4135" />
                    <RANKING order="9" place="9" resultid="3978" />
                    <RANKING order="10" place="10" resultid="3109" />
                    <RANKING order="11" place="11" resultid="3992" />
                    <RANKING order="12" place="12" resultid="3971" />
                    <RANKING order="13" place="13" resultid="3319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6217" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5051" />
                    <RANKING order="2" place="2" resultid="4535" />
                    <RANKING order="3" place="3" resultid="4784" />
                    <RANKING order="4" place="4" resultid="3400" />
                    <RANKING order="5" place="5" resultid="4908" />
                    <RANKING order="6" place="6" resultid="5206" />
                    <RANKING order="7" place="7" resultid="4190" />
                    <RANKING order="8" place="8" resultid="5242" />
                    <RANKING order="9" place="9" resultid="5210" />
                    <RANKING order="10" place="10" resultid="2979" />
                    <RANKING order="11" place="11" resultid="3873" />
                    <RANKING order="12" place="12" resultid="4277" />
                    <RANKING order="13" place="13" resultid="3924" />
                    <RANKING order="14" place="14" resultid="3130" />
                    <RANKING order="15" place="-1" resultid="5467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6218" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4994" />
                    <RANKING order="2" place="2" resultid="2804" />
                    <RANKING order="3" place="3" resultid="4508" />
                    <RANKING order="4" place="4" resultid="4225" />
                    <RANKING order="5" place="5" resultid="2830" />
                    <RANKING order="6" place="6" resultid="3168" />
                    <RANKING order="7" place="7" resultid="3393" />
                    <RANKING order="8" place="8" resultid="5215" />
                    <RANKING order="9" place="9" resultid="5001" />
                    <RANKING order="10" place="10" resultid="4679" />
                    <RANKING order="11" place="11" resultid="3920" />
                    <RANKING order="12" place="12" resultid="5561" />
                    <RANKING order="13" place="13" resultid="5105" />
                    <RANKING order="14" place="-1" resultid="3075" />
                    <RANKING order="15" place="-1" resultid="5230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6219" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2853" />
                    <RANKING order="2" place="2" resultid="3546" />
                    <RANKING order="3" place="3" resultid="4796" />
                    <RANKING order="4" place="4" resultid="2879" />
                    <RANKING order="5" place="5" resultid="4452" />
                    <RANKING order="6" place="6" resultid="4332" />
                    <RANKING order="7" place="7" resultid="4818" />
                    <RANKING order="8" place="8" resultid="5443" />
                    <RANKING order="9" place="9" resultid="4177" />
                    <RANKING order="10" place="10" resultid="5098" />
                    <RANKING order="11" place="11" resultid="5552" />
                    <RANKING order="12" place="12" resultid="4202" />
                    <RANKING order="13" place="13" resultid="4010" />
                    <RANKING order="14" place="14" resultid="5388" />
                    <RANKING order="15" place="15" resultid="3864" />
                    <RANKING order="16" place="-1" resultid="3654" />
                    <RANKING order="17" place="-1" resultid="4024" />
                    <RANKING order="18" place="-1" resultid="4673" />
                    <RANKING order="19" place="-1" resultid="5115" />
                    <RANKING order="20" place="-1" resultid="5360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6220" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5256" />
                    <RANKING order="2" place="2" resultid="3505" />
                    <RANKING order="3" place="3" resultid="3629" />
                    <RANKING order="4" place="4" resultid="3490" />
                    <RANKING order="5" place="5" resultid="4950" />
                    <RANKING order="6" place="6" resultid="3697" />
                    <RANKING order="7" place="7" resultid="4196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6221" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2726" />
                    <RANKING order="2" place="2" resultid="3378" />
                    <RANKING order="3" place="3" resultid="4809" />
                    <RANKING order="4" place="4" resultid="4584" />
                    <RANKING order="5" place="5" resultid="4790" />
                    <RANKING order="6" place="6" resultid="4050" />
                    <RANKING order="7" place="7" resultid="2846" />
                    <RANKING order="8" place="8" resultid="5458" />
                    <RANKING order="9" place="9" resultid="5267" />
                    <RANKING order="10" place="10" resultid="2868" />
                    <RANKING order="11" place="11" resultid="3136" />
                    <RANKING order="12" place="-1" resultid="3619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6222" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4623" />
                    <RANKING order="2" place="2" resultid="4716" />
                    <RANKING order="3" place="3" resultid="5038" />
                    <RANKING order="4" place="4" resultid="3362" />
                    <RANKING order="5" place="5" resultid="2935" />
                    <RANKING order="6" place="6" resultid="3705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6223" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4960" />
                    <RANKING order="2" place="2" resultid="3036" />
                    <RANKING order="3" place="3" resultid="5146" />
                    <RANKING order="4" place="4" resultid="4513" />
                    <RANKING order="5" place="5" resultid="2766" />
                    <RANKING order="6" place="6" resultid="4700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6224" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4036" />
                    <RANKING order="2" place="2" resultid="2751" />
                    <RANKING order="3" place="3" resultid="2922" />
                    <RANKING order="4" place="4" resultid="4553" />
                    <RANKING order="5" place="5" resultid="2942" />
                    <RANKING order="6" place="6" resultid="1678" />
                    <RANKING order="7" place="-1" resultid="3017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6225" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6226" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5157" />
                    <RANKING order="2" place="2" resultid="4086" />
                    <RANKING order="3" place="3" resultid="5745" />
                    <RANKING order="4" place="-1" resultid="3062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6227" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6228" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3498" />
                    <RANKING order="2" place="2" resultid="2773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6229" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5845" daytime="15:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5846" daytime="15:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5847" daytime="15:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5848" daytime="15:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5849" daytime="15:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5850" daytime="15:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5851" daytime="15:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5852" daytime="15:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5853" daytime="15:46" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5854" daytime="15:48" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5855" daytime="15:48" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5856" daytime="15:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5857" daytime="15:52" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5858" daytime="15:54" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1282" daytime="15:56" gender="F" number="14" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6230" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5311" />
                    <RANKING order="2" place="2" resultid="4912" />
                    <RANKING order="3" place="3" resultid="4829" />
                    <RANKING order="4" place="4" resultid="2791" />
                    <RANKING order="5" place="5" resultid="5438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6231" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6232" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3367" />
                    <RANKING order="2" place="2" resultid="3352" />
                    <RANKING order="3" place="3" resultid="3841" />
                    <RANKING order="4" place="4" resultid="5326" />
                    <RANKING order="5" place="-1" resultid="5761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6233" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4876" />
                    <RANKING order="2" place="2" resultid="5014" />
                    <RANKING order="3" place="3" resultid="5430" />
                    <RANKING order="4" place="4" resultid="4706" />
                    <RANKING order="5" place="5" resultid="4100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6234" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5505" />
                    <RANKING order="2" place="2" resultid="4781" />
                    <RANKING order="3" place="3" resultid="5373" />
                    <RANKING order="4" place="4" resultid="3525" />
                    <RANKING order="5" place="5" resultid="4642" />
                    <RANKING order="6" place="6" resultid="4577" />
                    <RANKING order="7" place="7" resultid="5092" />
                    <RANKING order="8" place="8" resultid="4634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6235" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5178" />
                    <RANKING order="2" place="2" resultid="4304" />
                    <RANKING order="3" place="3" resultid="4421" />
                    <RANKING order="4" place="4" resultid="5377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6236" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4604" />
                    <RANKING order="2" place="2" resultid="4258" />
                    <RANKING order="3" place="3" resultid="2860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6237" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4017" />
                    <RANKING order="2" place="2" resultid="4861" />
                    <RANKING order="3" place="3" resultid="2961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6238" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3889" />
                    <RANKING order="2" place="2" resultid="3713" />
                    <RANKING order="3" place="3" resultid="5163" />
                    <RANKING order="4" place="4" resultid="3861" />
                    <RANKING order="5" place="5" resultid="5170" />
                    <RANKING order="6" place="6" resultid="4110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6239" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3233" />
                    <RANKING order="2" place="2" resultid="3068" />
                    <RANKING order="3" place="3" resultid="4854" />
                    <RANKING order="4" place="-1" resultid="5401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6240" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5191" />
                    <RANKING order="2" place="2" resultid="2895" />
                    <RANKING order="3" place="-1" resultid="4918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6241" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5136" />
                    <RANKING order="2" place="2" resultid="4094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6242" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6243" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6244" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6245" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5859" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5860" daytime="15:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5861" daytime="16:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5862" daytime="16:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5863" daytime="16:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5864" daytime="16:06" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1299" daytime="16:08" gender="M" number="15" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6246" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4375" />
                    <RANKING order="2" place="2" resultid="5304" />
                    <RANKING order="3" place="3" resultid="3957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6247" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4842" />
                    <RANKING order="2" place="2" resultid="4542" />
                    <RANKING order="3" place="3" resultid="4985" />
                    <RANKING order="4" place="4" resultid="4660" />
                    <RANKING order="5" place="5" resultid="3113" />
                    <RANKING order="6" place="6" resultid="2998" />
                    <RANKING order="7" place="7" resultid="5293" />
                    <RANKING order="8" place="8" resultid="4498" />
                    <RANKING order="9" place="9" resultid="3100" />
                    <RANKING order="10" place="10" resultid="5348" />
                    <RANKING order="11" place="11" resultid="4082" />
                    <RANKING order="12" place="12" resultid="3274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6248" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5020" />
                    <RANKING order="2" place="2" resultid="3569" />
                    <RANKING order="3" place="3" resultid="4126" />
                    <RANKING order="4" place="4" resultid="4076" />
                    <RANKING order="5" place="5" resultid="3979" />
                    <RANKING order="6" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6249" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3042" />
                    <RANKING order="2" place="2" resultid="3358" />
                    <RANKING order="3" place="3" resultid="3964" />
                    <RANKING order="4" place="4" resultid="4183" />
                    <RANKING order="5" place="5" resultid="1658" />
                    <RANKING order="6" place="6" resultid="3315" />
                    <RANKING order="7" place="7" resultid="3985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6250" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4427" />
                    <RANKING order="2" place="2" resultid="3394" />
                    <RANKING order="3" place="3" resultid="4616" />
                    <RANKING order="4" place="4" resultid="5516" />
                    <RANKING order="5" place="5" resultid="4219" />
                    <RANKING order="6" place="6" resultid="2825" />
                    <RANKING order="7" place="7" resultid="4310" />
                    <RANKING order="8" place="8" resultid="4839" />
                    <RANKING order="9" place="9" resultid="3187" />
                    <RANKING order="10" place="10" resultid="5452" />
                    <RANKING order="11" place="11" resultid="5002" />
                    <RANKING order="12" place="12" resultid="5056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6251" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5528" />
                    <RANKING order="2" place="2" resultid="5444" />
                    <RANKING order="3" place="3" resultid="4025" />
                    <RANKING order="4" place="4" resultid="4655" />
                    <RANKING order="5" place="5" resultid="3692" />
                    <RANKING order="6" place="6" resultid="3290" />
                    <RANKING order="7" place="7" resultid="4761" />
                    <RANKING order="8" place="8" resultid="4315" />
                    <RANKING order="9" place="9" resultid="3865" />
                    <RANKING order="10" place="10" resultid="3269" />
                    <RANKING order="11" place="-1" resultid="3614" />
                    <RANKING order="12" place="-1" resultid="4674" />
                    <RANKING order="13" place="-1" resultid="5007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6252" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3553" />
                    <RANKING order="2" place="2" resultid="4070" />
                    <RANKING order="3" place="3" resultid="3506" />
                    <RANKING order="4" place="4" resultid="2929" />
                    <RANKING order="5" place="5" resultid="3286" />
                    <RANKING order="6" place="6" resultid="4197" />
                    <RANKING order="7" place="7" resultid="4265" />
                    <RANKING order="8" place="8" resultid="4548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6253" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5282" />
                    <RANKING order="2" place="2" resultid="5031" />
                    <RANKING order="3" place="3" resultid="5026" />
                    <RANKING order="4" place="4" resultid="4043" />
                    <RANKING order="5" place="5" resultid="4935" />
                    <RANKING order="6" place="6" resultid="4446" />
                    <RANKING order="7" place="-1" resultid="3620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6254" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3304" />
                    <RANKING order="2" place="2" resultid="5315" />
                    <RANKING order="3" place="3" resultid="5262" />
                    <RANKING order="4" place="4" resultid="3212" />
                    <RANKING order="5" place="5" resultid="4663" />
                    <RANKING order="6" place="6" resultid="4400" />
                    <RANKING order="7" place="7" resultid="4029" />
                    <RANKING order="8" place="8" resultid="4668" />
                    <RANKING order="9" place="9" resultid="4406" />
                    <RANKING order="10" place="10" resultid="2936" />
                    <RANKING order="11" place="11" resultid="3706" />
                    <RANKING order="12" place="-1" resultid="3517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6255" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3406" />
                    <RANKING order="2" place="2" resultid="4590" />
                    <RANKING order="3" place="3" resultid="3237" />
                    <RANKING order="4" place="4" resultid="3037" />
                    <RANKING order="5" place="5" resultid="5417" />
                    <RANKING order="6" place="6" resultid="5569" />
                    <RANKING order="7" place="7" resultid="3709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6256" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4648" />
                    <RANKING order="2" place="2" resultid="3018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6257" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3339" />
                    <RANKING order="2" place="2" resultid="4464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6258" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5131" />
                    <RANKING order="2" place="2" resultid="3462" />
                    <RANKING order="3" place="3" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6259" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6260" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3499" />
                    <RANKING order="2" place="2" resultid="2774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6261" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5865" daytime="16:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5866" daytime="16:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5867" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5868" daytime="16:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5869" daytime="16:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5870" daytime="16:16" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5871" daytime="16:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5872" daytime="16:18" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5873" daytime="16:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5874" daytime="16:20" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1316" daytime="16:22" gender="F" number="16" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6262" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2992" />
                    <RANKING order="2" place="2" resultid="4913" />
                    <RANKING order="3" place="3" resultid="5423" />
                    <RANKING order="4" place="4" resultid="3434" />
                    <RANKING order="5" place="5" resultid="4939" />
                    <RANKING order="6" place="6" resultid="4830" />
                    <RANKING order="7" place="7" resultid="2792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6263" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2798" />
                    <RANKING order="2" place="2" resultid="4362" />
                    <RANKING order="3" place="3" resultid="3430" />
                    <RANKING order="4" place="4" resultid="3122" />
                    <RANKING order="5" place="5" resultid="3855" />
                    <RANKING order="6" place="6" resultid="4345" />
                    <RANKING order="7" place="7" resultid="4835" />
                    <RANKING order="8" place="-1" resultid="3006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6264" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3368" />
                    <RANKING order="2" place="2" resultid="3422" />
                    <RANKING order="3" place="3" resultid="3575" />
                    <RANKING order="4" place="4" resultid="3353" />
                    <RANKING order="5" place="5" resultid="5075" />
                    <RANKING order="6" place="6" resultid="4337" />
                    <RANKING order="7" place="7" resultid="5344" />
                    <RANKING order="8" place="8" resultid="5327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6265" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5015" />
                    <RANKING order="2" place="2" resultid="5298" />
                    <RANKING order="3" place="3" resultid="4877" />
                    <RANKING order="4" place="4" resultid="4104" />
                    <RANKING order="5" place="5" resultid="3931" />
                    <RANKING order="6" place="6" resultid="3725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6266" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4571" />
                    <RANKING order="2" place="2" resultid="4740" />
                    <RANKING order="3" place="3" resultid="5506" />
                    <RANKING order="4" place="4" resultid="3900" />
                    <RANKING order="5" place="5" resultid="3526" />
                    <RANKING order="6" place="6" resultid="3581" />
                    <RANKING order="7" place="7" resultid="4643" />
                    <RANKING order="8" place="8" resultid="3564" />
                    <RANKING order="9" place="-1" resultid="4578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6267" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4691" />
                    <RANKING order="2" place="2" resultid="3850" />
                    <RANKING order="3" place="3" resultid="4924" />
                    <RANKING order="4" place="4" resultid="3676" />
                    <RANKING order="5" place="5" resultid="2875" />
                    <RANKING order="6" place="6" resultid="4065" />
                    <RANKING order="7" place="7" resultid="4286" />
                    <RANKING order="8" place="-1" resultid="4765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6268" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4605" />
                    <RANKING order="2" place="2" resultid="4259" />
                    <RANKING order="3" place="3" resultid="2861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6269" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4018" />
                    <RANKING order="2" place="2" resultid="4610" />
                    <RANKING order="3" place="3" resultid="5070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6270" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4321" />
                    <RANKING order="2" place="2" resultid="3714" />
                    <RANKING order="3" place="3" resultid="3261" />
                    <RANKING order="4" place="4" resultid="5171" />
                    <RANKING order="5" place="5" resultid="4111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6271" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3234" />
                    <RANKING order="2" place="2" resultid="4239" />
                    <RANKING order="3" place="3" resultid="2915" />
                    <RANKING order="4" place="4" resultid="2909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6272" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5186" />
                    <RANKING order="2" place="2" resultid="3456" />
                    <RANKING order="3" place="3" resultid="5192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6273" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6274" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6275" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6276" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6277" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5875" daytime="16:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5876" daytime="16:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5877" daytime="16:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5878" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5879" daytime="16:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5880" daytime="16:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5881" daytime="16:38" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1333" daytime="16:40" gender="M" number="17" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6278" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5305" />
                    <RANKING order="2" place="2" resultid="3443" />
                    <RANKING order="3" place="3" resultid="3951" />
                    <RANKING order="4" place="4" resultid="3477" />
                    <RANKING order="5" place="5" resultid="3206" />
                    <RANKING order="6" place="6" resultid="3958" />
                    <RANKING order="7" place="-1" resultid="3220" />
                    <RANKING order="8" place="-1" resultid="4252" />
                    <RANKING order="9" place="-1" resultid="5648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6279" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4476" />
                    <RANKING order="2" place="2" resultid="4164" />
                    <RANKING order="3" place="3" resultid="4543" />
                    <RANKING order="4" place="4" resultid="2985" />
                    <RANKING order="5" place="5" resultid="4524" />
                    <RANKING order="6" place="6" resultid="2999" />
                    <RANKING order="7" place="7" resultid="4843" />
                    <RANKING order="8" place="8" resultid="4930" />
                    <RANKING order="9" place="9" resultid="3114" />
                    <RANKING order="10" place="10" resultid="3101" />
                    <RANKING order="11" place="11" resultid="3388" />
                    <RANKING order="12" place="-1" resultid="3281" />
                    <RANKING order="13" place="-1" resultid="5723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6280" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5121" />
                    <RANKING order="2" place="2" resultid="5021" />
                    <RANKING order="3" place="3" resultid="3265" />
                    <RANKING order="4" place="4" resultid="3570" />
                    <RANKING order="5" place="5" resultid="4077" />
                    <RANKING order="6" place="6" resultid="3944" />
                    <RANKING order="7" place="7" resultid="2732" />
                    <RANKING order="8" place="8" resultid="4773" />
                    <RANKING order="9" place="-1" resultid="3972" />
                    <RANKING order="10" place="-1" resultid="3993" />
                    <RANKING order="11" place="-1" resultid="4272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6281" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3043" />
                    <RANKING order="2" place="2" resultid="3687" />
                    <RANKING order="3" place="3" resultid="4750" />
                    <RANKING order="4" place="4" resultid="3030" />
                    <RANKING order="5" place="5" resultid="3965" />
                    <RANKING order="6" place="6" resultid="3323" />
                    <RANKING order="7" place="7" resultid="3874" />
                    <RANKING order="8" place="8" resultid="3131" />
                    <RANKING order="9" place="9" resultid="3986" />
                    <RANKING order="10" place="10" resultid="1659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6282" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3731" />
                    <RANKING order="2" place="2" resultid="4617" />
                    <RANKING order="3" place="3" resultid="4470" />
                    <RANKING order="4" place="4" resultid="3049" />
                    <RANKING order="5" place="5" resultid="4685" />
                    <RANKING order="6" place="6" resultid="2826" />
                    <RANKING order="7" place="7" resultid="4813" />
                    <RANKING order="8" place="8" resultid="5453" />
                    <RANKING order="9" place="9" resultid="2812" />
                    <RANKING order="10" place="10" resultid="5226" />
                    <RANKING order="11" place="11" resultid="3148" />
                    <RANKING order="12" place="12" resultid="5045" />
                    <RANKING order="13" place="13" resultid="4680" />
                    <RANKING order="14" place="14" resultid="3076" />
                    <RANKING order="15" place="15" resultid="3188" />
                    <RANKING order="16" place="16" resultid="3182" />
                    <RANKING order="17" place="-1" resultid="2758" />
                    <RANKING order="18" place="-1" resultid="5231" />
                    <RANKING order="19" place="-1" resultid="5517" />
                    <RANKING order="20" place="-1" resultid="5521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6283" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2854" />
                    <RANKING order="2" place="2" resultid="3547" />
                    <RANKING order="3" place="3" resultid="4529" />
                    <RANKING order="4" place="4" resultid="4316" />
                    <RANKING order="5" place="5" resultid="4011" />
                    <RANKING order="6" place="6" resultid="5389" />
                    <RANKING order="7" place="-1" resultid="3615" />
                    <RANKING order="8" place="-1" resultid="4769" />
                    <RANKING order="9" place="-1" resultid="5361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6284" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                    <RANKING order="2" place="2" resultid="5237" />
                    <RANKING order="3" place="3" resultid="5257" />
                    <RANKING order="4" place="4" resultid="4071" />
                    <RANKING order="5" place="5" resultid="3630" />
                    <RANKING order="6" place="6" resultid="4973" />
                    <RANKING order="7" place="7" resultid="4629" />
                    <RANKING order="8" place="8" resultid="3383" />
                    <RANKING order="9" place="9" resultid="4266" />
                    <RANKING order="10" place="-1" resultid="3491" />
                    <RANKING order="11" place="-1" resultid="3698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6285" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3379" />
                    <RANKING order="2" place="2" resultid="5283" />
                    <RANKING order="3" place="3" resultid="5032" />
                    <RANKING order="4" place="4" resultid="4585" />
                    <RANKING order="5" place="5" resultid="4791" />
                    <RANKING order="6" place="6" resultid="4051" />
                    <RANKING order="7" place="7" resultid="2847" />
                    <RANKING order="8" place="8" resultid="3895" />
                    <RANKING order="9" place="9" resultid="4447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6286" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2786" />
                    <RANKING order="2" place="2" resultid="4353" />
                    <RANKING order="3" place="3" resultid="3305" />
                    <RANKING order="4" place="4" resultid="4214" />
                    <RANKING order="5" place="5" resultid="3213" />
                    <RANKING order="6" place="6" resultid="5219" />
                    <RANKING order="7" place="7" resultid="4669" />
                    <RANKING order="8" place="8" resultid="4411" />
                    <RANKING order="9" place="9" resultid="3884" />
                    <RANKING order="10" place="-1" resultid="3518" />
                    <RANKING order="11" place="-1" resultid="4407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6287" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3407" />
                    <RANKING order="2" place="2" resultid="4944" />
                    <RANKING order="3" place="3" resultid="5147" />
                    <RANKING order="4" place="4" resultid="4514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6288" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4711" />
                    <RANKING order="2" place="2" resultid="5141" />
                    <RANKING order="3" place="3" resultid="2923" />
                    <RANKING order="4" place="4" resultid="5752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6289" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3340" />
                    <RANKING order="2" place="2" resultid="4465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6290" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3463" />
                    <RANKING order="2" place="-1" resultid="5738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6291" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6292" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6293" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5882" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5883" daytime="16:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5884" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5885" daytime="16:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5886" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5887" daytime="16:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5888" daytime="16:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5889" daytime="16:56" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5890" daytime="16:58" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5891" daytime="17:00" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5892" daytime="17:02" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5893" daytime="17:04" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" daytime="17:06" gender="F" number="18" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6294" agemax="24" agemin="20" name="Kategoria 0" />
                <AGEGROUP agegroupid="6295" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="6296" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3533" />
                    <RANKING order="2" place="2" resultid="5510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6297" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3660" />
                    <RANKING order="2" place="2" resultid="4395" />
                    <RANKING order="3" place="3" resultid="3176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6298" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3152" />
                    <RANKING order="2" place="2" resultid="3162" />
                    <RANKING order="3" place="-1" resultid="5759" />
                    <RANKING order="4" place="-1" resultid="5374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6299" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6300" agemax="54" agemin="50" name="Kategoria F" />
                <AGEGROUP agegroupid="6301" agemax="59" agemin="55" name="Kategoria G" />
                <AGEGROUP agegroupid="6302" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6303" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="6304" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="6305" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6306" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6307" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6308" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6309" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5894" daytime="17:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5895" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1367" daytime="17:16" gender="M" number="19" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6310" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5653" />
                    <RANKING order="2" place="2" resultid="3296" />
                    <RANKING order="3" place="3" resultid="4369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6311" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6312" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5354" />
                    <RANKING order="2" place="2" resultid="3845" />
                    <RANKING order="3" place="3" resultid="4127" />
                    <RANKING order="4" place="4" resultid="3241" />
                    <RANKING order="5" place="5" resultid="5395" />
                    <RANKING order="6" place="6" resultid="3311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6313" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5052" />
                    <RANKING order="2" place="2" resultid="4184" />
                    <RANKING order="3" place="-1" resultid="4956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6314" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2805" />
                    <RANKING order="2" place="2" resultid="5522" />
                    <RANKING order="3" place="3" resultid="4487" />
                    <RANKING order="4" place="4" resultid="4686" />
                    <RANKING order="5" place="5" resultid="3702" />
                    <RANKING order="6" place="-1" resultid="3169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6315" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4171" />
                    <RANKING order="2" place="2" resultid="4890" />
                    <RANKING order="3" place="3" resultid="5099" />
                    <RANKING order="4" place="4" resultid="4292" />
                    <RANKING order="5" place="5" resultid="3539" />
                    <RANKING order="6" place="6" resultid="3560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6316" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4974" />
                    <RANKING order="2" place="2" resultid="4384" />
                    <RANKING order="3" place="3" resultid="4756" />
                    <RANKING order="4" place="4" resultid="1666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6317" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4433" />
                    <RANKING order="2" place="2" resultid="3092" />
                    <RANKING order="3" place="3" resultid="4245" />
                    <RANKING order="4" place="4" resultid="4723" />
                    <RANKING order="5" place="-1" resultid="2869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6318" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4391" />
                    <RANKING order="2" place="2" resultid="4030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6319" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5731" />
                    <RANKING order="2" place="2" resultid="4701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6320" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5753" />
                    <RANKING order="2" place="2" resultid="4037" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="-1" resultid="3056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6321" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6322" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6323" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6324" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6325" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5896" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5897" daytime="17:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5898" daytime="17:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5899" daytime="17:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5900" daytime="17:36" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1384" daytime="17:40" gender="F" number="20" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6326" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6327" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4558" />
                    <RANKING order="2" place="2" resultid="3347" />
                    <RANKING order="3" place="3" resultid="4898" />
                    <RANKING order="4" place="4" resultid="5080" />
                    <RANKING order="5" place="5" resultid="4346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6328" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5250" />
                    <RANKING order="2" place="2" resultid="3682" />
                    <RANKING order="3" place="3" resultid="5511" />
                    <RANKING order="4" place="-1" resultid="4805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6329" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5299" />
                    <RANKING order="2" place="2" resultid="3661" />
                    <RANKING order="3" place="3" resultid="4105" />
                    <RANKING order="4" place="4" resultid="3932" />
                    <RANKING order="5" place="-1" resultid="3645" />
                    <RANKING order="6" place="-1" resultid="4707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6330" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3901" />
                    <RANKING order="2" place="2" resultid="5321" />
                    <RANKING order="3" place="3" resultid="3163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6331" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6332" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6333" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4482" />
                    <RANKING order="2" place="2" resultid="2962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6334" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4322" />
                    <RANKING order="2" place="2" resultid="5164" />
                    <RANKING order="3" place="3" resultid="3890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6335" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3069" />
                    <RANKING order="2" place="2" resultid="2916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6336" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="6337" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6338" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6339" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6340" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6341" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5901" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5902" daytime="17:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5903" daytime="17:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1401" daytime="17:56" gender="M" number="21" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6342" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4884" />
                    <RANKING order="2" place="2" resultid="3444" />
                    <RANKING order="3" place="3" resultid="3297" />
                    <RANKING order="4" place="4" resultid="2740" />
                    <RANKING order="5" place="5" resultid="3221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6343" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4165" />
                    <RANKING order="2" place="2" resultid="5534" />
                    <RANKING order="3" place="3" resultid="3275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6344" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6345" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3031" />
                    <RANKING order="2" place="2" resultid="5243" />
                    <RANKING order="3" place="-1" resultid="5468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6346" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                    <RANKING order="2" place="2" resultid="5046" />
                    <RANKING order="3" place="3" resultid="4226" />
                    <RANKING order="4" place="-1" resultid="2759" />
                    <RANKING order="5" place="-1" resultid="3050" />
                    <RANKING order="6" place="-1" resultid="4995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6347" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4453" />
                    <RANKING order="2" place="2" resultid="4327" />
                    <RANKING order="3" place="3" resultid="4178" />
                    <RANKING order="4" place="4" resultid="4848" />
                    <RANKING order="5" place="5" resultid="3540" />
                    <RANKING order="6" place="6" resultid="4203" />
                    <RANKING order="7" place="-1" resultid="5008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6348" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2883" />
                    <RANKING order="2" place="2" resultid="2930" />
                    <RANKING order="3" place="3" resultid="4951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6349" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4459" />
                    <RANKING order="2" place="2" resultid="4044" />
                    <RANKING order="3" place="3" resultid="3093" />
                    <RANKING order="4" place="4" resultid="3137" />
                    <RANKING order="5" place="-1" resultid="4724" />
                    <RANKING order="6" place="-1" resultid="4810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6350" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4354" />
                    <RANKING order="2" place="2" resultid="4870" />
                    <RANKING order="3" place="3" resultid="5039" />
                    <RANKING order="4" place="4" resultid="4695" />
                    <RANKING order="5" place="-1" resultid="4412" />
                    <RANKING order="6" place="-1" resultid="4624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6351" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4945" />
                    <RANKING order="2" place="2" resultid="5732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6352" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4649" />
                    <RANKING order="2" place="2" resultid="5127" />
                    <RANKING order="3" place="3" resultid="2943" />
                    <RANKING order="4" place="4" resultid="3057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6353" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6354" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3063" />
                    <RANKING order="2" place="2" resultid="5746" />
                    <RANKING order="3" place="-1" resultid="5739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6355" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6356" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6357" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5904" daytime="17:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5905" daytime="18:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5906" daytime="18:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5907" daytime="18:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5908" daytime="18:14" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1418" daytime="18:18" gender="F" number="22" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6518" agemax="-1" agemin="-1" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6519" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL" />
                <AGEGROUP agegroupid="6520" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3450" />
                    <RANKING order="2" place="2" resultid="3914" />
                    <RANKING order="3" place="3" resultid="3740" />
                    <RANKING order="4" place="4" resultid="5082" />
                    <RANKING order="5" place="5" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6521" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3719" />
                    <RANKING order="2" place="2" resultid="5332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6522" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4729" />
                    <RANKING order="2" place="2" resultid="4115" />
                    <RANKING order="3" place="3" resultid="3912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6523" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL" />
                <AGEGROUP agegroupid="6524" agemax="-1" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5195" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5909" daytime="18:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5910" daytime="18:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1442" daytime="18:24" gender="M" number="23" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6525" agemax="-1" agemin="-1" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6526" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5725" />
                    <RANKING order="2" place="2" resultid="5765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6527" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5060" />
                    <RANKING order="2" place="2" resultid="4229" />
                    <RANKING order="3" place="3" resultid="3736" />
                    <RANKING order="4" place="4" resultid="4538" />
                    <RANKING order="5" place="5" resultid="2833" />
                    <RANKING order="6" place="6" resultid="4964" />
                    <RANKING order="7" place="7" resultid="3996" />
                    <RANKING order="8" place="-1" resultid="3078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6528" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4490" />
                    <RANKING order="2" place="2" resultid="5564" />
                    <RANKING order="3" place="3" resultid="5334" />
                    <RANKING order="4" place="4" resultid="3588" />
                    <RANKING order="5" place="5" resultid="4230" />
                    <RANKING order="6" place="6" resultid="5061" />
                    <RANKING order="7" place="7" resultid="5335" />
                    <RANKING order="8" place="8" resultid="5221" />
                    <RANKING order="9" place="9" resultid="3192" />
                    <RANKING order="10" place="10" resultid="4119" />
                    <RANKING order="11" place="11" resultid="4775" />
                    <RANKING order="12" place="12" resultid="3721" />
                    <RANKING order="13" place="13" resultid="3916" />
                    <RANKING order="14" place="-1" resultid="4730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6529" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4491" />
                    <RANKING order="2" place="2" resultid="3737" />
                    <RANKING order="3" place="3" resultid="4280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6530" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4731" />
                    <RANKING order="2" place="-1" resultid="4117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6531" agemax="-1" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5196" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5911" daytime="18:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5912" daytime="18:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5913" daytime="18:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5914" daytime="18:34" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-12-12" daytime="08:30" number="3">
          <EVENTS>
            <EVENT eventid="1451" daytime="08:30" gender="F" number="24" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6358" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2993" />
                    <RANKING order="2" place="2" resultid="3435" />
                    <RANKING order="3" place="3" resultid="3650" />
                    <RANKING order="4" place="4" resultid="3438" />
                    <RANKING order="5" place="5" resultid="4940" />
                    <RANKING order="6" place="6" resultid="4831" />
                    <RANKING order="7" place="7" resultid="5439" />
                    <RANKING order="8" place="-1" resultid="4721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6359" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="2799" />
                    <RANKING order="3" place="3" resultid="4363" />
                    <RANKING order="4" place="4" resultid="3881" />
                    <RANKING order="5" place="5" resultid="3123" />
                    <RANKING order="6" place="6" resultid="4836" />
                    <RANKING order="7" place="7" resultid="3007" />
                    <RANKING order="8" place="-1" resultid="3348" />
                    <RANKING order="9" place="-1" resultid="3856" />
                    <RANKING order="10" place="-1" resultid="4347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6360" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3369" />
                    <RANKING order="2" place="2" resultid="3354" />
                    <RANKING order="3" place="3" resultid="4338" />
                    <RANKING order="4" place="4" resultid="3228" />
                    <RANKING order="5" place="5" resultid="3623" />
                    <RANKING order="6" place="-1" resultid="5512" />
                    <RANKING order="7" place="-1" resultid="5641" />
                    <RANKING order="8" place="-1" resultid="5762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6361" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4878" />
                    <RANKING order="2" place="2" resultid="5300" />
                    <RANKING order="3" place="3" resultid="3609" />
                    <RANKING order="4" place="-1" resultid="3726" />
                    <RANKING order="5" place="-1" resultid="5016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6362" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4572" />
                    <RANKING order="2" place="2" resultid="4741" />
                    <RANKING order="3" place="3" resultid="3144" />
                    <RANKING order="4" place="4" resultid="4782" />
                    <RANKING order="5" place="5" resultid="3582" />
                    <RANKING order="6" place="6" resultid="2957" />
                    <RANKING order="7" place="7" resultid="3449" />
                    <RANKING order="8" place="8" resultid="4579" />
                    <RANKING order="9" place="9" resultid="5093" />
                    <RANKING order="10" place="-1" resultid="2951" />
                    <RANKING order="11" place="-1" resultid="3565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6363" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3851" />
                    <RANKING order="2" place="2" resultid="4305" />
                    <RANKING order="3" place="3" resultid="3677" />
                    <RANKING order="4" place="4" resultid="3668" />
                    <RANKING order="5" place="5" resultid="3673" />
                    <RANKING order="6" place="6" resultid="4422" />
                    <RANKING order="7" place="7" resultid="3869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6364" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2862" />
                    <RANKING order="2" place="2" resultid="2969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6365" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4019" />
                    <RANKING order="2" place="2" resultid="4611" />
                    <RANKING order="3" place="3" resultid="4862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6366" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4059" />
                    <RANKING order="2" place="2" resultid="4595" />
                    <RANKING order="3" place="3" resultid="3262" />
                    <RANKING order="4" place="4" resultid="3862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6367" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4903" />
                    <RANKING order="2" place="2" resultid="5402" />
                    <RANKING order="3" place="3" resultid="4240" />
                    <RANKING order="4" place="4" resultid="4855" />
                    <RANKING order="5" place="5" resultid="2910" />
                    <RANKING order="6" place="6" resultid="2917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6368" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3457" />
                    <RANKING order="2" place="2" resultid="5425" />
                    <RANKING order="3" place="3" resultid="4919" />
                    <RANKING order="4" place="4" resultid="2896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6369" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2903" />
                    <RANKING order="2" place="2" resultid="4095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6370" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6371" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6372" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6373" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5915" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5916" daytime="08:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5917" daytime="08:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5918" daytime="08:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5919" daytime="08:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5920" daytime="08:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5921" daytime="08:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5922" daytime="08:40" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1469" daytime="08:42" gender="M" number="25" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6374" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5306" />
                    <RANKING order="2" place="2" resultid="4376" />
                    <RANKING order="3" place="3" resultid="4885" />
                    <RANKING order="4" place="4" resultid="4826" />
                    <RANKING order="5" place="5" resultid="3640" />
                    <RANKING order="6" place="6" resultid="5201" />
                    <RANKING order="7" place="7" resultid="3952" />
                    <RANKING order="8" place="8" resultid="3025" />
                    <RANKING order="9" place="9" resultid="3478" />
                    <RANKING order="10" place="10" resultid="3207" />
                    <RANKING order="11" place="-1" resultid="4253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6375" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4477" />
                    <RANKING order="2" place="2" resultid="3908" />
                    <RANKING order="3" place="3" resultid="4525" />
                    <RANKING order="4" place="4" resultid="2986" />
                    <RANKING order="5" place="5" resultid="4544" />
                    <RANKING order="6" place="6" resultid="5541" />
                    <RANKING order="7" place="7" resultid="4563" />
                    <RANKING order="8" place="8" resultid="3102" />
                    <RANKING order="9" place="9" resultid="4566" />
                    <RANKING order="10" place="10" resultid="3282" />
                    <RANKING order="11" place="11" resultid="4931" />
                    <RANKING order="12" place="12" resultid="4499" />
                    <RANKING order="13" place="13" resultid="2821" />
                    <RANKING order="14" place="14" resultid="5368" />
                    <RANKING order="15" place="15" resultid="5349" />
                    <RANKING order="16" place="16" resultid="4083" />
                    <RANKING order="17" place="17" resultid="5382" />
                    <RANKING order="18" place="-1" resultid="3000" />
                    <RANKING order="19" place="-1" resultid="3389" />
                    <RANKING order="20" place="-1" resultid="4133" />
                    <RANKING order="21" place="-1" resultid="4844" />
                    <RANKING order="22" place="-1" resultid="5535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6376" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4438" />
                    <RANKING order="2" place="2" resultid="3266" />
                    <RANKING order="3" place="3" resultid="3512" />
                    <RANKING order="4" place="4" resultid="2733" />
                    <RANKING order="5" place="5" resultid="2974" />
                    <RANKING order="6" place="6" resultid="3945" />
                    <RANKING order="7" place="7" resultid="4136" />
                    <RANKING order="8" place="8" resultid="3110" />
                    <RANKING order="9" place="9" resultid="4774" />
                    <RANKING order="10" place="10" resultid="3980" />
                    <RANKING order="11" place="11" resultid="5110" />
                    <RANKING order="12" place="12" resultid="3973" />
                    <RANKING order="13" place="-1" resultid="3994" />
                    <RANKING order="14" place="-1" resultid="4209" />
                    <RANKING order="15" place="-1" resultid="4273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6377" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5059" />
                    <RANKING order="2" place="2" resultid="4536" />
                    <RANKING order="3" place="3" resultid="5053" />
                    <RANKING order="4" place="4" resultid="4785" />
                    <RANKING order="5" place="5" resultid="4751" />
                    <RANKING order="6" place="6" resultid="5207" />
                    <RANKING order="7" place="7" resultid="5211" />
                    <RANKING order="8" place="8" resultid="3359" />
                    <RANKING order="9" place="9" resultid="4191" />
                    <RANKING order="10" place="10" resultid="3966" />
                    <RANKING order="11" place="11" resultid="5350" />
                    <RANKING order="12" place="12" resultid="3875" />
                    <RANKING order="13" place="13" resultid="3987" />
                    <RANKING order="14" place="14" resultid="3925" />
                    <RANKING order="15" place="-1" resultid="3401" />
                    <RANKING order="16" place="-1" resultid="4278" />
                    <RANKING order="17" place="-1" resultid="4909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6378" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3732" />
                    <RANKING order="2" place="2" resultid="5523" />
                    <RANKING order="3" place="3" resultid="4428" />
                    <RANKING order="4" place="4" resultid="3395" />
                    <RANKING order="5" place="5" resultid="5518" />
                    <RANKING order="6" place="6" resultid="3051" />
                    <RANKING order="7" place="7" resultid="4471" />
                    <RANKING order="8" place="8" resultid="4618" />
                    <RANKING order="9" place="9" resultid="4509" />
                    <RANKING order="10" place="10" resultid="2831" />
                    <RANKING order="11" place="11" resultid="3170" />
                    <RANKING order="12" place="12" resultid="4220" />
                    <RANKING order="13" place="13" resultid="5454" />
                    <RANKING order="14" place="14" resultid="5216" />
                    <RANKING order="15" place="15" resultid="3189" />
                    <RANKING order="16" place="16" resultid="3149" />
                    <RANKING order="17" place="17" resultid="5003" />
                    <RANKING order="18" place="18" resultid="3077" />
                    <RANKING order="19" place="19" resultid="4681" />
                    <RANKING order="20" place="20" resultid="3921" />
                    <RANKING order="21" place="21" resultid="5057" />
                    <RANKING order="22" place="22" resultid="5562" />
                    <RANKING order="23" place="23" resultid="5106" />
                    <RANKING order="24" place="-1" resultid="4996" />
                    <RANKING order="25" place="-1" resultid="5232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6379" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4172" />
                    <RANKING order="2" place="2" resultid="2855" />
                    <RANKING order="3" place="3" resultid="4797" />
                    <RANKING order="4" place="4" resultid="2880" />
                    <RANKING order="5" place="5" resultid="3548" />
                    <RANKING order="6" place="6" resultid="4530" />
                    <RANKING order="7" place="7" resultid="4333" />
                    <RANKING order="8" place="8" resultid="4819" />
                    <RANKING order="9" place="9" resultid="4520" />
                    <RANKING order="10" place="10" resultid="3541" />
                    <RANKING order="11" place="11" resultid="4849" />
                    <RANKING order="12" place="12" resultid="4012" />
                    <RANKING order="13" place="13" resultid="5553" />
                    <RANKING order="14" place="14" resultid="4204" />
                    <RANKING order="15" place="15" resultid="3866" />
                    <RANKING order="16" place="-1" resultid="3655" />
                    <RANKING order="17" place="-1" resultid="4675" />
                    <RANKING order="18" place="-1" resultid="5009" />
                    <RANKING order="19" place="-1" resultid="5116" />
                    <RANKING order="20" place="-1" resultid="5362" />
                    <RANKING order="21" place="-1" resultid="5390" />
                    <RANKING order="22" place="-1" resultid="5529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6380" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4072" />
                    <RANKING order="2" place="2" resultid="5258" />
                    <RANKING order="3" place="3" resultid="3631" />
                    <RANKING order="4" place="4" resultid="3012" />
                    <RANKING order="5" place="5" resultid="4385" />
                    <RANKING order="6" place="6" resultid="4952" />
                    <RANKING order="7" place="7" resultid="4630" />
                    <RANKING order="8" place="8" resultid="3699" />
                    <RANKING order="9" place="9" resultid="4198" />
                    <RANKING order="10" place="10" resultid="4757" />
                    <RANKING order="11" place="11" resultid="4267" />
                    <RANKING order="12" place="12" resultid="4549" />
                    <RANKING order="13" place="13" resultid="1667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6381" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="5033" />
                    <RANKING order="3" place="3" resultid="4586" />
                    <RANKING order="4" place="4" resultid="4792" />
                    <RANKING order="5" place="5" resultid="5463" />
                    <RANKING order="6" place="6" resultid="4052" />
                    <RANKING order="7" place="7" resultid="3896" />
                    <RANKING order="8" place="8" resultid="2848" />
                    <RANKING order="9" place="9" resultid="5459" />
                    <RANKING order="10" place="10" resultid="2870" />
                    <RANKING order="11" place="11" resultid="3138" />
                    <RANKING order="12" place="12" resultid="2781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6382" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3306" />
                    <RANKING order="2" place="2" resultid="4625" />
                    <RANKING order="3" place="3" resultid="4717" />
                    <RANKING order="4" place="4" resultid="3214" />
                    <RANKING order="5" place="5" resultid="4670" />
                    <RANKING order="6" place="6" resultid="4413" />
                    <RANKING order="7" place="7" resultid="4401" />
                    <RANKING order="8" place="8" resultid="3519" />
                    <RANKING order="9" place="9" resultid="4408" />
                    <RANKING order="10" place="10" resultid="3363" />
                    <RANKING order="11" place="11" resultid="2937" />
                    <RANKING order="12" place="12" resultid="3707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6383" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3038" />
                    <RANKING order="2" place="2" resultid="4961" />
                    <RANKING order="3" place="3" resultid="4515" />
                    <RANKING order="4" place="4" resultid="4591" />
                    <RANKING order="5" place="5" resultid="5148" />
                    <RANKING order="6" place="6" resultid="2767" />
                    <RANKING order="7" place="7" resultid="5418" />
                    <RANKING order="8" place="8" resultid="3710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6384" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5142" />
                    <RANKING order="2" place="2" resultid="4038" />
                    <RANKING order="3" place="3" resultid="4554" />
                    <RANKING order="4" place="4" resultid="2924" />
                    <RANKING order="5" place="5" resultid="2752" />
                    <RANKING order="6" place="6" resultid="2944" />
                    <RANKING order="7" place="7" resultid="1680" />
                    <RANKING order="8" place="8" resultid="4712" />
                    <RANKING order="9" place="9" resultid="3019" />
                    <RANKING order="10" place="-1" resultid="5182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6385" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3341" />
                    <RANKING order="2" place="2" resultid="4466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6386" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5158" />
                    <RANKING order="2" place="2" resultid="3064" />
                    <RANKING order="3" place="3" resultid="4088" />
                    <RANKING order="4" place="4" resultid="3464" />
                    <RANKING order="5" place="5" resultid="5747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6387" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6388" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6389" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5923" daytime="08:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5924" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5925" daytime="08:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5926" daytime="08:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5927" daytime="08:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5928" daytime="08:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5929" daytime="08:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5930" daytime="08:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5931" daytime="08:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5932" daytime="08:54" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5933" daytime="08:56" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5934" daytime="08:58" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5935" daytime="08:58" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5936" daytime="09:00" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="5937" daytime="09:00" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="5938" daytime="09:02" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="5939" daytime="09:02" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="5940" daytime="09:04" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1486" daytime="09:06" gender="F" number="26" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6390" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4914" />
                    <RANKING order="2" place="2" resultid="5312" />
                    <RANKING order="3" place="3" resultid="5424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6391" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2800" />
                    <RANKING order="2" place="2" resultid="3606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6392" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3534" />
                    <RANKING order="2" place="2" resultid="3624" />
                    <RANKING order="3" place="3" resultid="5328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6393" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5086" />
                    <RANKING order="2" place="2" resultid="5431" />
                    <RANKING order="3" place="3" resultid="4101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6394" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5375" />
                    <RANKING order="2" place="2" resultid="3527" />
                    <RANKING order="3" place="3" resultid="4644" />
                    <RANKING order="4" place="4" resultid="3164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6395" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5179" />
                    <RANKING order="2" place="2" resultid="4925" />
                    <RANKING order="3" place="3" resultid="2876" />
                    <RANKING order="4" place="4" resultid="4288" />
                    <RANKING order="5" place="5" resultid="4423" />
                    <RANKING order="6" place="6" resultid="4443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6396" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="2863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6397" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6398" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3891" />
                    <RANKING order="2" place="2" resultid="3715" />
                    <RANKING order="3" place="3" resultid="5172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6399" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5403" />
                    <RANKING order="2" place="2" resultid="4856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6400" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5193" />
                    <RANKING order="2" place="2" resultid="2897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6401" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6402" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6403" agemax="89" agemin="85" name="Kategoria M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6404" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6405" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5941" daytime="09:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5942" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5943" daytime="09:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5944" daytime="09:24" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1503" daytime="09:30" gender="M" number="27" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6406" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3298" />
                    <RANKING order="2" place="2" resultid="3959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6407" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4987" />
                    <RANKING order="2" place="2" resultid="3001" />
                    <RANKING order="3" place="3" resultid="3115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6408" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3571" />
                    <RANKING order="2" place="2" resultid="4128" />
                    <RANKING order="3" place="-1" resultid="4274" />
                    <RANKING order="4" place="-1" resultid="5397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6409" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3044" />
                    <RANKING order="2" place="2" resultid="5244" />
                    <RANKING order="3" place="3" resultid="1660" />
                    <RANKING order="4" place="-1" resultid="4185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6410" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2806" />
                    <RANKING order="2" place="2" resultid="4687" />
                    <RANKING order="3" place="3" resultid="2827" />
                    <RANKING order="4" place="4" resultid="4311" />
                    <RANKING order="5" place="5" resultid="4221" />
                    <RANKING order="6" place="6" resultid="3190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6411" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4891" />
                    <RANKING order="2" place="2" resultid="5445" />
                    <RANKING order="3" place="3" resultid="4026" />
                    <RANKING order="4" place="4" resultid="3693" />
                    <RANKING order="5" place="5" resultid="3291" />
                    <RANKING order="6" place="6" resultid="4317" />
                    <RANKING order="7" place="7" resultid="4656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6412" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3555" />
                    <RANKING order="2" place="2" resultid="3507" />
                    <RANKING order="3" place="3" resultid="3287" />
                    <RANKING order="4" place="-1" resultid="2931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6413" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5284" />
                    <RANKING order="2" place="2" resultid="5027" />
                    <RANKING order="3" place="3" resultid="4936" />
                    <RANKING order="4" place="4" resultid="4448" />
                    <RANKING order="5" place="5" resultid="5288" />
                    <RANKING order="6" place="6" resultid="4053" />
                    <RANKING order="7" place="7" resultid="4246" />
                    <RANKING order="8" place="-1" resultid="3621" />
                    <RANKING order="9" place="-1" resultid="5034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6414" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2787" />
                    <RANKING order="2" place="2" resultid="5316" />
                    <RANKING order="3" place="3" resultid="5263" />
                    <RANKING order="4" place="4" resultid="4215" />
                    <RANKING order="5" place="5" resultid="4031" />
                    <RANKING order="6" place="6" resultid="4402" />
                    <RANKING order="7" place="7" resultid="4664" />
                    <RANKING order="8" place="8" resultid="2938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6415" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3408" />
                    <RANKING order="2" place="2" resultid="3238" />
                    <RANKING order="3" place="3" resultid="5570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6416" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4650" />
                    <RANKING order="2" place="2" resultid="5754" />
                    <RANKING order="3" place="3" resultid="3020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6417" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6418" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6419" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6420" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6421" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5945" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5946" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5947" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5948" daytime="09:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5949" daytime="09:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5950" daytime="09:52" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1520" daytime="09:56" gender="F" number="28" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6422" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6423" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3349" />
                    <RANKING order="2" place="2" resultid="3882" />
                    <RANKING order="3" place="3" resultid="4899" />
                    <RANKING order="4" place="4" resultid="3857" />
                    <RANKING order="5" place="5" resultid="3124" />
                    <RANKING order="6" place="-1" resultid="4348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6424" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5251" />
                    <RANKING order="2" place="2" resultid="3683" />
                    <RANKING order="3" place="3" resultid="3576" />
                    <RANKING order="4" place="4" resultid="3229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6425" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5301" />
                    <RANKING order="2" place="2" resultid="4879" />
                    <RANKING order="3" place="3" resultid="3662" />
                    <RANKING order="4" place="4" resultid="4106" />
                    <RANKING order="5" place="5" resultid="3177" />
                    <RANKING order="6" place="6" resultid="3933" />
                    <RANKING order="7" place="7" resultid="3610" />
                    <RANKING order="8" place="-1" resultid="5017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6426" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4573" />
                    <RANKING order="2" place="2" resultid="3902" />
                    <RANKING order="3" place="3" resultid="5322" />
                    <RANKING order="4" place="-1" resultid="2952" />
                    <RANKING order="5" place="-1" resultid="3583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6427" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4692" />
                    <RANKING order="2" place="2" resultid="4766" />
                    <RANKING order="3" place="3" resultid="4066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6428" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6429" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4020" />
                    <RANKING order="2" place="2" resultid="4863" />
                    <RANKING order="3" place="3" resultid="4483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6430" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4323" />
                    <RANKING order="2" place="2" resultid="5165" />
                    <RANKING order="3" place="3" resultid="4596" />
                    <RANKING order="4" place="4" resultid="4112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6431" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4241" />
                    <RANKING order="2" place="2" resultid="4904" />
                    <RANKING order="3" place="3" resultid="3070" />
                    <RANKING order="4" place="4" resultid="2911" />
                    <RANKING order="5" place="5" resultid="2918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6432" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5187" />
                    <RANKING order="2" place="2" resultid="3458" />
                    <RANKING order="3" place="3" resultid="5154" />
                    <RANKING order="4" place="4" resultid="4920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6433" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2904" />
                    <RANKING order="2" place="2" resultid="4096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6434" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6435" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6436" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6437" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5951" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5952" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5953" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5954" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5955" daytime="10:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1537" daytime="10:12" gender="M" number="29" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6438" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4886" />
                    <RANKING order="2" place="2" resultid="3445" />
                    <RANKING order="3" place="3" resultid="2741" />
                    <RANKING order="4" place="4" resultid="3222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6439" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5536" />
                    <RANKING order="2" place="2" resultid="3276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6440" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5122" />
                    <RANKING order="2" place="2" resultid="2975" />
                    <RANKING order="3" place="3" resultid="4078" />
                    <RANKING order="4" place="-1" resultid="3974" />
                    <RANKING order="5" place="-1" resultid="3995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6441" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3402" />
                    <RANKING order="2" place="2" resultid="3688" />
                    <RANKING order="3" place="3" resultid="5212" />
                    <RANKING order="4" place="4" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6442" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3733" />
                    <RANKING order="2" place="2" resultid="3158" />
                    <RANKING order="3" place="3" resultid="3052" />
                    <RANKING order="4" place="4" resultid="4472" />
                    <RANKING order="5" place="5" resultid="4619" />
                    <RANKING order="6" place="6" resultid="4227" />
                    <RANKING order="7" place="7" resultid="5047" />
                    <RANKING order="8" place="8" resultid="4814" />
                    <RANKING order="9" place="9" resultid="2813" />
                    <RANKING order="10" place="10" resultid="3635" />
                    <RANKING order="11" place="-1" resultid="2760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6443" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4454" />
                    <RANKING order="2" place="2" resultid="4531" />
                    <RANKING order="3" place="3" resultid="4328" />
                    <RANKING order="4" place="4" resultid="4762" />
                    <RANKING order="5" place="5" resultid="4850" />
                    <RANKING order="6" place="-1" resultid="4205" />
                    <RANKING order="7" place="-1" resultid="4770" />
                    <RANKING order="8" place="-1" resultid="5100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6444" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2884" />
                    <RANKING order="2" place="2" resultid="3492" />
                    <RANKING order="3" place="3" resultid="4953" />
                    <RANKING order="4" place="4" resultid="4550" />
                    <RANKING order="5" place="5" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6445" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4460" />
                    <RANKING order="2" place="2" resultid="4045" />
                    <RANKING order="3" place="3" resultid="3094" />
                    <RANKING order="4" place="4" resultid="3139" />
                    <RANKING order="5" place="-1" resultid="4725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6446" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4355" />
                    <RANKING order="2" place="2" resultid="4871" />
                    <RANKING order="3" place="3" resultid="5220" />
                    <RANKING order="4" place="4" resultid="5040" />
                    <RANKING order="5" place="-1" resultid="3307" />
                    <RANKING order="6" place="-1" resultid="3520" />
                    <RANKING order="7" place="-1" resultid="4414" />
                    <RANKING order="8" place="-1" resultid="4626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6447" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4946" />
                    <RANKING order="2" place="2" resultid="5733" />
                    <RANKING order="3" place="3" resultid="4702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6448" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4651" />
                    <RANKING order="2" place="2" resultid="5128" />
                    <RANKING order="3" place="3" resultid="2945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6449" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6450" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3465" />
                    <RANKING order="2" place="2" resultid="3065" />
                    <RANKING order="3" place="3" resultid="5748" />
                    <RANKING order="4" place="-1" resultid="5740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6451" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6452" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6453" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5956" daytime="10:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5957" daytime="10:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5958" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5959" daytime="10:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5960" daytime="10:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5961" daytime="10:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5962" daytime="10:30" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1554" daytime="10:32" gender="F" number="30" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6454" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6455" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3431" />
                    <RANKING order="2" place="2" resultid="3008" />
                    <RANKING order="3" place="3" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6456" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3370" />
                    <RANKING order="2" place="2" resultid="3684" />
                    <RANKING order="3" place="3" resultid="3535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6457" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3663" />
                    <RANKING order="2" place="2" resultid="3178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6458" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3153" />
                    <RANKING order="2" place="2" resultid="5376" />
                    <RANKING order="3" place="3" resultid="3528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6459" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4638" />
                    <RANKING order="2" place="2" resultid="3678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6460" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6461" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6462" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4060" />
                    <RANKING order="2" place="2" resultid="5173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6463" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="6464" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="6465" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6466" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6467" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6468" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6469" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5963" daytime="10:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5964" daytime="10:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1571" daytime="10:38" gender="M" number="31" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6470" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5654" />
                    <RANKING order="2" place="2" resultid="4371" />
                    <RANKING order="3" place="3" resultid="3953" />
                    <RANKING order="4" place="4" resultid="3026" />
                    <RANKING order="5" place="5" resultid="3960" />
                    <RANKING order="6" place="-1" resultid="5649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6471" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4478" />
                    <RANKING order="2" place="2" resultid="4166" />
                    <RANKING order="3" place="3" resultid="2987" />
                    <RANKING order="4" place="4" resultid="5650" />
                    <RANKING order="5" place="5" resultid="3116" />
                    <RANKING order="6" place="-1" resultid="5724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6472" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4210" />
                    <RANKING order="2" place="2" resultid="5355" />
                    <RANKING order="3" place="3" resultid="4439" />
                    <RANKING order="4" place="4" resultid="3846" />
                    <RANKING order="5" place="5" resultid="3946" />
                    <RANKING order="6" place="6" resultid="4129" />
                    <RANKING order="7" place="7" resultid="2734" />
                    <RANKING order="8" place="8" resultid="3981" />
                    <RANKING order="9" place="-1" resultid="4502" />
                    <RANKING order="10" place="-1" resultid="5022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6473" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4537" />
                    <RANKING order="2" place="2" resultid="5413" />
                    <RANKING order="3" place="3" resultid="3967" />
                    <RANKING order="4" place="4" resultid="3988" />
                    <RANKING order="5" place="-1" resultid="4186" />
                    <RANKING order="6" place="-1" resultid="4957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6474" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5524" />
                    <RANKING order="2" place="2" resultid="3703" />
                    <RANKING order="3" place="3" resultid="5455" />
                    <RANKING order="4" place="4" resultid="5233" />
                    <RANKING order="5" place="5" resultid="3396" />
                    <RANKING order="6" place="6" resultid="3183" />
                    <RANKING order="7" place="-1" resultid="3171" />
                    <RANKING order="8" place="-1" resultid="4429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6475" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2856" />
                    <RANKING order="2" place="2" resultid="3549" />
                    <RANKING order="3" place="3" resultid="5101" />
                    <RANKING order="4" place="4" resultid="4820" />
                    <RANKING order="5" place="5" resultid="4293" />
                    <RANKING order="6" place="6" resultid="3561" />
                    <RANKING order="7" place="7" resultid="5554" />
                    <RANKING order="8" place="-1" resultid="5010" />
                    <RANKING order="9" place="-1" resultid="5363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6476" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3556" />
                    <RANKING order="2" place="2" resultid="5238" />
                    <RANKING order="3" place="3" resultid="4975" />
                    <RANKING order="4" place="4" resultid="4386" />
                    <RANKING order="5" place="5" resultid="3384" />
                    <RANKING order="6" place="6" resultid="1668" />
                    <RANKING order="7" place="-1" resultid="4073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6477" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4587" />
                    <RANKING order="2" place="2" resultid="5285" />
                    <RANKING order="3" place="3" resultid="4434" />
                    <RANKING order="4" place="4" resultid="4247" />
                    <RANKING order="5" place="5" resultid="4726" />
                    <RANKING order="6" place="-1" resultid="4046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6478" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3215" />
                    <RANKING order="2" place="2" resultid="4392" />
                    <RANKING order="3" place="3" resultid="4032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6479" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5734" />
                    <RANKING order="2" place="2" resultid="4703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6480" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4039" />
                    <RANKING order="2" place="2" resultid="1681" />
                    <RANKING order="3" place="3" resultid="3058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6481" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6482" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6483" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6484" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6485" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5965" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5966" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5967" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5968" daytime="10:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5969" daytime="10:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5970" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5971" daytime="10:52" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1588" daytime="10:54" gender="F" number="32" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6486" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6487" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4559" />
                    <RANKING order="2" place="2" resultid="4364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6488" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5345" />
                    <RANKING order="2" place="2" resultid="4339" />
                    <RANKING order="3" place="3" resultid="5252" />
                    <RANKING order="4" place="4" resultid="3355" />
                    <RANKING order="5" place="5" resultid="3842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6489" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3934" />
                    <RANKING order="2" place="2" resultid="4396" />
                    <RANKING order="3" place="3" resultid="4708" />
                    <RANKING order="4" place="4" resultid="3727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6490" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3903" />
                    <RANKING order="2" place="2" resultid="5323" />
                    <RANKING order="3" place="3" resultid="5760" />
                    <RANKING order="4" place="4" resultid="3165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6491" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5180" />
                    <RANKING order="2" place="2" resultid="3852" />
                    <RANKING order="3" place="3" resultid="4306" />
                    <RANKING order="4" place="4" resultid="3669" />
                    <RANKING order="5" place="5" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6492" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6493" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3246" />
                    <RANKING order="2" place="2" resultid="4484" />
                    <RANKING order="3" place="-1" resultid="2964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6494" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4324" />
                    <RANKING order="2" place="2" resultid="5166" />
                    <RANKING order="3" place="3" resultid="3892" />
                    <RANKING order="4" place="4" resultid="4113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6495" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6496" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6497" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="6498" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="6499" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6500" agemax="94" agemin="90" name="Kategoria N" />
                <AGEGROUP agegroupid="6501" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5972" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5973" daytime="11:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5974" daytime="11:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5975" daytime="11:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1605" daytime="11:26" gender="M" number="33" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6502" agemax="24" agemin="20" name="Kategoria 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5307" />
                    <RANKING order="2" place="2" resultid="3299" />
                    <RANKING order="3" place="3" resultid="4380" />
                    <RANKING order="4" place="4" resultid="3446" />
                    <RANKING order="5" place="5" resultid="5202" />
                    <RANKING order="6" place="6" resultid="2742" />
                    <RANKING order="7" place="-1" resultid="3223" />
                    <RANKING order="8" place="-1" resultid="4254" />
                    <RANKING order="9" place="-1" resultid="4372" />
                    <RANKING order="10" place="-1" resultid="5655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6503" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4988" />
                    <RANKING order="2" place="2" resultid="4167" />
                    <RANKING order="3" place="3" resultid="4932" />
                    <RANKING order="4" place="4" resultid="5383" />
                    <RANKING order="5" place="-1" resultid="3277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6504" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5356" />
                    <RANKING order="2" place="2" resultid="3572" />
                    <RANKING order="3" place="3" resultid="3242" />
                    <RANKING order="4" place="4" resultid="5111" />
                    <RANKING order="5" place="-1" resultid="5398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6505" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5054" />
                    <RANKING order="2" place="2" resultid="3045" />
                    <RANKING order="3" place="3" resultid="4192" />
                    <RANKING order="4" place="4" resultid="3033" />
                    <RANKING order="5" place="5" resultid="5351" />
                    <RANKING order="6" place="6" resultid="3876" />
                    <RANKING order="7" place="7" resultid="3926" />
                    <RANKING order="8" place="8" resultid="1661" />
                    <RANKING order="9" place="-1" resultid="4279" />
                    <RANKING order="10" place="-1" resultid="4958" />
                    <RANKING order="11" place="-1" resultid="5245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6506" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2807" />
                    <RANKING order="2" place="2" resultid="4228" />
                    <RANKING order="3" place="3" resultid="4488" />
                    <RANKING order="4" place="4" resultid="4688" />
                    <RANKING order="5" place="5" resultid="5048" />
                    <RANKING order="6" place="6" resultid="3636" />
                    <RANKING order="7" place="7" resultid="5107" />
                    <RANKING order="8" place="-1" resultid="2761" />
                    <RANKING order="9" place="-1" resultid="4312" />
                    <RANKING order="10" place="-1" resultid="4997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6507" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4173" />
                    <RANKING order="2" place="2" resultid="4798" />
                    <RANKING order="3" place="3" resultid="4455" />
                    <RANKING order="4" place="4" resultid="5446" />
                    <RANKING order="5" place="5" resultid="4179" />
                    <RANKING order="6" place="6" resultid="3542" />
                    <RANKING order="7" place="7" resultid="4657" />
                    <RANKING order="8" place="-1" resultid="4892" />
                    <RANKING order="9" place="-1" resultid="5117" />
                    <RANKING order="10" place="-1" resultid="5391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6508" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5259" />
                    <RANKING order="2" place="2" resultid="3508" />
                    <RANKING order="3" place="3" resultid="3632" />
                    <RANKING order="4" place="4" resultid="4976" />
                    <RANKING order="5" place="5" resultid="3493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6509" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5028" />
                    <RANKING order="2" place="2" resultid="4793" />
                    <RANKING order="3" place="3" resultid="5289" />
                    <RANKING order="4" place="4" resultid="3095" />
                    <RANKING order="5" place="5" resultid="2871" />
                    <RANKING order="6" place="-1" resultid="2782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6510" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4216" />
                    <RANKING order="2" place="2" resultid="4718" />
                    <RANKING order="3" place="3" resultid="5041" />
                    <RANKING order="4" place="4" resultid="3364" />
                    <RANKING order="5" place="5" resultid="4393" />
                    <RANKING order="6" place="6" resultid="3885" />
                    <RANKING order="7" place="7" resultid="4696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6511" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5149" />
                    <RANKING order="2" place="2" resultid="4516" />
                    <RANKING order="3" place="3" resultid="2768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6512" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4713" />
                    <RANKING order="2" place="2" resultid="5755" />
                    <RANKING order="3" place="3" resultid="2925" />
                    <RANKING order="4" place="4" resultid="2753" />
                    <RANKING order="5" place="-1" resultid="3059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6513" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6514" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5159" />
                    <RANKING order="2" place="2" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6515" agemax="89" agemin="85" name="Kategoria M" />
                <AGEGROUP agegroupid="6516" agemax="94" agemin="90" name="Kategoria N">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6517" agemax="99" agemin="95" name="Kategoria O" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5976" daytime="11:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5977" daytime="11:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5978" daytime="11:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5979" daytime="11:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5980" daytime="12:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5981" daytime="12:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5982" daytime="12:18" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5983" daytime="12:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5984" daytime="12:30" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1622" daytime="12:36" gender="F" number="34" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6532" agemax="-1" agemin="-1" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6533" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL" />
                <AGEGROUP agegroupid="6534" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3451" />
                    <RANKING order="2" place="2" resultid="3915" />
                    <RANKING order="3" place="3" resultid="3739" />
                    <RANKING order="4" place="4" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6535" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3720" />
                    <RANKING order="2" place="2" resultid="5338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6536" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4732" />
                    <RANKING order="2" place="2" resultid="4116" />
                    <RANKING order="3" place="3" resultid="4966" />
                    <RANKING order="4" place="4" resultid="3913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6537" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL" />
                <AGEGROUP agegroupid="6538" agemax="-1" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5197" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5985" daytime="12:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5986" daytime="12:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1646" daytime="12:44" gender="M" number="35" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6539" agemax="-1" agemin="-1" name="Kategoria 0" calculate="TOTAL" />
                <AGEGROUP agegroupid="6540" agemax="119" agemin="100" name="Kategoria A" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6541" agemax="159" agemin="120" name="Kategoria B" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4231" />
                    <RANKING order="2" place="2" resultid="3738" />
                    <RANKING order="3" place="3" resultid="4539" />
                    <RANKING order="4" place="4" resultid="2832" />
                    <RANKING order="5" place="5" resultid="3998" />
                    <RANKING order="6" place="-1" resultid="3079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6542" agemax="199" agemin="160" name="Kategoria C" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5062" />
                    <RANKING order="2" place="2" resultid="4492" />
                    <RANKING order="3" place="3" resultid="5565" />
                    <RANKING order="4" place="4" resultid="3589" />
                    <RANKING order="5" place="5" resultid="5339" />
                    <RANKING order="6" place="6" resultid="4733" />
                    <RANKING order="7" place="7" resultid="3193" />
                    <RANKING order="8" place="8" resultid="3722" />
                    <RANKING order="9" place="9" resultid="5340" />
                    <RANKING order="10" place="10" resultid="5222" />
                    <RANKING order="11" place="11" resultid="3917" />
                    <RANKING order="12" place="-1" resultid="4120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6543" agemax="239" agemin="200" name="Kategoria D" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5063" />
                    <RANKING order="2" place="2" resultid="4493" />
                    <RANKING order="3" place="3" resultid="4968" />
                    <RANKING order="4" place="-1" resultid="4281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6544" agemax="279" agemin="240" name="Kategoria E" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6545" agemax="-1" agemin="280" name="Kategoria F" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5198" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5987" daytime="12:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5988" daytime="12:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5989" daytime="12:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="2971" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Malak" birthdate="1988-01-01" gender="M" nation="POL" swrid="4060740" athleteid="2970">
              <RESULTS>
                <RESULT eventid="1144" points="383" reactiontime="+69" swimtime="00:00:30.59" resultid="2972" heatid="5811" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1265" points="432" swimtime="00:00:59.43" resultid="2973" heatid="5857" lane="9" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="426" reactiontime="+72" swimtime="00:00:26.79" resultid="2974" heatid="5939" lane="1" entrytime="00:00:25.00" />
                <RESULT eventid="1537" points="378" reactiontime="+67" swimtime="00:01:06.81" resultid="2975" heatid="5962" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="2724" name="Ilgaplaukiai">
          <ATHLETES>
            <ATHLETE firstname="Vaidotas" lastname="Gumbis" birthdate="1966-01-01" gender="M" nation="POL" athleteid="2723">
              <RESULTS>
                <RESULT eventid="1212" points="413" reactiontime="+66" swimtime="00:02:13.39" resultid="2725" heatid="5834" lane="7" entrytime="00:02:14.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:02.35" />
                    <SPLIT distance="150" swimtime="00:01:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="432" reactiontime="+67" swimtime="00:00:59.43" resultid="2726" heatid="5856" lane="8" entrytime="00:00:59.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="403" reactiontime="+67" swimtime="00:00:27.29" resultid="2727" heatid="5936" lane="1" entrytime="00:00:26.93" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="4894" name="Uks Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-04-07" gender="M" nation="POL" license="503415700182" swrid="4187282" athleteid="4941">
              <RESULTS>
                <RESULT eventid="1144" points="128" reactiontime="+92" swimtime="00:00:44.04" resultid="4942" heatid="5805" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1178" points="159" reactiontime="+95" swimtime="00:03:22.21" resultid="4943" heatid="5817" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.76" />
                    <SPLIT distance="100" swimtime="00:01:39.43" />
                    <SPLIT distance="150" swimtime="00:02:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="158" reactiontime="+92" swimtime="00:01:31.04" resultid="4944" heatid="5886" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="150" reactiontime="+90" swimtime="00:03:18.71" resultid="4945" heatid="5905" lane="6" entrytime="00:03:19.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                    <SPLIT distance="150" swimtime="00:02:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="146" reactiontime="+92" swimtime="00:01:31.74" resultid="4946" heatid="5959" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Rybak-Starczak" birthdate="1975-01-16" gender="F" nation="POL" license="503415600144" swrid="5439532" athleteid="4921">
              <RESULTS>
                <RESULT eventid="1093" points="320" swimtime="00:01:31.17" resultid="4922" heatid="5787" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="278" reactiontime="+107" swimtime="00:03:06.54" resultid="4923" heatid="5813" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:31.56" />
                    <SPLIT distance="150" swimtime="00:02:23.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="302" swimtime="00:01:24.17" resultid="4924" heatid="5879" lane="7" entrytime="00:01:23.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="308" reactiontime="+108" swimtime="00:03:19.26" resultid="4925" heatid="5944" lane="1" entrytime="00:03:20.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:36.45" />
                    <SPLIT distance="150" swimtime="00:02:28.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Barczyk" birthdate="2001-02-13" gender="F" nation="POL" license="103415600129" swrid="4757023" athleteid="4937">
              <RESULTS>
                <RESULT eventid="1127" points="512" reactiontime="+70" swimtime="00:00:31.98" resultid="4938" heatid="5802" lane="7" entrytime="00:00:32.97" entrycourse="SCM" />
                <RESULT eventid="1316" points="426" reactiontime="+77" swimtime="00:01:15.05" resultid="4939" heatid="5880" lane="1" entrytime="00:01:15.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="444" swimtime="00:00:30.04" resultid="4940" heatid="5916" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Kozanecka" birthdate="2001-06-08" gender="F" nation="POL" license="503415600361" swrid="4749880" athleteid="4910">
              <RESULTS>
                <RESULT eventid="1093" points="487" reactiontime="+74" swimtime="00:01:19.21" resultid="4911" heatid="5784" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="493" reactiontime="+70" swimtime="00:00:36.15" resultid="4912" heatid="5859" lane="4" />
                <RESULT eventid="1316" points="491" reactiontime="+75" swimtime="00:01:11.63" resultid="4913" heatid="5876" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="471" reactiontime="+77" swimtime="00:02:52.90" resultid="4914" heatid="5941" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:02:08.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Radzik" birthdate="1995-05-25" gender="F" nation="POL" license="503415600359" swrid="4229123" athleteid="4895">
              <RESULTS>
                <RESULT eventid="1059" points="436" reactiontime="+73" swimtime="00:00:32.15" resultid="4896" heatid="5766" lane="3" />
                <RESULT eventid="1127" points="471" reactiontime="+69" swimtime="00:00:32.88" resultid="4897" heatid="5798" lane="9" />
                <RESULT eventid="1384" points="464" reactiontime="+60" swimtime="00:02:33.54" resultid="4898" heatid="5901" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="150" swimtime="00:01:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="461" reactiontime="+62" swimtime="00:01:11.04" resultid="4899" heatid="5952" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska-Błachowicz" birthdate="1954-07-13" gender="F" nation="POL" license="503415600184" swrid="5471727" athleteid="4900">
              <RESULTS>
                <RESULT eventid="1059" points="70" reactiontime="+108" swimtime="00:00:58.93" resultid="4901" heatid="5768" lane="9" entrytime="00:00:59.00" />
                <RESULT eventid="1127" points="83" reactiontime="+90" swimtime="00:00:58.47" resultid="4902" heatid="5799" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1451" points="109" reactiontime="+99" swimtime="00:00:47.91" resultid="4903" heatid="5917" lane="5" entrytime="00:00:46.00" />
                <RESULT eventid="1520" points="72" reactiontime="+97" swimtime="00:02:11.89" resultid="4904" heatid="5953" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Masłek" birthdate="1953-01-01" gender="F" nation="POL" athleteid="5399">
              <RESULTS>
                <RESULT eventid="1093" points="105" reactiontime="+135" swimtime="00:02:12.18" resultid="5400" heatid="5786" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" status="DNS" swimtime="00:00:00.00" resultid="5401" heatid="5861" lane="4" entrytime="00:00:56.00" />
                <RESULT eventid="1451" points="93" swimtime="00:00:50.49" resultid="5402" heatid="5917" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1486" points="114" reactiontime="+100" swimtime="00:04:36.91" resultid="5403" heatid="5943" lane="8" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.14" />
                    <SPLIT distance="100" swimtime="00:02:12.85" />
                    <SPLIT distance="150" swimtime="00:03:24.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" license="503415700353" swrid="5471729" athleteid="4947">
              <RESULTS>
                <RESULT eventid="1144" points="176" reactiontime="+87" swimtime="00:00:39.62" resultid="4948" heatid="5806" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1212" points="224" reactiontime="+94" swimtime="00:02:43.55" resultid="4949" heatid="5831" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="267" reactiontime="+93" swimtime="00:01:09.76" resultid="4950" heatid="5851" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="154" reactiontime="+81" swimtime="00:03:16.75" resultid="4951" heatid="5905" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:02:25.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="309" reactiontime="+85" swimtime="00:00:29.79" resultid="4952" heatid="5933" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1537" points="154" reactiontime="+83" swimtime="00:01:30.00" resultid="4953" heatid="5958" lane="4" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Barełkowska" birthdate="1948-08-02" gender="F" nation="POL" license="503415600350" swrid="4920301" athleteid="4915">
              <RESULTS>
                <RESULT eventid="1093" points="69" reactiontime="+115" swimtime="00:02:31.70" resultid="4916" heatid="5786" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="42" reactiontime="+83" swimtime="00:01:13.39" resultid="4917" heatid="5799" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1282" status="DNS" swimtime="00:00:00.00" resultid="4918" heatid="5861" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1451" points="37" reactiontime="+117" swimtime="00:01:08.54" resultid="4919" heatid="5917" lane="3" entrytime="00:00:47.00" />
                <RESULT eventid="1520" points="42" reactiontime="+89" swimtime="00:02:36.79" resultid="4920" heatid="5952" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Szczesiak" birthdate="1955-05-22" gender="M" nation="POL" license="503415700271" athleteid="4959">
              <RESULTS>
                <RESULT eventid="1265" points="204" reactiontime="+121" swimtime="00:01:16.29" resultid="4960" heatid="5849" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="202" reactiontime="+88" swimtime="00:00:34.32" resultid="4961" heatid="5928" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Sęczkowski" birthdate="1995-11-15" gender="M" nation="POL" license="503415700363" athleteid="4926">
              <RESULTS>
                <RESULT eventid="1110" points="480" reactiontime="+65" swimtime="00:01:10.65" resultid="4927" heatid="5795" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="453" reactiontime="+67" swimtime="00:02:09.30" resultid="4928" heatid="5834" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="150" swimtime="00:01:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="492" swimtime="00:00:56.90" resultid="4929" heatid="5857" lane="7" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="452" reactiontime="+63" swimtime="00:01:04.20" resultid="4930" heatid="5891" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="472" reactiontime="+63" swimtime="00:00:25.88" resultid="4931" heatid="5938" lane="2" entrytime="00:00:25.50" />
                <RESULT eventid="1605" points="422" reactiontime="+70" swimtime="00:04:42.94" resultid="4932" heatid="5983" lane="6" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:39.35" />
                    <SPLIT distance="200" swimtime="00:02:15.18" />
                    <SPLIT distance="250" swimtime="00:02:51.87" />
                    <SPLIT distance="300" swimtime="00:03:28.93" />
                    <SPLIT distance="350" swimtime="00:04:06.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Gołembiewski" birthdate="1985-03-14" gender="M" nation="POL" license="503415700164" swrid="4061025" athleteid="4954">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="4955" heatid="5834" lane="3" entrytime="00:02:08.00" />
                <RESULT eventid="1367" status="DNS" swimtime="00:00:00.00" resultid="4956" heatid="5900" lane="9" entrytime="00:02:26.00" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4957" heatid="5970" lane="9" entrytime="00:01:07.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4958" heatid="5983" lane="3" entrytime="00:04:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Orłowski" birthdate="1982-12-11" gender="M" nation="POL" license="503415700360" athleteid="4905">
              <RESULTS>
                <RESULT eventid="1076" points="365" reactiontime="+69" swimtime="00:00:30.43" resultid="4906" heatid="5773" lane="1" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="4907" heatid="5826" lane="5" />
                <RESULT eventid="1265" points="388" reactiontime="+74" swimtime="00:01:01.61" resultid="4908" heatid="5846" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4909" heatid="5924" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Cybertowicz" birthdate="1966-01-12" gender="M" nation="POL" license="503415700177" swrid="4269915" athleteid="4933">
              <RESULTS>
                <RESULT eventid="1110" points="289" reactiontime="+79" swimtime="00:01:23.62" resultid="4934" heatid="5793" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="316" reactiontime="+78" swimtime="00:00:37.04" resultid="4935" heatid="5871" lane="0" entrytime="00:00:37.70" entrycourse="SCM" />
                <RESULT eventid="1503" points="254" swimtime="00:03:09.54" resultid="4936" heatid="5948" lane="9" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:20.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="408" reactiontime="+73" swimtime="00:01:50.20" resultid="4964" heatid="5912" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                    <SPLIT distance="150" swimtime="00:01:22.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4905" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4947" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="4926" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="4954" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" points="217" reactiontime="+85" swimtime="00:02:30.34" resultid="4968" heatid="5987" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:01:56.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4941" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="4933" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="4947" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4959" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1622" points="174" reactiontime="+95" swimtime="00:03:03.14" resultid="4966" heatid="5986" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.46" />
                    <SPLIT distance="100" swimtime="00:01:56.28" />
                    <SPLIT distance="150" swimtime="00:02:28.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4900" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="5399" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4895" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4921" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="145" reactiontime="+86" swimtime="00:03:02.84" resultid="4962" heatid="5837" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.73" />
                    <SPLIT distance="100" swimtime="00:01:48.50" />
                    <SPLIT distance="150" swimtime="00:02:26.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4915" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="4933" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="4921" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4941" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5465" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Fidurski" birthdate="1986-01-01" gender="M" nation="POL" athleteid="5464">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="5466" heatid="5831" lane="2" entrytime="00:02:46.00" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="5467" heatid="5853" lane="8" entrytime="00:01:06.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="5468" heatid="5905" lane="5" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2966" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-01-01" gender="F" nation="POL" athleteid="2965">
              <RESULTS>
                <RESULT eventid="1059" points="176" reactiontime="+117" swimtime="00:00:43.46" resultid="2967" heatid="5768" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1451" points="237" swimtime="00:00:37.05" resultid="2969" heatid="5918" lane="9" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5427" name="Swim2tri">
          <ATHLETES>
            <ATHLETE firstname="Norbert" lastname="Giecewicz" birthdate="1990-03-14" gender="M" nation="POL" athleteid="5432">
              <RESULTS>
                <RESULT eventid="1076" points="365" reactiontime="+86" swimtime="00:00:30.43" resultid="5433" heatid="5781" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1178" points="345" reactiontime="+90" swimtime="00:02:36.29" resultid="5434" heatid="5820" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="388" swimtime="00:01:01.59" resultid="5435" heatid="5855" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Mazur" birthdate="1984-10-05" gender="F" nation="POL" athleteid="5428">
              <RESULTS>
                <RESULT eventid="1093" points="292" reactiontime="+88" swimtime="00:01:33.95" resultid="5429" heatid="5787" lane="3" entrytime="00:01:34.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="321" swimtime="00:00:41.68" resultid="5430" heatid="5863" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1486" points="263" reactiontime="+95" swimtime="00:03:29.93" resultid="5431" heatid="5944" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:37.29" />
                    <SPLIT distance="150" swimtime="00:02:33.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Gągola" birthdate="2000-02-02" gender="F" nation="POL" athleteid="5436">
              <RESULTS>
                <RESULT eventid="1059" points="128" reactiontime="+97" swimtime="00:00:48.28" resultid="5437" heatid="5769" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1282" points="214" reactiontime="+85" swimtime="00:00:47.68" resultid="5438" heatid="5863" lane="0" entrytime="00:00:43.00" />
                <RESULT eventid="1451" points="221" reactiontime="+94" swimtime="00:00:37.87" resultid="5439" heatid="5918" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5420" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Bartniak" birthdate="1997-01-01" gender="F" nation="POL" athleteid="5419">
              <RESULTS>
                <RESULT eventid="1093" points="451" reactiontime="+80" swimtime="00:01:21.30" resultid="5421" heatid="5788" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="446" reactiontime="+81" swimtime="00:02:39.46" resultid="5422" heatid="5814" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:02:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="482" reactiontime="+79" swimtime="00:01:12.05" resultid="5423" heatid="5881" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="440" reactiontime="+81" swimtime="00:02:56.84" resultid="5424" heatid="5944" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                    <SPLIT distance="150" swimtime="00:02:11.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02902" nation="POL" region="02" clubid="4969" name="Uks Czwórka Nakło">
          <ATHLETES>
            <ATHLETE firstname="Radosław" lastname="Staszkiewicz" birthdate="1968-04-21" gender="M" nation="POL" license="102902700326" swrid="5337392" athleteid="4970">
              <RESULTS>
                <RESULT eventid="1076" points="268" reactiontime="+84" swimtime="00:00:33.72" resultid="4971" heatid="5778" lane="3" entrytime="00:00:31.89" />
                <RESULT eventid="1178" points="281" reactiontime="+111" swimtime="00:02:47.36" resultid="4972" heatid="5818" lane="1" entrytime="00:02:49.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                    <SPLIT distance="150" swimtime="00:02:08.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="259" swimtime="00:01:17.30" resultid="4973" heatid="5888" lane="7" entrytime="00:01:17.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="252" reactiontime="+123" swimtime="00:02:51.34" resultid="4974" heatid="5899" lane="2" entrytime="00:02:45.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="288" reactiontime="+96" swimtime="00:01:12.27" resultid="4975" heatid="5968" lane="5" entrytime="00:01:10.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="283" reactiontime="+101" swimtime="00:05:23.01" resultid="4976" heatid="5981" lane="2" entrytime="00:05:23.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="150" swimtime="00:01:53.73" />
                    <SPLIT distance="200" swimtime="00:02:35.28" />
                    <SPLIT distance="250" swimtime="00:03:17.30" />
                    <SPLIT distance="300" swimtime="00:03:59.59" />
                    <SPLIT distance="350" swimtime="00:04:41.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Spychalski" birthdate="1980-09-05" gender="M" nation="POL" license="102902700357" swrid="5337379" athleteid="4977">
              <RESULTS>
                <RESULT eventid="1144" points="183" reactiontime="+88" swimtime="00:00:39.10" resultid="4978" heatid="5806" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1212" points="310" reactiontime="+83" swimtime="00:02:26.81" resultid="4979" heatid="5832" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:47.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3643" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Stoińska" birthdate="1983-01-01" gender="F" nation="POL" athleteid="3642">
              <RESULTS>
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="3644" heatid="5798" lane="7" />
                <RESULT eventid="1384" status="DNS" swimtime="00:00:00.00" resultid="3645" heatid="5901" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5412" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Nowicki" birthdate="1984-01-01" gender="M" nation="POL" athleteid="5411">
              <RESULTS>
                <RESULT eventid="1571" points="222" reactiontime="+95" swimtime="00:01:18.87" resultid="5413" heatid="5965" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="337" reactiontime="+92" swimtime="00:00:31.23" resultid="5414" heatid="5772" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1663" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Łopuszyński" birthdate="1969-01-01" gender="M" nation="POL" athleteid="1662">
              <RESULTS>
                <RESULT eventid="1076" points="105" reactiontime="+105" swimtime="00:00:46.09" resultid="1664" heatid="5774" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1178" points="105" swimtime="00:03:51.83" resultid="1665" heatid="5816" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:53.81" />
                    <SPLIT distance="150" swimtime="00:02:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="97" reactiontime="+121" swimtime="00:03:54.83" resultid="1666" heatid="5897" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:49.55" />
                    <SPLIT distance="150" swimtime="00:02:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="108" reactiontime="+119" swimtime="00:00:42.26" resultid="1667" heatid="5925" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1571" points="90" reactiontime="+105" swimtime="00:01:46.57" resultid="1668" heatid="5966" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2715" name="niezrzeszony" />
        <CLUB type="CLUB" code="03210" nation="POL" region="10" clubid="4540" name="MKP Gdańsk">
          <ATHLETES>
            <ATHLETE firstname="Aleksander" lastname="Weiss" birthdate="1994-08-11" gender="M" nation="POL" license="103210700095" swrid="4104763" athleteid="4541">
              <RESULTS>
                <RESULT eventid="1299" points="589" swimtime="00:00:30.12" resultid="4542" heatid="5865" lane="2" />
                <RESULT eventid="1333" points="502" swimtime="00:01:01.99" resultid="4543" heatid="5883" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="540" reactiontime="+78" swimtime="00:00:24.75" resultid="4544" heatid="5924" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5385" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-01-01" gender="M" nation="POL" athleteid="5384">
              <RESULTS>
                <RESULT eventid="1144" points="163" reactiontime="+103" swimtime="00:00:40.63" resultid="5386" heatid="5804" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1212" points="168" reactiontime="+97" swimtime="00:02:59.88" resultid="5387" heatid="5830" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:19.93" />
                    <SPLIT distance="150" swimtime="00:02:08.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="193" reactiontime="+93" swimtime="00:01:17.70" resultid="5388" heatid="5849" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="139" reactiontime="+93" swimtime="00:01:35.00" resultid="5389" heatid="5884" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5390" heatid="5926" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="5391" heatid="5979" lane="7" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Kubiak" birthdate="1989-01-01" gender="M" nation="POL" athleteid="5392">
              <RESULTS>
                <RESULT eventid="1178" points="155" swimtime="00:03:23.79" resultid="5393" heatid="5816" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                    <SPLIT distance="100" swimtime="00:01:43.98" />
                    <SPLIT distance="150" swimtime="00:02:45.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="248" swimtime="00:02:38.01" resultid="5394" heatid="5831" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:01:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="139" swimtime="00:03:28.77" resultid="5395" heatid="5898" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:40.42" />
                    <SPLIT distance="150" swimtime="00:02:36.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="82" reactiontime="+143" swimtime="00:04:03.05" resultid="5396" heatid="5905" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                    <SPLIT distance="100" swimtime="00:01:58.43" />
                    <SPLIT distance="150" swimtime="00:03:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="5397" heatid="5946" lane="8" entrytime="00:04:00.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="5398" heatid="5980" lane="1" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" clubid="3521" name="Uks Delfin Masters Tarnobrzeg">
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Urbaniak" birthdate="1991-03-03" gender="F" nation="POL" license="500408600214" swrid="4072332" athleteid="3529">
              <RESULTS>
                <RESULT eventid="1059" points="366" reactiontime="+73" swimtime="00:00:34.07" resultid="3530" heatid="5771" lane="9" entrytime="00:00:32.80" />
                <RESULT eventid="1195" points="403" reactiontime="+76" swimtime="00:02:29.39" resultid="3531" heatid="5824" lane="3" entrytime="00:02:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                    <SPLIT distance="150" swimtime="00:01:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="396" swimtime="00:01:08.38" resultid="3532" heatid="5843" lane="9" entrytime="00:01:12.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="255" reactiontime="+79" swimtime="00:03:08.45" resultid="3533" heatid="5895" lane="5" entrytime="00:03:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:16.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="370" reactiontime="+77" swimtime="00:03:07.39" resultid="3534" heatid="5943" lane="4" entrytime="00:03:25.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:30.21" />
                    <SPLIT distance="150" swimtime="00:02:18.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="279" reactiontime="+46" swimtime="00:01:23.57" resultid="3535" heatid="5964" lane="8" entrytime="00:01:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Meksuła" birthdate="1977-03-28" gender="F" nation="POL" license="500408600207" swrid="4992937" athleteid="3577">
              <RESULTS>
                <RESULT eventid="1059" points="261" reactiontime="+77" swimtime="00:00:38.12" resultid="3578" heatid="5769" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1127" points="264" reactiontime="+72" swimtime="00:00:39.89" resultid="3579" heatid="5800" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1247" points="315" reactiontime="+73" swimtime="00:01:13.85" resultid="3580" heatid="5842" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="274" swimtime="00:01:26.94" resultid="3581" heatid="5879" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="333" reactiontime="+78" swimtime="00:00:33.05" resultid="3582" heatid="5919" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1520" status="DNS" swimtime="00:00:00.00" resultid="3583" heatid="5954" lane="9" entrytime="00:01:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelika" lastname="Rozmus" birthdate="1978-03-30" gender="F" nation="POL" license="500408600206" swrid="4992936" athleteid="3522">
              <RESULTS>
                <RESULT eventid="1093" points="296" reactiontime="+83" swimtime="00:01:33.48" resultid="3523" heatid="5787" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="287" reactiontime="+85" swimtime="00:03:04.74" resultid="3524" heatid="5813" lane="4" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:28.81" />
                    <SPLIT distance="150" swimtime="00:02:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="293" swimtime="00:00:43.00" resultid="3525" heatid="5863" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="1316" points="288" reactiontime="+91" swimtime="00:01:25.50" resultid="3526" heatid="5878" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="275" reactiontime="+98" swimtime="00:03:26.87" resultid="3527" heatid="5944" lane="8" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.69" />
                    <SPLIT distance="100" swimtime="00:01:40.66" />
                    <SPLIT distance="150" swimtime="00:02:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="192" reactiontime="+96" swimtime="00:01:34.64" resultid="3528" heatid="5963" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kunicki" birthdate="1972-03-14" gender="M" nation="POL" license="500408700202" swrid="4992901" athleteid="3557">
              <RESULTS>
                <RESULT eventid="1076" points="281" reactiontime="+81" swimtime="00:00:33.20" resultid="3558" heatid="5776" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1178" points="220" reactiontime="+81" swimtime="00:03:01.34" resultid="3559" heatid="5817" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:22.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="174" reactiontime="+96" swimtime="00:03:13.64" resultid="3560" heatid="5898" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:33.86" />
                    <SPLIT distance="150" swimtime="00:02:24.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="220" reactiontime="+84" swimtime="00:01:19.13" resultid="3561" heatid="5967" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Tobiasz" birthdate="1979-02-01" gender="F" nation="POL" license="500408600203" athleteid="3562">
              <RESULTS>
                <RESULT eventid="1059" points="132" reactiontime="+81" swimtime="00:00:47.82" resultid="3563" heatid="5768" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1316" points="146" swimtime="00:01:47.29" resultid="3564" heatid="5877" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3565" heatid="5918" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Zieliński" birthdate="1989-04-27" gender="M" nation="POL" license="500408700239" swrid="4071551" athleteid="3566">
              <RESULTS>
                <RESULT eventid="1110" points="474" reactiontime="+82" swimtime="00:01:10.96" resultid="3567" heatid="5795" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="382" reactiontime="+90" swimtime="00:02:31.03" resultid="3568" heatid="5819" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="475" reactiontime="+77" swimtime="00:00:32.34" resultid="3569" heatid="5874" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1333" points="377" reactiontime="+80" swimtime="00:01:08.20" resultid="3570" heatid="5890" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="439" reactiontime="+85" swimtime="00:02:38.04" resultid="3571" heatid="5948" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="388" swimtime="00:04:50.90" resultid="3572" heatid="5982" lane="7" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:45.84" />
                    <SPLIT distance="200" swimtime="00:02:23.07" />
                    <SPLIT distance="250" swimtime="00:03:00.47" />
                    <SPLIT distance="300" swimtime="00:03:37.62" />
                    <SPLIT distance="350" swimtime="00:04:14.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ślęczka" birthdate="1974-10-23" gender="M" nation="POL" license="500408700205" swrid="4992942" athleteid="3543">
              <RESULTS>
                <RESULT eventid="1076" points="385" reactiontime="+80" swimtime="00:00:29.88" resultid="3544" heatid="5776" lane="9" entrytime="00:00:36.74" />
                <RESULT eventid="1110" points="413" reactiontime="+75" swimtime="00:01:14.26" resultid="3545" heatid="5795" lane="0" entrytime="00:01:16.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="444" reactiontime="+77" swimtime="00:00:58.89" resultid="3546" heatid="5852" lane="0" entrytime="00:01:08.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="371" reactiontime="+70" swimtime="00:01:08.54" resultid="3547" heatid="5890" lane="1" entrytime="00:01:10.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="438" reactiontime="+73" swimtime="00:00:26.53" resultid="3548" heatid="5931" lane="3" entrytime="00:00:30.74" />
                <RESULT eventid="1571" points="337" swimtime="00:01:08.64" resultid="3549" heatid="5968" lane="7" entrytime="00:01:12.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Darowski" birthdate="1971-01-14" gender="M" nation="POL" license="500408700211" swrid="5465834" athleteid="3550">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1110" points="466" reactiontime="+72" swimtime="00:01:11.34" resultid="3551" heatid="5795" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="421" reactiontime="+82" swimtime="00:02:26.24" resultid="3552" heatid="5819" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="455" reactiontime="+68" swimtime="00:00:32.81" resultid="3553" heatid="5873" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1333" points="388" reactiontime="+71" swimtime="00:01:07.51" resultid="3554" heatid="5891" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1503" points="445" reactiontime="+74" swimtime="00:02:37.34" resultid="3555" heatid="5950" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="329" reactiontime="+75" swimtime="00:01:09.16" resultid="3556" heatid="5969" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Janus" birthdate="1987-10-02" gender="F" nation="POL" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1127" points="375" reactiontime="+64" swimtime="00:00:35.47" resultid="3574" heatid="5800" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1316" points="414" reactiontime="+78" swimtime="00:01:15.82" resultid="3575" heatid="5878" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="351" reactiontime="+68" swimtime="00:01:17.78" resultid="3576" heatid="5954" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Płaneta" birthdate="1974-09-12" gender="M" nation="POL" license="500408700210" swrid="4992944" athleteid="3536">
              <RESULTS>
                <RESULT eventid="1144" points="221" reactiontime="+81" swimtime="00:00:36.70" resultid="3537" heatid="5807" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1212" points="279" reactiontime="+76" swimtime="00:02:32.04" resultid="3538" heatid="5832" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="177" reactiontime="+85" swimtime="00:03:12.63" resultid="3539" heatid="5898" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:32.76" />
                    <SPLIT distance="150" swimtime="00:02:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="194" reactiontime="+84" swimtime="00:03:02.25" resultid="3540" heatid="5905" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:18.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="288" reactiontime="+70" swimtime="00:00:30.51" resultid="3541" heatid="5932" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1605" points="266" swimtime="00:05:29.86" resultid="3542" heatid="5980" lane="7" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                    <SPLIT distance="150" swimtime="00:01:58.23" />
                    <SPLIT distance="200" swimtime="00:02:40.13" />
                    <SPLIT distance="250" swimtime="00:03:23.14" />
                    <SPLIT distance="300" swimtime="00:04:06.46" />
                    <SPLIT distance="350" swimtime="00:04:49.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="378" reactiontime="+71" swimtime="00:01:53.10" resultid="3588" heatid="5911" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="100" swimtime="00:00:56.09" />
                    <SPLIT distance="150" swimtime="00:01:26.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3550" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3566" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3557" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3543" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="377" reactiontime="+84" swimtime="00:02:05.18" resultid="3589" heatid="5987" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:06.19" />
                    <SPLIT distance="150" swimtime="00:01:38.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3550" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3566" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3557" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3543" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="360" reactiontime="+81" swimtime="00:02:09.98" resultid="3586" heatid="5909" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:06.56" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3522" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3529" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3573" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3577" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="340" reactiontime="+69" swimtime="00:02:26.57" resultid="3587" heatid="5985" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:17.88" />
                    <SPLIT distance="150" swimtime="00:01:53.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3573" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3522" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3529" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3577" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1229" reactiontime="+65" status="DSQ" swimtime="00:00:00.00" resultid="3584" heatid="5836" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:41.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3573" number="1" reactiontime="+65" status="DSQ" />
                    <RELAYPOSITION athleteid="3566" number="2" reactiontime="-16" status="DSQ" />
                    <RELAYPOSITION athleteid="3529" number="3" reactiontime="+43" status="DSQ" />
                    <RELAYPOSITION athleteid="3543" number="4" reactiontime="+28" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="317" reactiontime="+75" swimtime="00:02:21.00" resultid="3585" heatid="5837" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3577" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3550" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3557" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3522" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5227" name="START Poznań">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Kaczmarek" birthdate="1982-10-03" gender="M" nation="POL" athleteid="5239">
              <RESULTS>
                <RESULT eventid="1110" points="297" reactiontime="+91" swimtime="00:01:22.94" resultid="5240" heatid="5794" lane="9" entrytime="00:01:22.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="345" reactiontime="+89" swimtime="00:01:04.07" resultid="5242" heatid="5854" lane="0" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="235" reactiontime="+94" swimtime="00:02:51.04" resultid="5243" heatid="5906" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:23.42" />
                    <SPLIT distance="150" swimtime="00:02:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="286" swimtime="00:03:02.28" resultid="5244" heatid="5949" lane="7" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="150" swimtime="00:02:14.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="5245" heatid="5980" lane="4" entrytime="00:05:30.00" entrycourse="SCM" />
                <RESULT eventid="1178" points="263" reactiontime="+102" swimtime="00:02:51.02" resultid="5720" heatid="5817" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:09.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Parysek" birthdate="1977-12-17" gender="M" nation="POL" athleteid="5228">
              <RESULTS>
                <RESULT eventid="1076" points="327" reactiontime="+75" swimtime="00:00:31.56" resultid="5229" heatid="5779" lane="9" entrytime="00:00:31.13" entrycourse="SCM" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="5230" heatid="5853" lane="0" entrytime="00:01:06.11" entrycourse="SCM" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5231" heatid="5889" lane="8" entrytime="00:01:13.41" entrycourse="SCM" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5232" heatid="5933" lane="9" entrytime="00:00:29.03" entrycourse="SCM" />
                <RESULT eventid="1571" points="279" reactiontime="+78" swimtime="00:01:13.10" resultid="5233" heatid="5967" lane="2" entrytime="00:01:16.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Wróbel" birthdate="1967-02-06" gender="M" nation="POL" athleteid="5234">
              <RESULTS>
                <RESULT eventid="1076" points="400" reactiontime="+76" swimtime="00:00:29.50" resultid="5235" heatid="5779" lane="5" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1178" points="333" swimtime="00:02:38.07" resultid="5236" heatid="5819" lane="2" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:59.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="338" reactiontime="+85" swimtime="00:01:10.74" resultid="5237" heatid="5890" lane="6" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="313" reactiontime="+85" swimtime="00:01:10.30" resultid="5238" heatid="5968" lane="6" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Kostencka" birthdate="1987-03-06" gender="F" nation="POL" athleteid="5246">
              <RESULTS>
                <RESULT eventid="1127" points="377" reactiontime="+73" swimtime="00:00:35.43" resultid="5247" heatid="5801" lane="2" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1195" points="373" reactiontime="+83" swimtime="00:02:33.33" resultid="5248" heatid="5825" lane="9" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="369" reactiontime="+81" swimtime="00:01:10.03" resultid="5249" heatid="5843" lane="7" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="362" reactiontime="+82" swimtime="00:02:46.77" resultid="5250" heatid="5903" lane="2" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="150" swimtime="00:02:03.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="371" reactiontime="+77" swimtime="00:01:16.38" resultid="5251" heatid="5954" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="352" reactiontime="+82" swimtime="00:05:31.25" resultid="5252" heatid="5974" lane="4" entrytime="00:05:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:00.32" />
                    <SPLIT distance="200" swimtime="00:02:42.29" />
                    <SPLIT distance="250" swimtime="00:03:24.84" />
                    <SPLIT distance="300" swimtime="00:04:07.11" />
                    <SPLIT distance="350" swimtime="00:04:49.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Dmytrów" birthdate="1961-07-15" gender="M" nation="POL" athleteid="5260">
              <RESULTS>
                <RESULT eventid="1110" points="311" reactiontime="+78" swimtime="00:01:21.65" resultid="5261" heatid="5793" lane="6" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="329" reactiontime="+73" swimtime="00:00:36.55" resultid="5262" heatid="5870" lane="0" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1503" points="280" reactiontime="+80" swimtime="00:03:03.49" resultid="5263" heatid="5947" lane="6" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:16.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Monczak" birthdate="1967-11-03" gender="M" nation="POL" athleteid="5253">
              <RESULTS>
                <RESULT eventid="1178" points="351" reactiontime="+85" swimtime="00:02:35.35" resultid="5254" heatid="5816" lane="6" entrytime="00:03:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="422" reactiontime="+60" swimtime="00:02:12.44" resultid="5255" heatid="5834" lane="2" entrytime="00:02:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="416" reactiontime="+72" swimtime="00:01:00.19" resultid="5256" heatid="5856" lane="1" entrytime="00:00:59.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="336" reactiontime="+74" swimtime="00:01:10.84" resultid="5257" heatid="5891" lane="9" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="388" reactiontime="+70" swimtime="00:00:27.64" resultid="5258" heatid="5935" lane="2" entrytime="00:00:27.03" entrycourse="SCM" />
                <RESULT eventid="1605" points="394" reactiontime="+77" swimtime="00:04:49.49" resultid="5259" heatid="5982" lane="4" entrytime="00:04:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:08.66" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                    <SPLIT distance="200" swimtime="00:02:23.03" />
                    <SPLIT distance="250" swimtime="00:03:00.30" />
                    <SPLIT distance="300" swimtime="00:03:37.76" />
                    <SPLIT distance="350" swimtime="00:04:14.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3283" name="Delfin Masters Łódź">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Gaede" birthdate="1974-01-24" gender="M" nation="POL" athleteid="3288">
              <RESULTS>
                <RESULT eventid="1110" points="239" reactiontime="+88" swimtime="00:01:29.09" resultid="3289" heatid="5792" lane="8" entrytime="00:01:32.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="262" swimtime="00:00:39.45" resultid="3290" heatid="5870" lane="7" entrytime="00:00:38.69" />
                <RESULT eventid="1503" points="237" reactiontime="+83" swimtime="00:03:13.99" resultid="3291" heatid="5947" lane="5" entrytime="00:03:11.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:32.61" />
                    <SPLIT distance="150" swimtime="00:02:23.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Kadłubiec" birthdate="1971-02-25" gender="M" nation="POL" athleteid="3284">
              <RESULTS>
                <RESULT eventid="1110" points="277" reactiontime="+87" swimtime="00:01:24.89" resultid="3285" heatid="5792" lane="5" entrytime="00:01:28.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="277" reactiontime="+86" swimtime="00:00:38.70" resultid="3286" heatid="5869" lane="5" entrytime="00:00:39.25" />
                <RESULT eventid="1503" points="280" swimtime="00:03:03.56" resultid="3287" heatid="5948" lane="7" entrytime="00:03:05.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:02:14.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5123" name="Weteran  Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Włodzimierz" lastname="Bosowski" birthdate="1948-05-22" gender="M" nation="POL" license="102611700014" athleteid="5181">
              <RESULTS>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5182" heatid="5925" lane="2" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Kosiak" birthdate="1940-04-20" gender="M" nation="POL" license="102611700027" athleteid="5155">
              <RESULTS>
                <RESULT eventid="1212" points="71" reactiontime="+114" swimtime="00:03:58.91" resultid="5156" heatid="5828" lane="6" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.12" />
                    <SPLIT distance="100" swimtime="00:01:59.65" />
                    <SPLIT distance="150" swimtime="00:03:03.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="80" swimtime="00:01:44.12" resultid="5157" heatid="5848" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="100" reactiontime="+127" swimtime="00:00:43.37" resultid="5158" heatid="5925" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1605" points="70" reactiontime="+142" swimtime="00:08:34.23" resultid="5159" heatid="5977" lane="5" entrytime="00:08:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.64" />
                    <SPLIT distance="100" swimtime="00:02:05.43" />
                    <SPLIT distance="150" swimtime="00:03:12.33" />
                    <SPLIT distance="200" swimtime="00:04:18.23" />
                    <SPLIT distance="250" swimtime="00:05:24.78" />
                    <SPLIT distance="300" swimtime="00:06:29.52" />
                    <SPLIT distance="350" swimtime="00:07:32.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystyna" lastname="Fecica" birthdate="1943-03-12" gender="F" nation="POL" license="102611600019" athleteid="5133">
              <RESULTS>
                <RESULT eventid="1059" points="98" swimtime="00:00:52.82" resultid="5134" heatid="5768" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="1093" points="129" swimtime="00:02:03.19" resultid="5135" heatid="5786" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="131" reactiontime="+89" swimtime="00:00:56.12" resultid="5136" heatid="5862" lane="0" entrytime="00:00:53.00" />
                <RESULT eventid="1486" points="119" reactiontime="+107" swimtime="00:04:33.09" resultid="5137" heatid="5942" lane="4" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.91" />
                    <SPLIT distance="100" swimtime="00:02:08.51" />
                    <SPLIT distance="150" swimtime="00:03:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="79" swimtime="00:02:06.79" resultid="5138" heatid="5963" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Kiszczak" birthdate="1950-02-18" gender="F" nation="POL" license="102611600039" athleteid="5183">
              <RESULTS>
                <RESULT eventid="1059" points="143" reactiontime="+81" swimtime="00:00:46.56" resultid="5184" heatid="5767" lane="6" />
                <RESULT eventid="1127" points="197" reactiontime="+80" swimtime="00:00:43.94" resultid="5185" heatid="5797" lane="3" />
                <RESULT eventid="1316" points="162" reactiontime="+83" swimtime="00:01:43.52" resultid="5186" heatid="5875" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1520" points="190" reactiontime="+79" swimtime="00:01:35.41" resultid="5187" heatid="5951" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" license="102611700032" athleteid="5124">
              <RESULTS>
                <RESULT eventid="1076" points="124" reactiontime="+75" swimtime="00:00:43.52" resultid="5125" heatid="5774" lane="9" entrytime="00:00:45.75" />
                <RESULT eventid="1144" points="115" reactiontime="+74" swimtime="00:00:45.67" resultid="5126" heatid="5805" lane="0" entrytime="00:00:44.80" />
                <RESULT eventid="1401" points="100" reactiontime="+70" swimtime="00:03:47.51" resultid="5127" heatid="5905" lane="8" entrytime="00:03:48.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.64" />
                    <SPLIT distance="100" swimtime="00:01:48.92" />
                    <SPLIT distance="150" swimtime="00:02:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="110" reactiontime="+78" swimtime="00:01:40.71" resultid="5128" heatid="5958" lane="7" entrytime="00:01:46.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" license="102611600029" athleteid="5150">
              <RESULTS>
                <RESULT eventid="1127" points="71" reactiontime="+73" swimtime="00:01:01.74" resultid="5151" heatid="5799" lane="0" entrytime="00:01:00.00" />
                <RESULT eventid="1247" points="72" swimtime="00:02:00.59" resultid="5152" heatid="5841" lane="0" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="68" reactiontime="+67" swimtime="00:02:14.16" resultid="5154" heatid="5952" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="80" swimtime="00:00:53.06" resultid="5425" heatid="5917" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Dąbrowska" birthdate="1958-02-05" gender="F" nation="POL" license="102611600028" athleteid="5167">
              <RESULTS>
                <RESULT eventid="1059" points="79" reactiontime="+88" swimtime="00:00:56.63" resultid="5168" heatid="5767" lane="0" />
                <RESULT eventid="1093" points="138" reactiontime="+87" swimtime="00:02:00.51" resultid="5169" heatid="5785" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="133" reactiontime="+90" swimtime="00:00:55.88" resultid="5170" heatid="5860" lane="8" />
                <RESULT eventid="1316" points="92" reactiontime="+92" swimtime="00:02:05.07" resultid="5171" heatid="5876" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="117" reactiontime="+92" swimtime="00:04:34.51" resultid="5172" heatid="5941" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                    <SPLIT distance="100" swimtime="00:02:11.65" />
                    <SPLIT distance="150" swimtime="00:03:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="63" reactiontime="+84" swimtime="00:02:16.83" resultid="5173" heatid="5963" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" license="502611700035" athleteid="5143">
              <RESULTS>
                <RESULT eventid="1144" points="138" reactiontime="+77" swimtime="00:00:42.93" resultid="5144" heatid="5805" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="179" reactiontime="+96" swimtime="00:02:56.01" resultid="5145" heatid="5828" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="196" reactiontime="+90" swimtime="00:01:17.32" resultid="5146" heatid="5850" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="149" reactiontime="+105" swimtime="00:01:32.77" resultid="5147" heatid="5885" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="173" swimtime="00:00:36.13" resultid="5148" heatid="5928" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1605" points="176" swimtime="00:06:18.66" resultid="5149" heatid="5979" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:02:13.74" />
                    <SPLIT distance="200" swimtime="00:03:02.46" />
                    <SPLIT distance="250" swimtime="00:03:51.78" />
                    <SPLIT distance="300" swimtime="00:04:41.12" />
                    <SPLIT distance="350" swimtime="00:05:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Zagała" birthdate="1959-06-24" gender="F" nation="POL" license="102611600043" athleteid="5160">
              <RESULTS>
                <RESULT eventid="1127" points="163" reactiontime="+74" swimtime="00:00:46.79" resultid="5161" heatid="5799" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1195" points="198" reactiontime="+79" swimtime="00:03:09.43" resultid="5162" heatid="5822" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="188" swimtime="00:00:49.81" resultid="5163" heatid="5861" lane="7" entrytime="00:01:00.00" />
                <RESULT eventid="1384" points="142" reactiontime="+81" swimtime="00:03:47.90" resultid="5164" heatid="5902" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.84" />
                    <SPLIT distance="100" swimtime="00:01:54.54" />
                    <SPLIT distance="150" swimtime="00:02:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="147" reactiontime="+77" swimtime="00:01:44.00" resultid="5165" heatid="5953" lane="8" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="185" reactiontime="+78" swimtime="00:06:50.00" resultid="5166" heatid="5973" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                    <SPLIT distance="150" swimtime="00:02:31.90" />
                    <SPLIT distance="200" swimtime="00:03:24.75" />
                    <SPLIT distance="250" swimtime="00:04:18.06" />
                    <SPLIT distance="300" swimtime="00:05:10.90" />
                    <SPLIT distance="350" swimtime="00:06:02.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" license="102611700015" athleteid="5139">
              <RESULTS>
                <RESULT eventid="1076" points="190" reactiontime="+90" swimtime="00:00:37.82" resultid="5140" heatid="5775" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1333" points="121" swimtime="00:01:39.48" resultid="5141" heatid="5886" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="247" reactiontime="+92" swimtime="00:00:32.10" resultid="5142" heatid="5929" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-18" gender="F" nation="POL" license="102611600033" athleteid="5188">
              <RESULTS>
                <RESULT eventid="1093" points="74" reactiontime="+104" swimtime="00:02:28.28" resultid="5189" heatid="5785" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="63" reactiontime="+77" swimtime="00:01:04.04" resultid="5190" heatid="5798" lane="5" entrytime="00:01:06.00" />
                <RESULT eventid="1282" points="95" swimtime="00:01:02.57" resultid="5191" heatid="5861" lane="9" entrytime="00:01:05.00" />
                <RESULT eventid="1316" points="68" swimtime="00:02:17.85" resultid="5192" heatid="5876" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="74" swimtime="00:05:19.64" resultid="5193" heatid="5942" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.64" />
                    <SPLIT distance="100" swimtime="00:02:35.57" />
                    <SPLIT distance="150" swimtime="00:04:00.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" license="102611600016" athleteid="5174">
              <RESULTS>
                <RESULT eventid="1093" points="386" reactiontime="+86" swimtime="00:01:25.63" resultid="5175" heatid="5788" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="385" reactiontime="+74" swimtime="00:02:31.76" resultid="5176" heatid="5825" lane="8" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="367" reactiontime="+77" swimtime="00:01:10.18" resultid="5177" heatid="5843" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="370" swimtime="00:00:39.78" resultid="5178" heatid="5864" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1486" points="376" reactiontime="+92" swimtime="00:03:06.39" resultid="5179" heatid="5941" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:30.73" />
                    <SPLIT distance="150" swimtime="00:02:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="384" reactiontime="+74" swimtime="00:05:21.72" resultid="5180" heatid="5975" lane="2" entrytime="00:05:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:56.45" />
                    <SPLIT distance="200" swimtime="00:02:37.60" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:04:00.14" />
                    <SPLIT distance="350" swimtime="00:04:41.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Fecica" birthdate="1940-11-29" gender="M" nation="POL" license="102611700018" athleteid="5129">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1110" points="137" reactiontime="+92" swimtime="00:01:47.14" resultid="5130" heatid="5790" lane="4" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="136" reactiontime="+99" swimtime="00:00:49.04" resultid="5131" heatid="5867" lane="3" entrytime="00:00:49.00" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1503" points="129" reactiontime="+112" swimtime="00:03:57.26" resultid="5132" heatid="5946" lane="6" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:54.45" />
                    <SPLIT distance="150" swimtime="00:02:56.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1442" points="148" reactiontime="+109" swimtime="00:02:34.52" resultid="5196" heatid="5911" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5143" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="5155" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="5124" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5139" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1646" points="151" reactiontime="+73" swimtime="00:02:49.52" resultid="5198" heatid="5987" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:35.05" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5124" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5129" number="2" />
                    <RELAYPOSITION athleteid="5139" number="3" />
                    <RELAYPOSITION athleteid="5143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1418" points="119" reactiontime="+92" swimtime="00:03:07.57" resultid="5195" heatid="5909" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.92" />
                    <SPLIT distance="100" swimtime="00:01:44.82" />
                    <SPLIT distance="150" swimtime="00:02:24.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5133" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="5150" number="2" />
                    <RELAYPOSITION athleteid="5160" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="5183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1622" points="113" reactiontime="+71" swimtime="00:03:31.20" resultid="5197" heatid="5985" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:40.59" />
                    <SPLIT distance="150" swimtime="00:02:38.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5183" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5133" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5167" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="5150" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="170" reactiontime="+85" swimtime="00:02:53.48" resultid="5194" heatid="5836" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:02:14.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5183" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5129" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="5139" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5160" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3270" name="Baza Pływania Mysłowice">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Czwartosz" birthdate="1993-04-15" gender="M" nation="POL" swrid="4086584" athleteid="3278">
              <RESULTS>
                <RESULT eventid="1076" points="477" reactiontime="+76" swimtime="00:00:27.83" resultid="3279" heatid="5782" lane="5" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1178" points="371" swimtime="00:02:32.55" resultid="3280" heatid="5820" lane="9" entrytime="00:02:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:06.06" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3281" heatid="5893" lane="9" entrytime="00:01:02.00" entrycourse="SCM" />
                <RESULT eventid="1469" points="481" swimtime="00:00:25.72" resultid="3282" heatid="5939" lane="7" entrytime="00:00:25.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kisiel" birthdate="1993-03-26" gender="M" nation="POL" swrid="4086753" athleteid="3271">
              <RESULTS>
                <RESULT eventid="1076" points="489" reactiontime="+67" swimtime="00:00:27.60" resultid="3272" heatid="5781" lane="6" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1144" points="372" reactiontime="+71" swimtime="00:00:30.87" resultid="3273" heatid="5811" lane="0" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1299" points="343" reactiontime="+73" swimtime="00:00:36.07" resultid="3274" heatid="5873" lane="6" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1401" points="384" reactiontime="+70" swimtime="00:02:25.21" resultid="3275" heatid="5908" lane="8" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="411" reactiontime="+69" swimtime="00:01:04.99" resultid="3276" heatid="5962" lane="5" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="3277" heatid="5983" lane="8" entrytime="00:04:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5119" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michael" lastname="Oleasz" birthdate="1991-01-01" gender="M" nation="POL" athleteid="5118">
              <RESULTS>
                <RESULT eventid="1144" points="472" reactiontime="+55" swimtime="00:00:28.53" resultid="5120" heatid="5811" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1333" points="476" reactiontime="+65" swimtime="00:01:03.10" resultid="5121" heatid="5891" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="482" reactiontime="+60" swimtime="00:01:01.63" resultid="5122" heatid="5962" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3321" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Patryk" lastname="Matysiak" birthdate="1982-01-01" gender="M" nation="POL" athleteid="3320">
              <RESULTS>
                <RESULT eventid="1110" points="234" reactiontime="+74" swimtime="00:01:29.73" resultid="3322" heatid="5792" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="202" reactiontime="+74" swimtime="00:01:23.93" resultid="3323" heatid="5885" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PWR" nation="POL" clubid="2946" name="Masters Politechnika Wrocławska">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Bajor-Traczyńska" birthdate="1977-07-08" gender="F" nation="POL" athleteid="2947">
              <RESULTS>
                <RESULT eventid="1127" points="321" reactiontime="+85" swimtime="00:00:37.36" resultid="2948" heatid="5801" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1195" points="307" reactiontime="+89" swimtime="00:02:43.54" resultid="2949" heatid="5824" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="354" reactiontime="+89" swimtime="00:01:11.02" resultid="2950" heatid="5843" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="2951" heatid="5921" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1520" status="DNS" swimtime="00:00:00.00" resultid="2952" heatid="5954" lane="6" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Kasprzak" birthdate="1979-01-29" gender="F" nation="POL" athleteid="2953">
              <RESULTS>
                <RESULT eventid="1059" points="228" reactiontime="+84" swimtime="00:00:39.85" resultid="2954" heatid="5770" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1127" points="209" reactiontime="+84" swimtime="00:00:43.08" resultid="2955" heatid="5800" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1247" points="292" reactiontime="+88" swimtime="00:01:15.74" resultid="2956" heatid="5842" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="300" reactiontime="+84" swimtime="00:00:34.25" resultid="2957" heatid="5920" lane="4" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Bogdan" birthdate="1966-10-30" gender="F" nation="POL" athleteid="2958">
              <RESULTS>
                <RESULT eventid="1127" points="168" reactiontime="+80" swimtime="00:00:46.37" resultid="2959" heatid="5800" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="2960" heatid="5823" lane="6" entrytime="00:03:00.00" />
                <RESULT eventid="1282" points="166" reactiontime="+105" swimtime="00:00:51.88" resultid="2961" heatid="5863" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1384" points="171" reactiontime="+89" swimtime="00:03:34.17" resultid="2962" heatid="5902" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.89" />
                    <SPLIT distance="100" swimtime="00:01:43.73" />
                    <SPLIT distance="150" swimtime="00:02:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="179" swimtime="00:03:58.62" resultid="2963" heatid="5944" lane="9" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                    <SPLIT distance="100" swimtime="00:01:53.61" />
                    <SPLIT distance="150" swimtime="00:02:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" status="DNS" swimtime="00:00:00.00" resultid="2964" heatid="5974" lane="0" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MMS" nation="POL" clubid="3939" name="Max Masters Szamotuły">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Sędrowicz" birthdate="1997-05-19" gender="M" nation="POL" swrid="4878673" athleteid="3954">
              <RESULTS>
                <RESULT eventid="1110" points="337" reactiontime="+72" swimtime="00:01:19.46" resultid="3955" heatid="5793" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="239" reactiontime="+72" swimtime="00:02:56.44" resultid="3956" heatid="5817" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="373" reactiontime="+68" swimtime="00:00:35.07" resultid="3957" heatid="5872" lane="8" entrytime="00:00:35.60" />
                <RESULT eventid="1333" points="283" reactiontime="+71" swimtime="00:01:15.02" resultid="3958" heatid="5888" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="305" reactiontime="+74" swimtime="00:02:58.49" resultid="3959" heatid="5947" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="210" reactiontime="+76" swimtime="00:01:20.35" resultid="3960" heatid="5967" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Błauciak" birthdate="1982-12-17" gender="M" nation="POL" athleteid="3961">
              <RESULTS>
                <RESULT eventid="1076" points="238" swimtime="00:00:35.07" resultid="3962" heatid="5776" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1178" points="204" reactiontime="+91" swimtime="00:03:06.12" resultid="3963" heatid="5817" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:27.86" />
                    <SPLIT distance="150" swimtime="00:02:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="314" reactiontime="+83" swimtime="00:00:37.13" resultid="3964" heatid="5869" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1333" points="220" reactiontime="+79" swimtime="00:01:21.53" resultid="3965" heatid="5887" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="299" reactiontime="+79" swimtime="00:00:30.13" resultid="3966" heatid="5931" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1571" points="157" reactiontime="+80" swimtime="00:01:28.51" resultid="3967" heatid="5966" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Powąska" birthdate="1990-07-26" gender="M" nation="POL" swrid="4752833" athleteid="3975">
              <RESULTS>
                <RESULT eventid="1076" points="365" reactiontime="+64" swimtime="00:00:30.43" resultid="3976" heatid="5780" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="1144" points="250" reactiontime="+67" swimtime="00:00:35.24" resultid="3977" heatid="5808" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1265" points="347" reactiontime="+52" swimtime="00:01:03.94" resultid="3978" heatid="5855" lane="5" entrytime="00:00:59.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="283" reactiontime="+70" swimtime="00:00:38.45" resultid="3979" heatid="5871" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1469" points="341" reactiontime="+67" swimtime="00:00:28.85" resultid="3980" heatid="5935" lane="1" entrytime="00:00:27.14" />
                <RESULT eventid="1571" points="247" reactiontime="+73" swimtime="00:01:16.05" resultid="3981" heatid="5969" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Cegielski" birthdate="1989-01-23" gender="M" nation="POL" athleteid="3989">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3990" heatid="5773" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3991" heatid="5805" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1265" points="210" reactiontime="+70" swimtime="00:01:15.59" resultid="3992" heatid="5848" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3993" heatid="5883" lane="3" entrytime="00:01:50.00" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="3994" heatid="5926" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="3995" heatid="5958" lane="6" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Pernak" birthdate="1990-11-06" gender="M" nation="POL" athleteid="3968">
              <RESULTS>
                <RESULT eventid="1076" points="175" reactiontime="+96" swimtime="00:00:38.83" resultid="3969" heatid="5774" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1144" points="98" reactiontime="+88" swimtime="00:00:48.16" resultid="3970" heatid="5806" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1265" points="174" swimtime="00:01:20.39" resultid="3971" heatid="5849" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3972" heatid="5884" lane="8" entrytime="00:01:45.00" />
                <RESULT eventid="1469" points="193" reactiontime="+90" swimtime="00:00:34.88" resultid="3973" heatid="5927" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="3974" heatid="5958" lane="8" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szmania" birthdate="1984-12-17" gender="M" nation="POL" athleteid="3982">
              <RESULTS>
                <RESULT eventid="1076" points="152" reactiontime="+80" swimtime="00:00:40.73" resultid="3983" heatid="5775" lane="5" entrytime="00:00:38.00" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1110" reactiontime="+79" status="DSQ" swimtime="00:00:00.00" resultid="3984" heatid="5793" lane="9" entrytime="00:01:28.00" />
                <RESULT eventid="1299" points="207" reactiontime="+80" swimtime="00:00:42.64" resultid="3985" heatid="5870" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1333" points="141" reactiontime="+75" swimtime="00:01:34.64" resultid="3986" heatid="5885" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="187" reactiontime="+77" swimtime="00:00:35.20" resultid="3987" heatid="5929" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1571" points="100" swimtime="00:01:42.79" resultid="3988" heatid="5966" lane="7" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Bartkowiak" birthdate="1988-01-25" gender="M" nation="POL" athleteid="3940">
              <RESULTS>
                <RESULT eventid="1076" points="393" reactiontime="+80" swimtime="00:00:29.69" resultid="3941" heatid="5780" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1144" points="322" reactiontime="+70" swimtime="00:00:32.41" resultid="3942" heatid="5810" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1265" points="381" reactiontime="+83" swimtime="00:01:01.96" resultid="3943" heatid="5855" lane="3" entrytime="00:00:59.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="326" reactiontime="+78" swimtime="00:01:11.53" resultid="3944" heatid="5891" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="378" reactiontime="+75" swimtime="00:00:27.86" resultid="3945" heatid="5935" lane="8" entrytime="00:00:27.14" />
                <RESULT eventid="1571" points="334" reactiontime="+72" swimtime="00:01:08.85" resultid="3946" heatid="5968" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Zajas" birthdate="1999-06-16" gender="M" nation="POL" swrid="4943288" athleteid="3947">
              <RESULTS>
                <RESULT eventid="1076" points="413" swimtime="00:00:29.19" resultid="3948" heatid="5780" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1144" points="359" reactiontime="+100" swimtime="00:00:31.24" resultid="3949" heatid="5810" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1265" points="415" reactiontime="+86" swimtime="00:01:00.22" resultid="3950" heatid="5855" lane="6" entrytime="00:00:59.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="357" reactiontime="+86" swimtime="00:01:09.45" resultid="3951" heatid="5891" lane="0" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="447" swimtime="00:00:26.35" resultid="3952" heatid="5936" lane="7" entrytime="00:00:26.92" />
                <RESULT eventid="1571" points="338" swimtime="00:01:08.57" resultid="3953" heatid="5969" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="311" reactiontime="+71" swimtime="00:02:00.65" resultid="3996" heatid="5912" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:00:56.32" />
                    <SPLIT distance="150" swimtime="00:01:30.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3975" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3940" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3982" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3961" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" points="342" reactiontime="+88" swimtime="00:02:09.28" resultid="3997" heatid="5987" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="150" swimtime="00:01:35.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3947" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3954" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3989" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3968" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1442" points="282" reactiontime="+87" swimtime="00:02:04.71" resultid="5765" heatid="5912" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.97" />
                    <SPLIT distance="100" swimtime="00:00:57.00" />
                    <SPLIT distance="150" swimtime="00:01:30.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3947" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3954" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="3989" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3968" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1646" points="286" reactiontime="+66" swimtime="00:02:17.23" resultid="3998" heatid="5988" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:42.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3940" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3961" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3975" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="3982" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03114" nation="POL" region="14" clubid="4880" name="Uks ,,Pingwiny&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Artur" lastname="Kostanowicz" birthdate="1998-04-03" gender="M" nation="POL" license="103114700307" swrid="4363163" athleteid="4881">
              <RESULTS>
                <RESULT eventid="1076" points="560" reactiontime="+78" swimtime="00:00:26.38" resultid="4882" heatid="5773" lane="9" />
                <RESULT eventid="1144" points="580" reactiontime="+62" swimtime="00:00:26.63" resultid="4883" heatid="5811" lane="5" entrytime="00:00:26.45" entrycourse="SCM" />
                <RESULT eventid="1401" points="498" reactiontime="+68" swimtime="00:02:13.20" resultid="4884" heatid="5908" lane="4" entrytime="00:02:05.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="553" reactiontime="+74" swimtime="00:00:24.56" resultid="4885" heatid="5940" lane="1" entrytime="00:00:24.15" entrycourse="SCM" />
                <RESULT eventid="1537" points="569" reactiontime="+65" swimtime="00:00:58.30" resultid="4886" heatid="5962" lane="4" entrytime="00:00:56.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3010" name="Najmowicz Triatlon Team Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Chodyna" birthdate="1967-01-01" gender="M" nation="POL" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1144" points="212" reactiontime="+75" swimtime="00:00:37.25" resultid="3011" heatid="5810" lane="9" entrytime="00:00:31.50" />
                <RESULT eventid="1469" points="352" reactiontime="+61" swimtime="00:00:28.53" resultid="3012" heatid="5936" lane="8" entrytime="00:00:26.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07414" nation="POL" region="14" clubid="4982" name="UKS Manta Warszawa Włochy">
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" license="507414700150" swrid="4806379" athleteid="4983">
              <RESULTS>
                <RESULT eventid="1110" points="586" reactiontime="+71" swimtime="00:01:06.11" resultid="4984" heatid="5796" lane="7" entrytime="00:01:05.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="581" swimtime="00:00:30.26" resultid="4985" heatid="5874" lane="7" entrytime="00:00:30.20" entrycourse="SCM" />
                <RESULT eventid="1367" points="534" reactiontime="+71" swimtime="00:02:13.34" resultid="4986" heatid="5900" lane="6" entrytime="00:02:15.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:02.90" />
                    <SPLIT distance="150" swimtime="00:01:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="570" reactiontime="+70" swimtime="00:02:24.88" resultid="4987" heatid="5950" lane="4" entrytime="00:02:21.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:47.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="598" reactiontime="+69" swimtime="00:04:11.93" resultid="4988" heatid="5984" lane="6" entrytime="00:04:18.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:33.84" />
                    <SPLIT distance="200" swimtime="00:02:06.13" />
                    <SPLIT distance="250" swimtime="00:02:38.18" />
                    <SPLIT distance="300" swimtime="00:03:10.09" />
                    <SPLIT distance="350" swimtime="00:03:41.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="5440" name="Plavecky klub Havirov">
          <ATHLETES>
            <ATHLETE firstname="Libor" lastname="Hracki" birthdate="1972-08-29" gender="M" nation="CZE" athleteid="5441">
              <RESULTS>
                <RESULT eventid="1212" points="341" reactiontime="+66" swimtime="00:02:22.15" resultid="5442" heatid="5832" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="150" swimtime="00:01:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="332" reactiontime="+66" swimtime="00:01:04.85" resultid="5443" heatid="5852" lane="8" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="337" reactiontime="+66" swimtime="00:00:36.28" resultid="5444" heatid="5869" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1503" points="326" reactiontime="+67" swimtime="00:02:54.55" resultid="5445" heatid="5948" lane="2" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                    <SPLIT distance="150" swimtime="00:02:08.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="327" reactiontime="+60" swimtime="00:05:07.78" resultid="5446" heatid="5981" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                    <SPLIT distance="200" swimtime="00:02:29.02" />
                    <SPLIT distance="250" swimtime="00:03:08.76" />
                    <SPLIT distance="300" swimtime="00:03:48.53" />
                    <SPLIT distance="350" swimtime="00:04:28.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRLOD" nation="POL" clubid="3292" name="MKS Trójka Łódź">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Szwedzki" birthdate="2000-12-12" gender="M" nation="POL" license="100905700604" swrid="4001538" athleteid="3293">
              <RESULTS>
                <RESULT eventid="1178" points="503" reactiontime="+70" swimtime="00:02:17.78" resultid="3294" heatid="5820" lane="3" entrytime="00:02:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="571" reactiontime="+69" swimtime="00:01:59.76" resultid="3295" heatid="5835" lane="5" entrytime="00:01:59.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                    <SPLIT distance="100" swimtime="00:00:58.77" />
                    <SPLIT distance="150" swimtime="00:01:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="478" reactiontime="+67" swimtime="00:02:18.35" resultid="3296" heatid="5900" lane="2" entrytime="00:02:19.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="426" reactiontime="+74" swimtime="00:02:20.30" resultid="3297" heatid="5908" lane="7" entrytime="00:02:18.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                    <SPLIT distance="150" swimtime="00:01:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="486" reactiontime="+69" swimtime="00:02:32.80" resultid="3298" heatid="5950" lane="3" entrytime="00:02:28.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="614" reactiontime="+71" swimtime="00:04:09.69" resultid="3299" heatid="5984" lane="3" entrytime="00:04:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:32.13" />
                    <SPLIT distance="200" swimtime="00:02:04.40" />
                    <SPLIT distance="250" swimtime="00:02:35.97" />
                    <SPLIT distance="300" swimtime="00:03:08.20" />
                    <SPLIT distance="350" swimtime="00:03:39.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" clubid="5302" name="Uks Wodnik 29 Katowice">
          <ATHLETES>
            <ATHLETE firstname="Agata" lastname="Kowalczyk" birthdate="2001-03-27" gender="F" nation="POL" athleteid="5308">
              <RESULTS>
                <RESULT eventid="1093" points="462" reactiontime="+71" swimtime="00:01:20.64" resultid="5309" heatid="5788" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="414" reactiontime="+70" swimtime="00:02:43.45" resultid="5310" heatid="5814" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:02:03.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="525" reactiontime="+68" swimtime="00:00:35.39" resultid="5311" heatid="5864" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1486" points="458" reactiontime="+75" swimtime="00:02:54.54" resultid="5312" heatid="5944" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:10.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Mróz" birthdate="1979-06-09" gender="F" nation="POL" athleteid="5317">
              <RESULTS>
                <RESULT eventid="1127" points="278" reactiontime="+90" swimtime="00:00:39.20" resultid="5318" heatid="5800" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1195" points="327" reactiontime="+81" swimtime="00:02:40.27" resultid="5319" heatid="5823" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:01:59.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="285" reactiontime="+93" swimtime="00:01:16.33" resultid="5320" heatid="5842" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="276" reactiontime="+96" swimtime="00:03:02.64" resultid="5321" heatid="5903" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:16.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="266" reactiontime="+96" swimtime="00:01:25.34" resultid="5322" heatid="5953" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="338" reactiontime="+99" swimtime="00:05:35.70" resultid="5323" heatid="5974" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:03.46" />
                    <SPLIT distance="200" swimtime="00:02:46.67" />
                    <SPLIT distance="250" swimtime="00:03:29.66" />
                    <SPLIT distance="300" swimtime="00:04:12.22" />
                    <SPLIT distance="350" swimtime="00:04:54.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Mrożiński" birthdate="1959-12-28" gender="M" nation="POL" athleteid="5313">
              <RESULTS>
                <RESULT eventid="1110" points="314" reactiontime="+81" swimtime="00:01:21.37" resultid="5314" heatid="5794" lane="3" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="345" reactiontime="+75" swimtime="00:00:35.97" resultid="5315" heatid="5872" lane="0" entrytime="00:00:35.70" />
                <RESULT eventid="1503" points="282" reactiontime="+82" swimtime="00:03:03.21" resultid="5316" heatid="5948" lane="6" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Koenig" birthdate="1987-04-21" gender="F" nation="POL" athleteid="5324">
              <RESULTS>
                <RESULT eventid="1093" points="104" swimtime="00:02:12.54" resultid="5325" heatid="5786" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="100" reactiontime="+71" swimtime="00:01:01.34" resultid="5326" heatid="5861" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1316" points="64" swimtime="00:02:20.69" resultid="5327" heatid="5877" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="102" swimtime="00:04:47.36" resultid="5328" heatid="5942" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.96" />
                    <SPLIT distance="100" swimtime="00:02:18.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Ogorzałek" birthdate="1999-08-22" gender="M" nation="POL" athleteid="5303">
              <RESULTS>
                <RESULT eventid="1299" points="560" reactiontime="+70" swimtime="00:00:30.63" resultid="5304" heatid="5873" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1333" points="534" reactiontime="+70" swimtime="00:01:00.73" resultid="5305" heatid="5892" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="632" swimtime="00:00:23.48" resultid="5306" heatid="5940" lane="7" entrytime="00:00:23.60" />
                <RESULT eventid="1605" points="614" reactiontime="+73" swimtime="00:04:09.61" resultid="5307" heatid="5984" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="150" swimtime="00:01:32.49" />
                    <SPLIT distance="200" swimtime="00:02:05.02" />
                    <SPLIT distance="250" swimtime="00:02:37.17" />
                    <SPLIT distance="300" swimtime="00:03:09.26" />
                    <SPLIT distance="350" swimtime="00:03:40.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="4282" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Pietrzak" birthdate="1996-01-01" gender="M" nation="POL" athleteid="5336">
              <RESULTS>
                <RESULT eventid="1110" points="380" reactiontime="+87" swimtime="00:01:16.40" resultid="5346" heatid="5793" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="404" swimtime="00:01:00.75" resultid="5347" heatid="5853" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="397" reactiontime="+79" swimtime="00:00:34.34" resultid="5348" heatid="5871" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1469" points="383" reactiontime="+81" swimtime="00:00:27.75" resultid="5349" heatid="5934" lane="6" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Pieślak" birthdate="1979-02-28" gender="M" nation="POL" license="102016700010" athleteid="4307">
              <RESULTS>
                <RESULT eventid="1110" points="338" reactiontime="+71" swimtime="00:01:19.43" resultid="4308" heatid="5794" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="4309" heatid="5833" lane="8" entrytime="00:02:28.00" />
                <RESULT eventid="1299" points="345" reactiontime="+70" swimtime="00:00:35.97" resultid="4310" heatid="5871" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1503" points="305" reactiontime="+76" swimtime="00:02:58.44" resultid="4311" heatid="5948" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                    <SPLIT distance="150" swimtime="00:02:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4312" heatid="5981" lane="9" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Mamrot" birthdate="1972-12-10" gender="M" nation="POL" license="102016700007" swrid="5471728" athleteid="4313">
              <RESULTS>
                <RESULT eventid="1110" points="224" reactiontime="+72" swimtime="00:01:31.10" resultid="4314" heatid="5791" lane="9" entrytime="00:01:41.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="239" reactiontime="+72" swimtime="00:00:40.67" resultid="4315" heatid="5868" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1333" points="204" reactiontime="+76" swimtime="00:01:23.64" resultid="4316" heatid="5885" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="211" reactiontime="+71" swimtime="00:03:21.68" resultid="4317" heatid="5947" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:32.80" />
                    <SPLIT distance="150" swimtime="00:02:26.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Gudaniec" birthdate="1960-08-26" gender="F" nation="POL" license="102016600015" swrid="4992893" athleteid="4318">
              <RESULTS>
                <RESULT eventid="1127" points="151" reactiontime="+65" swimtime="00:00:48.00" resultid="4319" heatid="5799" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1161" points="185" reactiontime="+85" swimtime="00:03:33.55" resultid="4320" heatid="5813" lane="1" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:42.75" />
                    <SPLIT distance="150" swimtime="00:02:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="179" reactiontime="+72" swimtime="00:01:40.19" resultid="4321" heatid="5878" lane="0" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="161" reactiontime="+69" swimtime="00:03:38.28" resultid="4322" heatid="5902" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.42" />
                    <SPLIT distance="100" swimtime="00:01:46.57" />
                    <SPLIT distance="150" swimtime="00:02:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="152" reactiontime="+72" swimtime="00:01:42.71" resultid="4323" heatid="5953" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="204" swimtime="00:06:37.05" resultid="4324" heatid="5974" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:31.23" />
                    <SPLIT distance="150" swimtime="00:02:21.93" />
                    <SPLIT distance="200" swimtime="00:03:13.25" />
                    <SPLIT distance="250" swimtime="00:04:04.60" />
                    <SPLIT distance="300" swimtime="00:04:56.22" />
                    <SPLIT distance="350" swimtime="00:05:47.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Winiarczyk" birthdate="1972-01-23" gender="M" nation="POL" license="102016700008" athleteid="4329">
              <RESULTS>
                <RESULT eventid="1144" points="249" reactiontime="+84" swimtime="00:00:35.31" resultid="4330" heatid="5807" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="4331" heatid="5833" lane="1" entrytime="00:02:25.00" />
                <RESULT eventid="1265" points="363" reactiontime="+75" swimtime="00:01:02.98" resultid="4332" heatid="5854" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="359" swimtime="00:00:28.35" resultid="4333" heatid="5934" lane="7" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Paziewska" birthdate="1974-09-05" gender="F" nation="POL" license="102016600012" swrid="5471732" athleteid="4300">
              <RESULTS>
                <RESULT eventid="1093" status="DNS" swimtime="00:00:00.00" resultid="4301" heatid="5787" lane="9" entrytime="00:01:44.00" />
                <RESULT eventid="1195" points="283" reactiontime="+87" swimtime="00:02:48.01" resultid="4302" heatid="5824" lane="9" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="323" reactiontime="+82" swimtime="00:01:13.19" resultid="4303" heatid="5842" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="248" reactiontime="+89" swimtime="00:00:45.41" resultid="4304" heatid="5862" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1451" points="332" swimtime="00:00:33.09" resultid="4305" heatid="5920" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1588" points="273" reactiontime="+95" swimtime="00:06:00.40" resultid="4306" heatid="5974" lane="3" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                    <SPLIT distance="200" swimtime="00:02:54.10" />
                    <SPLIT distance="250" swimtime="00:03:40.44" />
                    <SPLIT distance="300" swimtime="00:04:27.46" />
                    <SPLIT distance="350" swimtime="00:05:14.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Gudaniec" birthdate="1988-01-01" gender="F" nation="POL" athleteid="5333">
              <RESULTS>
                <RESULT eventid="1161" points="312" swimtime="00:02:59.55" resultid="5341" heatid="5814" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:16.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="345" reactiontime="+79" swimtime="00:02:37.36" resultid="5342" heatid="5824" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:55.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="352" reactiontime="+72" swimtime="00:01:11.14" resultid="5343" heatid="5843" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="322" reactiontime="+70" swimtime="00:01:22.41" resultid="5344" heatid="5879" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="359" reactiontime="+80" swimtime="00:05:28.91" resultid="5345" heatid="5975" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                    <SPLIT distance="200" swimtime="00:02:39.18" />
                    <SPLIT distance="250" swimtime="00:03:21.47" />
                    <SPLIT distance="300" swimtime="00:04:03.84" />
                    <SPLIT distance="350" swimtime="00:04:46.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Wróblewski" birthdate="1990-01-01" gender="M" nation="POL" athleteid="5331">
              <RESULTS>
                <RESULT eventid="1076" points="594" reactiontime="+70" swimtime="00:00:25.87" resultid="5352" heatid="5782" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1178" points="526" reactiontime="+75" swimtime="00:02:15.81" resultid="5353" heatid="5819" lane="4" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="100" swimtime="00:01:03.55" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="484" reactiontime="+75" swimtime="00:02:17.82" resultid="5354" heatid="5900" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="150" swimtime="00:01:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="584" reactiontime="+70" swimtime="00:00:57.15" resultid="5355" heatid="5970" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="517" reactiontime="+72" swimtime="00:04:24.35" resultid="5356" heatid="5983" lane="2" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:39.60" />
                    <SPLIT distance="200" swimtime="00:02:13.82" />
                    <SPLIT distance="250" swimtime="00:02:47.98" />
                    <SPLIT distance="300" swimtime="00:03:21.49" />
                    <SPLIT distance="350" swimtime="00:03:53.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Stankiewicz-Majkowska" birthdate="1972-12-06" gender="F" nation="POL" license="102016600011" swrid="4992894" athleteid="4283">
              <RESULTS>
                <RESULT eventid="1059" points="150" swimtime="00:00:45.80" resultid="4284" heatid="5768" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1161" points="188" swimtime="00:03:32.47" resultid="4285" heatid="5813" lane="7" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:41.37" />
                    <SPLIT distance="150" swimtime="00:02:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="177" swimtime="00:01:40.48" resultid="4286" heatid="5878" lane="9" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="152" reactiontime="+102" swimtime="00:03:42.63" resultid="4287" heatid="5902" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.77" />
                    <SPLIT distance="100" swimtime="00:01:51.20" />
                    <SPLIT distance="150" swimtime="00:02:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="213" reactiontime="+95" swimtime="00:03:45.26" resultid="4288" heatid="5943" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                    <SPLIT distance="100" swimtime="00:01:48.54" />
                    <SPLIT distance="150" swimtime="00:02:47.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Rutkowski" birthdate="1974-02-20" gender="M" nation="POL" license="102016700018" swrid="4992794" athleteid="4289">
              <RESULTS>
                <RESULT eventid="1076" points="327" reactiontime="+88" swimtime="00:00:31.57" resultid="4290" heatid="5777" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1178" points="264" reactiontime="+87" swimtime="00:02:50.73" resultid="4291" heatid="5818" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:02:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="223" reactiontime="+88" swimtime="00:02:58.33" resultid="4292" heatid="5899" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:11.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="255" swimtime="00:01:15.30" resultid="4293" heatid="5967" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kruk" birthdate="1982-01-01" gender="M" nation="POL" athleteid="5337">
              <RESULTS>
                <RESULT eventid="1469" points="297" reactiontime="+75" swimtime="00:00:30.19" resultid="5350" heatid="5932" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1605" points="242" reactiontime="+75" swimtime="00:05:40.14" resultid="5351" heatid="5980" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:56.41" />
                    <SPLIT distance="200" swimtime="00:02:39.52" />
                    <SPLIT distance="250" swimtime="00:03:23.82" />
                    <SPLIT distance="300" swimtime="00:04:08.84" />
                    <SPLIT distance="350" swimtime="00:04:55.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lidia" lastname="Mikołajczyk" birthdate="1987-04-29" gender="F" nation="POL" license="102016600013" swrid="5471730" athleteid="4334">
              <RESULTS>
                <RESULT eventid="1195" points="367" swimtime="00:02:34.23" resultid="4335" heatid="5824" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="391" reactiontime="+102" swimtime="00:01:08.69" resultid="4336" heatid="5843" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="385" reactiontime="+97" swimtime="00:01:17.66" resultid="4337" heatid="5878" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="401" reactiontime="+85" swimtime="00:00:31.09" resultid="4338" heatid="5920" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1588" points="355" reactiontime="+95" swimtime="00:05:30.07" resultid="4339" heatid="5975" lane="0" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:57.97" />
                    <SPLIT distance="200" swimtime="00:02:40.41" />
                    <SPLIT distance="250" swimtime="00:03:23.26" />
                    <SPLIT distance="300" swimtime="00:04:06.57" />
                    <SPLIT distance="350" swimtime="00:04:49.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Ćwikła" birthdate="1974-08-22" gender="M" nation="POL" license="102016700002" athleteid="4325">
              <RESULTS>
                <RESULT eventid="1144" points="295" reactiontime="+65" swimtime="00:00:33.36" resultid="4326" heatid="5808" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1401" points="273" reactiontime="+68" swimtime="00:02:42.64" resultid="4327" heatid="5906" lane="3" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:00.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="265" reactiontime="+63" swimtime="00:01:15.18" resultid="4328" heatid="5960" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="398" reactiontime="+75" swimtime="00:01:51.15" resultid="5334" heatid="5913" lane="4" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.79" />
                    <SPLIT distance="100" swimtime="00:00:53.48" />
                    <SPLIT distance="150" swimtime="00:01:23.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5331" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4307" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4325" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4329" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="369" reactiontime="+62" swimtime="00:02:06.06" resultid="5339" heatid="5988" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4325" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="4307" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4289" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="5331" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="325" reactiontime="+80" swimtime="00:01:58.92" resultid="5335" heatid="5913" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="100" swimtime="00:00:59.08" />
                    <SPLIT distance="150" swimtime="00:01:28.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5336" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4313" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4289" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5337" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="296" reactiontime="+80" swimtime="00:02:15.62" resultid="5340" heatid="5988" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:01:45.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5336" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="4313" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4329" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="5337" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="294" swimtime="00:02:19.03" resultid="5332" heatid="5910" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:15.26" />
                    <SPLIT distance="150" swimtime="00:01:46.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4318" number="1" />
                    <RELAYPOSITION athleteid="5333" number="2" />
                    <RELAYPOSITION athleteid="4334" number="3" />
                    <RELAYPOSITION athleteid="4300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="269" reactiontime="+89" swimtime="00:02:38.51" resultid="5338" heatid="5986" lane="7" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                    <SPLIT distance="150" swimtime="00:02:05.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4283" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="4334" number="2" />
                    <RELAYPOSITION athleteid="5333" number="3" />
                    <RELAYPOSITION athleteid="4300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="274" reactiontime="+72" swimtime="00:02:27.98" resultid="5329" heatid="5838" lane="8" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                    <SPLIT distance="150" swimtime="00:01:55.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4325" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4318" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4289" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4300" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="287" reactiontime="+75" swimtime="00:02:25.77" resultid="5330" heatid="5838" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:00.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4329" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4283" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4334" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="5331" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="2873" name="SPK Kupele Piestany">
          <ATHLETES>
            <ATHLETE firstname="Miroslava" lastname="Samuhelova" birthdate="1975-01-01" gender="F" nation="SVK" swrid="5448431" athleteid="2872">
              <RESULTS>
                <RESULT eventid="1093" points="296" reactiontime="+83" swimtime="00:01:33.57" resultid="2874" heatid="5787" lane="2" entrytime="00:01:35.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="242" reactiontime="+82" swimtime="00:01:30.67" resultid="2875" heatid="5878" lane="2" entrytime="00:01:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="266" swimtime="00:03:29.17" resultid="2876" heatid="5944" lane="7" entrytime="00:03:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:37.45" />
                    <SPLIT distance="150" swimtime="00:02:33.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martin" lastname="Babsky" birthdate="1972-01-01" gender="M" nation="SVK" swrid="5439025" athleteid="2877">
              <RESULTS>
                <RESULT eventid="1076" points="359" reactiontime="+83" swimtime="00:00:30.60" resultid="2878" heatid="5780" lane="8" entrytime="00:00:29.90" />
                <RESULT eventid="1265" points="423" reactiontime="+79" swimtime="00:00:59.84" resultid="2879" heatid="5855" lane="1" entrytime="00:01:00.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="440" reactiontime="+75" swimtime="00:00:26.50" resultid="2880" heatid="5936" lane="4" entrytime="00:00:26.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pavel" lastname="Škodný" birthdate="1969-01-01" gender="M" nation="SVK" swrid="4688816" athleteid="2881">
              <RESULTS>
                <RESULT eventid="1178" points="329" swimtime="00:02:38.71" resultid="2882" heatid="5819" lane="9" entrytime="00:02:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:02:02.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="281" reactiontime="+81" swimtime="00:02:41.13" resultid="2883" heatid="5907" lane="8" entrytime="00:02:39.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:02:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="270" reactiontime="+82" swimtime="00:01:14.69" resultid="2884" heatid="5960" lane="6" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5224" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Rólczyński" birthdate="1977-01-01" gender="M" nation="POL" athleteid="5223">
              <RESULTS>
                <RESULT eventid="1144" points="247" reactiontime="+71" swimtime="00:00:35.40" resultid="5225" heatid="5808" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1333" points="277" reactiontime="+68" swimtime="00:01:15.56" resultid="5226" heatid="5890" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="14" clubid="4505" name="Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Wilczęga" birthdate="1981-10-24" gender="M" nation="POL" license="106614700042" swrid="4992879" athleteid="4506">
              <RESULTS>
                <RESULT eventid="1076" points="367" reactiontime="+71" swimtime="00:00:30.37" resultid="4507" heatid="5780" lane="0" entrytime="00:00:29.95" />
                <RESULT eventid="1265" points="441" reactiontime="+69" swimtime="00:00:59.02" resultid="4508" heatid="5856" lane="6" entrytime="00:00:58.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="445" swimtime="00:00:26.39" resultid="4509" heatid="5937" lane="7" entrytime="00:00:26.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" license="506614700212" swrid="4992696" athleteid="4510">
              <RESULTS>
                <RESULT eventid="1144" points="123" reactiontime="+83" swimtime="00:00:44.64" resultid="4511" heatid="5803" lane="2" />
                <RESULT eventid="1212" points="139" reactiontime="+94" swimtime="00:03:11.49" resultid="4512" heatid="5827" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                    <SPLIT distance="150" swimtime="00:02:19.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="160" reactiontime="+62" swimtime="00:01:22.70" resultid="4513" heatid="5846" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="133" reactiontime="+76" swimtime="00:01:36.49" resultid="4514" heatid="5882" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="189" reactiontime="+79" swimtime="00:00:35.10" resultid="4515" heatid="5923" lane="5" />
                <RESULT eventid="1605" points="125" reactiontime="+88" swimtime="00:07:03.87" resultid="4516" heatid="5976" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:33.34" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                    <SPLIT distance="200" swimtime="00:03:18.48" />
                    <SPLIT distance="250" swimtime="00:04:14.67" />
                    <SPLIT distance="300" swimtime="00:05:13.13" />
                    <SPLIT distance="350" swimtime="00:06:10.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="4416" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" swrid="4595659" athleteid="4485">
              <RESULTS>
                <RESULT eventid="1212" points="391" reactiontime="+87" swimtime="00:02:15.81" resultid="4486" heatid="5833" lane="4" entrytime="00:02:16.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="150" swimtime="00:01:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="311" reactiontime="+81" swimtime="00:02:39.66" resultid="4487" heatid="5899" lane="6" entrytime="00:02:41.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="367" reactiontime="+90" swimtime="00:04:56.36" resultid="4488" heatid="5982" lane="6" entrytime="00:04:58.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                    <SPLIT distance="200" swimtime="00:02:24.07" />
                    <SPLIT distance="250" swimtime="00:03:01.49" />
                    <SPLIT distance="300" swimtime="00:03:39.28" />
                    <SPLIT distance="350" swimtime="00:04:16.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Osik" birthdate="1976-01-02" gender="M" nation="POL" license="500115700521" athleteid="4449">
              <RESULTS>
                <RESULT eventid="1144" points="318" reactiontime="+67" swimtime="00:00:32.54" resultid="4450" heatid="5808" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1212" points="410" reactiontime="+93" swimtime="00:02:13.74" resultid="4451" heatid="5834" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.81" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="414" swimtime="00:01:00.28" resultid="4452" heatid="5855" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="328" reactiontime="+81" swimtime="00:02:33.06" resultid="4453" heatid="5907" lane="7" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:01:54.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="344" reactiontime="+78" swimtime="00:01:08.93" resultid="4454" heatid="5961" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="402" reactiontime="+93" swimtime="00:04:47.41" resultid="4455" heatid="5982" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:45.73" />
                    <SPLIT distance="200" swimtime="00:02:22.88" />
                    <SPLIT distance="250" swimtime="00:02:59.90" />
                    <SPLIT distance="300" swimtime="00:03:36.70" />
                    <SPLIT distance="350" swimtime="00:04:12.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuca" birthdate="1994-07-23" gender="M" nation="POL" license="100115700396" swrid="4213120" athleteid="4473">
              <RESULTS>
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="4474" heatid="5820" lane="5" entrytime="00:02:10.50" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="4475" heatid="5858" lane="3" entrytime="00:00:52.32" entrycourse="SCM" />
                <RESULT eventid="1333" points="564" reactiontime="+63" swimtime="00:00:59.64" resultid="4476" heatid="5893" lane="2" entrytime="00:00:59.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="617" reactiontime="+62" swimtime="00:00:23.68" resultid="4477" heatid="5940" lane="3" entrytime="00:00:23.30" />
                <RESULT eventid="1571" points="583" reactiontime="+64" swimtime="00:00:57.19" resultid="4478" heatid="5971" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" swrid="4754727" athleteid="4479">
              <RESULTS>
                <RESULT eventid="1195" points="228" reactiontime="+100" swimtime="00:03:00.72" resultid="4480" heatid="5821" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:27.30" />
                    <SPLIT distance="150" swimtime="00:02:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="219" reactiontime="+107" swimtime="00:01:23.24" resultid="4481" heatid="5840" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="199" reactiontime="+127" swimtime="00:03:23.60" resultid="4482" heatid="5901" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                    <SPLIT distance="100" swimtime="00:01:40.87" />
                    <SPLIT distance="150" swimtime="00:02:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="178" reactiontime="+134" swimtime="00:01:37.49" resultid="4483" heatid="5951" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="245" reactiontime="+97" swimtime="00:06:13.60" resultid="4484" heatid="5974" lane="8" entrytime="00:06:15.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:28.88" />
                    <SPLIT distance="150" swimtime="00:02:16.50" />
                    <SPLIT distance="200" swimtime="00:03:04.17" />
                    <SPLIT distance="250" swimtime="00:03:52.25" />
                    <SPLIT distance="300" swimtime="00:04:39.65" />
                    <SPLIT distance="350" swimtime="00:05:27.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dowgiert" birthdate="1990-01-01" gender="F" nation="POL" swrid="4071947" athleteid="5638">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1059" points="827" reactiontime="+62" status="EXH" swimtime="00:00:25.97" resultid="5639" heatid="5771" lane="4" entrytime="00:00:25.69" entrycourse="SCM" />
                <RESULT eventid="1247" reactiontime="+65" status="DNF" swimtime="00:00:00.00" resultid="5640" heatid="5844" lane="4" entrytime="00:00:54.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="5641" heatid="5922" lane="4" entrytime="00:00:24.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Lesiński" birthdate="1944-04-13" gender="M" nation="POL" license="500115700616" swrid="4188190" athleteid="4461">
              <RESULTS>
                <RESULT eventid="1144" points="103" reactiontime="+77" swimtime="00:00:47.29" resultid="4462" heatid="5804" lane="3" entrytime="00:00:51.06" entrycourse="SCM" />
                <RESULT eventid="1212" points="97" reactiontime="+115" swimtime="00:03:35.87" resultid="4463" heatid="5827" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                    <SPLIT distance="100" swimtime="00:01:41.25" />
                    <SPLIT distance="150" swimtime="00:02:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="107" reactiontime="+103" swimtime="00:00:53.16" resultid="4464" heatid="5867" lane="2" entrytime="00:00:54.00" />
                <RESULT eventid="1333" points="95" reactiontime="+112" swimtime="00:01:47.93" resultid="4465" heatid="5883" lane="4" entrytime="00:01:49.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="106" reactiontime="+112" swimtime="00:00:42.48" resultid="4466" heatid="5926" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1537" points="90" reactiontime="+81" swimtime="00:01:47.78" resultid="4467" heatid="5958" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" swrid="4992782" athleteid="4456">
              <RESULTS>
                <RESULT eventid="1144" points="325" reactiontime="+64" swimtime="00:00:32.29" resultid="4457" heatid="5809" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1212" points="369" reactiontime="+84" swimtime="00:02:18.49" resultid="4458" heatid="5833" lane="3" entrytime="00:02:18.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="296" reactiontime="+70" swimtime="00:02:38.37" resultid="4459" heatid="5907" lane="1" entrytime="00:02:36.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="319" reactiontime="+67" swimtime="00:01:10.72" resultid="4460" heatid="5961" lane="6" entrytime="00:01:09.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Smektała" birthdate="2004-01-01" gender="F" nation="POL" swrid="5114691" athleteid="5642">
              <RESULTS>
                <RESULT eventid="1059" points="574" reactiontime="+68" status="EXH" swimtime="00:00:29.32" resultid="5643" heatid="5771" lane="5" entrytime="00:00:28.64" entrycourse="SCM" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="5644" heatid="5921" lane="5" entrytime="00:00:28.14" entrycourse="SCM" />
                <RESULT eventid="1247" status="DNS" swimtime="00:00:00.00" resultid="5645" heatid="5844" lane="2" entrytime="00:01:00.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Wieja" birthdate="1978-09-08" gender="M" nation="POL" license="500115700467" swrid="5331775" athleteid="4468">
              <RESULTS>
                <RESULT eventid="1144" points="382" reactiontime="+59" swimtime="00:00:30.61" resultid="4469" heatid="5810" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1333" points="431" reactiontime="+67" swimtime="00:01:05.21" resultid="4470" heatid="5892" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="452" reactiontime="+66" swimtime="00:00:26.26" resultid="4471" heatid="5937" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1537" points="363" reactiontime="+62" swimtime="00:01:07.72" resultid="4472" heatid="5962" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Zajączek" birthdate="1976-07-17" gender="F" nation="POL" license="500115600524" swrid="5455051" athleteid="4417">
              <RESULTS>
                <RESULT eventid="1059" points="67" swimtime="00:00:59.80" resultid="4418" heatid="5767" lane="5" />
                <RESULT eventid="1093" points="130" swimtime="00:02:03.05" resultid="4419" heatid="5784" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="76" swimtime="00:01:58.17" resultid="4420" heatid="5839" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="129" swimtime="00:00:56.48" resultid="4421" heatid="5861" lane="3" entrytime="00:00:58.27" entrycourse="SCM" />
                <RESULT eventid="1451" points="86" swimtime="00:00:51.83" resultid="4422" heatid="5916" lane="2" />
                <RESULT eventid="1486" points="147" swimtime="00:04:14.49" resultid="4423" heatid="5943" lane="0" entrytime="00:04:25.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.65" />
                    <SPLIT distance="100" swimtime="00:02:04.17" />
                    <SPLIT distance="150" swimtime="00:03:11.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="4440">
              <RESULTS>
                <RESULT eventid="1093" points="110" reactiontime="+99" swimtime="00:02:10.05" resultid="4441" heatid="5786" lane="7" entrytime="00:02:08.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="112" swimtime="00:04:38.86" resultid="4443" heatid="5943" lane="9" entrytime="00:04:30.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.19" />
                    <SPLIT distance="100" swimtime="00:02:14.46" />
                    <SPLIT distance="150" swimtime="00:03:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="109" reactiontime="+103" swimtime="00:00:59.67" resultid="5377" heatid="5861" lane="5" entrytime="00:00:57.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="4444">
              <RESULTS>
                <RESULT eventid="1110" points="256" reactiontime="+88" swimtime="00:01:27.10" resultid="4445" heatid="5792" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="272" reactiontime="+84" swimtime="00:00:38.95" resultid="4446" heatid="5870" lane="1" entrytime="00:00:38.79" entrycourse="SCM" />
                <RESULT eventid="1333" points="199" swimtime="00:01:24.38" resultid="4447" heatid="5887" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="234" reactiontime="+85" swimtime="00:03:14.97" resultid="4448" heatid="5948" lane="0" entrytime="00:03:08.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:31.87" />
                    <SPLIT distance="150" swimtime="00:02:22.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Chudy" birthdate="1997-01-01" gender="M" nation="POL" swrid="4286914" athleteid="5646">
              <RESULTS>
                <RESULT eventid="1076" points="723" reactiontime="+65" status="EXH" swimtime="00:00:24.23" resultid="5647" heatid="5783" lane="4" entrytime="00:00:23.55" entrycourse="SCM" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5648" heatid="5893" lane="4" entrytime="00:00:53.61" entrycourse="SCM" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5649" heatid="5971" lane="4" entrytime="00:00:52.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" swrid="5312534" athleteid="4424">
              <RESULTS>
                <RESULT eventid="1076" points="476" reactiontime="+69" swimtime="00:00:27.84" resultid="4425" heatid="5782" lane="4" entrytime="00:00:26.90" entrycourse="SCM" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1110" points="561" reactiontime="+71" swimtime="00:01:07.06" resultid="4426" heatid="5796" lane="1" entrytime="00:01:06.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1299" points="623" reactiontime="+65" swimtime="00:00:29.55" resultid="4427" heatid="5874" lane="3" entrytime="00:00:29.20" entrycourse="SCM" />
                <RESULT eventid="1469" points="486" reactiontime="+68" swimtime="00:00:25.63" resultid="4428" heatid="5939" lane="6" entrytime="00:00:24.90" entrycourse="SCM" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4429" heatid="5970" lane="1" entrytime="00:01:03.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Thiem" birthdate="1963-02-17" gender="M" nation="POL" license="100115700345" swrid="4754725" athleteid="4430">
              <RESULTS>
                <RESULT eventid="1076" points="162" reactiontime="+98" swimtime="00:00:39.84" resultid="4431" heatid="5774" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1212" points="150" swimtime="00:03:06.81" resultid="4432" heatid="5830" lane="9" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:29.40" />
                    <SPLIT distance="150" swimtime="00:02:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="139" reactiontime="+106" swimtime="00:03:28.73" resultid="4433" heatid="5898" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:44.39" />
                    <SPLIT distance="150" swimtime="00:02:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="145" reactiontime="+102" swimtime="00:01:30.74" resultid="4434" heatid="5967" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" swrid="5062813" athleteid="4435">
              <RESULTS>
                <RESULT eventid="1076" points="517" reactiontime="+70" swimtime="00:00:27.09" resultid="4436" heatid="5783" lane="9" entrytime="00:00:26.81" entrycourse="SCM" />
                <RESULT eventid="1265" points="584" swimtime="00:00:53.76" resultid="4437" heatid="5858" lane="7" entrytime="00:00:53.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="606" reactiontime="+72" swimtime="00:00:23.82" resultid="4438" heatid="5940" lane="9" entrytime="00:00:24.45" entrycourse="SCM" />
                <RESULT eventid="1571" points="505" swimtime="00:00:59.98" resultid="4439" heatid="5970" lane="7" entrytime="00:01:03.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1442" points="529" reactiontime="+68" swimtime="00:01:41.14" resultid="4490" heatid="5914" lane="3" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.65" />
                    <SPLIT distance="100" swimtime="00:00:50.65" />
                    <SPLIT distance="150" swimtime="00:01:18.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4468" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4424" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4456" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4473" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="524" reactiontime="+59" swimtime="00:01:52.12" resultid="4492" heatid="5989" lane="5" entrytime="00:01:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                    <SPLIT distance="150" swimtime="00:01:24.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4468" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="4424" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="4473" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="4456" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="281" reactiontime="+82" swimtime="00:02:04.87" resultid="4491" heatid="5913" lane="0" entrytime="00:02:01.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:28.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4449" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="4485" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="4444" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4430" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="223" reactiontime="+77" swimtime="00:02:29.04" resultid="4493" heatid="5988" lane="0" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:47.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4435" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4444" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4430" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4461" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="172" reactiontime="+61" swimtime="00:02:52.90" resultid="4489" heatid="5836" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                    <SPLIT distance="150" swimtime="00:02:28.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4435" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4417" number="2" />
                    <RELAYPOSITION athleteid="4440" number="3" />
                    <RELAYPOSITION athleteid="4468" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3140" name="Masters Łódź">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Olejarczyk" birthdate="1979-06-12" gender="M" nation="POL" license="503605700007" swrid="4992959" athleteid="3166">
              <RESULTS>
                <RESULT eventid="1076" points="366" swimtime="00:00:30.40" resultid="3167" heatid="5780" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1265" points="391" swimtime="00:01:01.43" resultid="3168" heatid="5856" lane="7" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" status="DNS" swimtime="00:00:00.00" resultid="3169" heatid="5899" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="1469" points="384" swimtime="00:00:27.72" resultid="3170" heatid="5937" lane="9" entrytime="00:00:26.50" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="3171" heatid="5970" lane="0" entrytime="00:01:06.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kurstak-Jagiełło" birthdate="1981-06-30" gender="F" nation="POL" license="503605600022" athleteid="3141">
              <RESULTS>
                <RESULT eventid="1195" points="411" reactiontime="+89" swimtime="00:02:28.44" resultid="3142" heatid="5821" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="447" reactiontime="+87" swimtime="00:01:05.69" resultid="3143" heatid="5840" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="445" reactiontime="+84" swimtime="00:00:30.03" resultid="3144" heatid="5920" lane="3" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Karczmarczyk" birthdate="1980-04-16" gender="M" nation="POL" license="103605700004" swrid="4992955" athleteid="3184">
              <RESULTS>
                <RESULT eventid="1110" points="271" reactiontime="+90" swimtime="00:01:25.51" resultid="3185" heatid="5791" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="204" reactiontime="+97" swimtime="00:03:06.12" resultid="3186" heatid="5817" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="296" reactiontime="+91" swimtime="00:00:37.86" resultid="3187" heatid="5869" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1333" points="222" reactiontime="+91" swimtime="00:01:21.38" resultid="3188" heatid="5885" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="302" reactiontime="+90" swimtime="00:00:30.02" resultid="3189" heatid="5928" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1503" points="223" reactiontime="+91" swimtime="00:03:17.97" resultid="3190" heatid="5947" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                    <SPLIT distance="100" swimtime="00:01:33.45" />
                    <SPLIT distance="150" swimtime="00:02:29.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Woźniak" birthdate="1981-08-25" gender="M" nation="POL" license="503605700034" swrid="5484423" athleteid="3154">
              <RESULTS>
                <RESULT eventid="1076" points="448" reactiontime="+76" swimtime="00:00:28.41" resultid="3155" heatid="5782" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1144" points="409" reactiontime="+60" swimtime="00:00:29.91" resultid="3156" heatid="5811" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="1401" points="395" reactiontime="+59" swimtime="00:02:23.91" resultid="3157" heatid="5908" lane="0" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.48" />
                    <SPLIT distance="150" swimtime="00:01:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="430" reactiontime="+64" swimtime="00:01:04.01" resultid="3158" heatid="5962" lane="0" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="503605600029" swrid="5464091" athleteid="3159">
              <RESULTS>
                <RESULT eventid="1161" points="170" reactiontime="+102" swimtime="00:03:39.61" resultid="3160" heatid="5812" lane="4" entrytime="00:03:48.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                    <SPLIT distance="100" swimtime="00:01:51.85" />
                    <SPLIT distance="150" swimtime="00:02:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="186" swimtime="00:03:13.13" resultid="3161" heatid="5823" lane="9" entrytime="00:03:23.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                    <SPLIT distance="150" swimtime="00:02:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="146" reactiontime="+102" swimtime="00:03:46.96" resultid="3162" heatid="5895" lane="8" entrytime="00:04:02.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:46.36" />
                    <SPLIT distance="150" swimtime="00:02:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="110" reactiontime="+94" swimtime="00:04:08.23" resultid="3163" heatid="5901" lane="4" entrytime="00:04:27.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                    <SPLIT distance="100" swimtime="00:02:03.33" />
                    <SPLIT distance="150" swimtime="00:03:06.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="205" reactiontime="+103" swimtime="00:03:47.87" resultid="3164" heatid="5943" lane="1" entrytime="00:03:55.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.51" />
                    <SPLIT distance="100" swimtime="00:01:53.03" />
                    <SPLIT distance="150" swimtime="00:02:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="172" reactiontime="+110" swimtime="00:07:00.47" resultid="3165" heatid="5973" lane="2" entrytime="00:07:07.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:37.74" />
                    <SPLIT distance="150" swimtime="00:02:30.28" />
                    <SPLIT distance="200" swimtime="00:03:25.05" />
                    <SPLIT distance="250" swimtime="00:04:19.76" />
                    <SPLIT distance="300" swimtime="00:05:13.66" />
                    <SPLIT distance="350" swimtime="00:06:08.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Lipka" birthdate="1980-12-18" gender="M" nation="POL" license="503605700025" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1076" points="165" reactiontime="+95" swimtime="00:00:39.64" resultid="3180" heatid="5775" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1178" points="170" reactiontime="+98" swimtime="00:03:17.78" resultid="3181" heatid="5816" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                    <SPLIT distance="150" swimtime="00:02:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="166" reactiontime="+98" swimtime="00:01:29.55" resultid="3182" heatid="5885" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="106" reactiontime="+106" swimtime="00:01:40.78" resultid="3183" heatid="5966" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Wilińska-Nowak" birthdate="1980-04-16" gender="F" nation="POL" license="103605600002" athleteid="3150">
              <RESULTS>
                <RESULT eventid="1059" points="460" reactiontime="+96" swimtime="00:00:31.57" resultid="3151" heatid="5767" lane="7" />
                <RESULT eventid="1350" points="388" reactiontime="+94" swimtime="00:02:43.96" resultid="3152" heatid="5894" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:01:59.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="465" swimtime="00:01:10.46" resultid="3153" heatid="5963" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Kruszyna-Kotulski" birthdate="1979-05-25" gender="M" nation="POL" license="503605700044" athleteid="3145">
              <RESULTS>
                <RESULT eventid="1076" points="334" reactiontime="+73" swimtime="00:00:31.32" resultid="3146" heatid="5773" lane="0" />
                <RESULT eventid="1144" points="202" reactiontime="+74" swimtime="00:00:37.85" resultid="3147" heatid="5804" lane="0" />
                <RESULT eventid="1333" points="276" reactiontime="+75" swimtime="00:01:15.68" resultid="3148" heatid="5882" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="289" reactiontime="+76" swimtime="00:00:30.49" resultid="3149" heatid="5924" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Adamska" birthdate="1984-09-25" gender="F" nation="POL" license="503605600036" swrid="5464086" athleteid="3172">
              <RESULTS>
                <RESULT eventid="1059" points="302" swimtime="00:00:36.31" resultid="3173" heatid="5769" lane="5" entrytime="00:00:37.07" entrycourse="SCM" />
                <RESULT eventid="1127" points="235" reactiontime="+72" swimtime="00:00:41.43" resultid="3174" heatid="5800" lane="0" entrytime="00:00:40.12" entrycourse="SCM" />
                <RESULT eventid="1247" points="285" reactiontime="+65" swimtime="00:01:16.33" resultid="3175" heatid="5841" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="162" reactiontime="+74" swimtime="00:03:39.09" resultid="3176" heatid="5894" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:34.86" />
                    <SPLIT distance="150" swimtime="00:02:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="232" reactiontime="+69" swimtime="00:01:29.26" resultid="3177" heatid="5953" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="231" reactiontime="+71" swimtime="00:01:28.97" resultid="3178" heatid="5963" lane="5" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="305" reactiontime="+71" swimtime="00:02:01.48" resultid="3192" heatid="5913" lane="6" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:01:02.70" />
                    <SPLIT distance="150" swimtime="00:01:32.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3166" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3179" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3184" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3145" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1646" points="326" reactiontime="+49" swimtime="00:02:11.29" resultid="3193" heatid="5989" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3154" number="1" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3184" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3166" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3179" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="342" reactiontime="+60" swimtime="00:02:17.46" resultid="3191" heatid="5838" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:48.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3154" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3159" number="2" />
                    <RELAYPOSITION athleteid="3166" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3141" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="3301" name="KPS Nereus Žilina">
          <ATHLETES>
            <ATHLETE firstname="Rastislav" lastname="Pavlik" birthdate="1960-01-01" gender="M" nation="SVK" swrid="4269975" athleteid="3300">
              <RESULTS>
                <RESULT eventid="1076" points="364" reactiontime="+78" swimtime="00:00:30.44" resultid="3302" heatid="5779" lane="7" entrytime="00:00:30.49" />
                <RESULT eventid="1144" points="337" reactiontime="+80" swimtime="00:00:31.91" resultid="3303" heatid="5810" lane="0" entrytime="00:00:31.49" />
                <RESULT eventid="1299" points="382" reactiontime="+79" swimtime="00:00:34.79" resultid="3304" heatid="5872" lane="5" entrytime="00:00:34.49" />
                <RESULT eventid="1333" points="307" swimtime="00:01:12.99" resultid="3305" heatid="5891" lane="7" entrytime="00:01:08.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="364" reactiontime="+74" swimtime="00:00:28.22" resultid="3306" heatid="5935" lane="0" entrytime="00:00:27.49" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="3307" heatid="5961" lane="3" entrytime="00:01:08.49" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2707" name="niezrzeszona" />
        <CLUB type="CLUB" nation="POL" clubid="1675" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Płonka" birthdate="1948-01-01" gender="M" nation="POL" swrid="4754750" athleteid="1674">
              <RESULTS>
                <RESULT eventid="1076" points="48" reactiontime="+103" swimtime="00:00:59.79" resultid="1676" heatid="5773" lane="7" entrytime="00:01:00.00" />
                <RESULT eventid="1212" points="39" reactiontime="+105" swimtime="00:04:51.85" resultid="1677" heatid="5828" lane="0" entrytime="00:04:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.32" />
                    <SPLIT distance="100" swimtime="00:02:21.31" />
                    <SPLIT distance="150" swimtime="00:03:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="40" reactiontime="+134" swimtime="00:02:10.79" resultid="1678" heatid="5847" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="25" reactiontime="+107" swimtime="00:06:09.83" resultid="1679" heatid="5896" lane="4" entrytime="00:05:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.32" />
                    <SPLIT distance="100" swimtime="00:02:57.25" />
                    <SPLIT distance="150" swimtime="00:04:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="66" reactiontime="+103" swimtime="00:00:49.64" resultid="1680" heatid="5925" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1571" points="24" reactiontime="+113" swimtime="00:02:45.59" resultid="1681" heatid="5965" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GER" clubid="2755" name="BerlinerTSC">
          <ATHLETES>
            <ATHLETE firstname="Martin" lastname="Klein" birthdate="1979-01-01" gender="M" nation="GER" swrid="4125319" athleteid="2754">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2756" heatid="5782" lane="8" entrytime="00:00:27.60" />
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="2757" heatid="5820" lane="2" entrytime="00:02:19.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="2758" heatid="5892" lane="3" entrytime="00:01:03.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="2759" heatid="5908" lane="6" entrytime="00:02:16.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="2760" heatid="5962" lane="7" entrytime="00:01:02.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="2761" heatid="5983" lane="0" entrytime="00:04:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="2784" name="Dzukijos vandenis">
          <ATHLETES>
            <ATHLETE firstname="Sigitas" lastname="Katkevicius" birthdate="1957-01-01" gender="M" nation="LTU" swrid="4418116" athleteid="2783">
              <RESULTS>
                <RESULT eventid="1178" points="327" reactiontime="+77" swimtime="00:02:39.09" resultid="2785" heatid="5818" lane="6" entrytime="00:02:40.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:02:00.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="327" reactiontime="+79" swimtime="00:01:11.48" resultid="2786" heatid="5889" lane="5" entrytime="00:01:11.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="335" reactiontime="+85" swimtime="00:02:52.87" resultid="2787" heatid="5948" lane="4" entrytime="00:02:59.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:22.98" />
                    <SPLIT distance="150" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="5508" name="Energoatom Varash">
          <ATHLETES>
            <ATHLETE firstname="Anastasiia" lastname="Zaichyk" birthdate="1989-01-01" gender="F" nation="UKR" athleteid="5507">
              <RESULTS>
                <RESULT eventid="1161" points="280" reactiontime="+96" swimtime="00:03:06.13" resultid="5509" heatid="5813" lane="6" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="169" reactiontime="+94" swimtime="00:03:36.19" resultid="5510" heatid="5895" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:37.83" />
                    <SPLIT distance="150" swimtime="00:02:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="223" swimtime="00:03:15.95" resultid="5511" heatid="5902" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="5512" heatid="5919" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3209" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Seweryński" birthdate="1961-01-01" gender="M" nation="POL" athleteid="3208">
              <RESULTS>
                <RESULT eventid="1076" points="211" reactiontime="+108" swimtime="00:00:36.49" resultid="3210" heatid="5775" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1110" points="194" reactiontime="+105" swimtime="00:01:35.45" resultid="3211" heatid="5791" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="220" reactiontime="+103" swimtime="00:00:41.82" resultid="3212" heatid="5869" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1333" points="164" reactiontime="+100" swimtime="00:01:29.91" resultid="3213" heatid="5886" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="219" reactiontime="+107" swimtime="00:00:33.40" resultid="3214" heatid="5930" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1571" points="139" reactiontime="+103" swimtime="00:01:32.12" resultid="3215" heatid="5966" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5513" name="iSwim Białystok">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Markowski" birthdate="1977-09-21" gender="M" nation="POL" athleteid="5559">
              <RESULTS>
                <RESULT eventid="1212" points="194" reactiontime="+95" swimtime="00:02:51.38" resultid="5560" heatid="5831" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:18.65" />
                    <SPLIT distance="150" swimtime="00:02:04.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="204" reactiontime="+88" swimtime="00:01:16.24" resultid="5561" heatid="5851" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="201" reactiontime="+89" swimtime="00:00:34.39" resultid="5562" heatid="5930" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Bocheń" birthdate="1999-12-29" gender="M" nation="POL" athleteid="5563">
              <RESULTS>
                <RESULT eventid="1076" points="574" reactiontime="+63" swimtime="00:00:26.17" resultid="5651" heatid="5783" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1144" points="501" reactiontime="+64" swimtime="00:00:27.97" resultid="5652" heatid="5811" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1367" points="536" reactiontime="+68" swimtime="00:02:13.18" resultid="5653" heatid="5900" lane="5" entrytime="00:02:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="591" reactiontime="+65" swimtime="00:00:56.92" resultid="5654" heatid="5971" lane="5" entrytime="00:00:56.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="5655" heatid="5984" lane="9" entrytime="00:04:27.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Butkiewicz" birthdate="1989-02-25" gender="F" nation="POL" athleteid="5542">
              <RESULTS>
                <RESULT eventid="1282" status="DNS" swimtime="00:00:00.00" resultid="5761" heatid="5864" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="5762" heatid="5921" lane="7" entrytime="00:00:29.90" />
                <RESULT eventid="1093" status="DNS" swimtime="00:00:00.00" resultid="5763" heatid="5788" lane="5" entrytime="00:01:18.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wienczysław" lastname="Safrończyk" birthdate="1954-08-27" gender="M" nation="POL" athleteid="5567">
              <RESULTS>
                <RESULT eventid="1110" points="102" reactiontime="+141" swimtime="00:01:58.13" resultid="5568" heatid="5790" lane="7" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="89" reactiontime="+124" swimtime="00:00:56.52" resultid="5569" heatid="5867" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1503" points="109" swimtime="00:04:11.52" resultid="5570" heatid="5946" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.65" />
                    <SPLIT distance="100" swimtime="00:02:00.61" />
                    <SPLIT distance="150" swimtime="00:03:06.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Chomicki" birthdate="1975-11-07" gender="M" nation="POL" athleteid="5550">
              <RESULTS>
                <RESULT eventid="1076" points="245" reactiontime="+80" swimtime="00:00:34.75" resultid="5551" heatid="5777" lane="8" entrytime="00:00:33.90" />
                <RESULT eventid="1265" points="220" reactiontime="+77" swimtime="00:01:14.37" resultid="5552" heatid="5850" lane="6" entrytime="00:01:16.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="225" reactiontime="+74" swimtime="00:00:33.14" resultid="5553" heatid="5930" lane="1" entrytime="00:00:32.90" />
                <RESULT eventid="1571" points="173" reactiontime="+82" swimtime="00:01:25.64" resultid="5554" heatid="5967" lane="8" entrytime="00:01:19.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Perkowski" birthdate="1996-06-10" gender="M" nation="POL" athleteid="5537">
              <RESULTS>
                <RESULT eventid="1076" points="545" reactiontime="+64" swimtime="00:00:26.62" resultid="5538" heatid="5783" lane="1" entrytime="00:00:26.20" />
                <RESULT eventid="1265" points="580" reactiontime="+63" swimtime="00:00:53.87" resultid="5539" heatid="5857" lane="1" entrytime="00:00:56.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="521" reactiontime="+62" swimtime="00:00:25.05" resultid="5541" heatid="5939" lane="2" entrytime="00:00:24.90" />
                <RESULT eventid="1571" points="541" swimtime="00:00:58.62" resultid="5650" heatid="5971" lane="7" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Humbla" birthdate="1979-01-24" gender="M" nation="POL" athleteid="5514">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5515" heatid="5781" lane="7" entrytime="00:00:28.20" />
                <RESULT eventid="1299" points="433" swimtime="00:00:33.36" resultid="5516" heatid="5873" lane="9" entrytime="00:00:33.90" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5517" heatid="5890" lane="4" entrytime="00:01:09.00" />
                <RESULT eventid="1469" points="465" reactiontime="+62" swimtime="00:00:26.01" resultid="5518" heatid="5937" lane="2" entrytime="00:00:26.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Iłendo" birthdate="1993-02-09" gender="M" nation="POL" athleteid="5530">
              <RESULTS>
                <RESULT eventid="1144" points="460" reactiontime="+69" swimtime="00:00:28.78" resultid="5531" heatid="5811" lane="7" entrytime="00:00:28.90" />
                <RESULT eventid="1212" points="547" swimtime="00:02:01.44" resultid="5532" heatid="5835" lane="2" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                    <SPLIT distance="100" swimtime="00:00:59.62" />
                    <SPLIT distance="150" swimtime="00:01:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="452" reactiontime="+74" swimtime="00:02:17.56" resultid="5534" heatid="5908" lane="1" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5535" heatid="5939" lane="9" entrytime="00:00:25.10" />
                <RESULT eventid="1537" points="478" reactiontime="+69" swimtime="00:01:01.79" resultid="5536" heatid="5962" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="575" reactiontime="+61" swimtime="00:00:54.04" resultid="5663" heatid="5858" lane="0" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Daszuta" birthdate="1973-03-12" gender="M" nation="POL" athleteid="5525">
              <RESULTS>
                <RESULT eventid="1076" points="399" reactiontime="+76" swimtime="00:00:29.54" resultid="5526" heatid="5781" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1144" points="318" reactiontime="+76" swimtime="00:00:32.53" resultid="5527" heatid="5809" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1299" points="424" swimtime="00:00:33.59" resultid="5528" heatid="5873" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5529" heatid="5936" lane="6" entrytime="00:00:26.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" athleteid="5519">
              <RESULTS>
                <RESULT eventid="1076" points="503" reactiontime="+75" swimtime="00:00:27.34" resultid="5520" heatid="5782" lane="1" entrytime="00:00:27.30" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5521" heatid="5892" lane="8" entrytime="00:01:06.00" />
                <RESULT eventid="1367" points="406" reactiontime="+81" swimtime="00:02:26.11" resultid="5522" heatid="5900" lane="0" entrytime="00:02:25.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="504" reactiontime="+74" swimtime="00:00:25.32" resultid="5523" heatid="5938" lane="1" entrytime="00:00:25.85" />
                <RESULT eventid="1571" points="466" reactiontime="+76" swimtime="00:01:01.60" resultid="5524" heatid="5970" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Markowska" birthdate="1981-03-20" gender="F" nation="POL" athleteid="5555">
              <RESULTS>
                <RESULT eventid="1161" points="165" reactiontime="+97" swimtime="00:03:42.07" resultid="5758" heatid="5813" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                    <SPLIT distance="100" swimtime="00:01:53.53" />
                    <SPLIT distance="150" swimtime="00:02:50.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="5759" heatid="5895" lane="7" entrytime="00:03:45.00" />
                <RESULT eventid="1588" points="190" reactiontime="+97" swimtime="00:06:46.74" resultid="5760" heatid="5973" lane="4" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                    <SPLIT distance="150" swimtime="00:02:22.46" />
                    <SPLIT distance="200" swimtime="00:03:15.67" />
                    <SPLIT distance="250" swimtime="00:04:08.85" />
                    <SPLIT distance="300" swimtime="00:05:01.84" />
                    <SPLIT distance="350" swimtime="00:05:55.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="497" reactiontime="+64" swimtime="00:01:43.20" resultid="5564" heatid="5914" lane="2" entrytime="00:01:43.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="100" swimtime="00:00:50.17" />
                    <SPLIT distance="150" swimtime="00:01:17.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5530" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5519" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="5525" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5514" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" points="493" reactiontime="+71" swimtime="00:01:54.46" resultid="5565" heatid="5989" lane="4" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:01:01.56" />
                    <SPLIT distance="150" swimtime="00:01:28.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5530" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="5519" number="2" reactiontime="+5" />
                    <RELAYPOSITION athleteid="5525" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="5514" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1229" status="DNS" swimtime="00:00:00.00" resultid="5566" heatid="5838" lane="6" entrytime="00:02:07.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5555" number="1" />
                    <RELAYPOSITION athleteid="5542" number="2" />
                    <RELAYPOSITION athleteid="5514" number="3" />
                    <RELAYPOSITION athleteid="5525" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5405" name="niezrzeszony" />
        <CLUB type="CLUB" nation="POL" clubid="4008" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Paszkiewicz" birthdate="1975-01-01" gender="M" nation="POL" athleteid="4007">
              <RESULTS>
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1076" reactiontime="+74" status="DSQ" swimtime="00:00:00.00" resultid="4009" heatid="5775" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1265" points="196" swimtime="00:01:17.33" resultid="4010" heatid="5851" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="144" reactiontime="+81" swimtime="00:01:33.90" resultid="4011" heatid="5886" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="242" reactiontime="+69" swimtime="00:00:32.33" resultid="4012" heatid="5932" lane="8" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" nation="POL" region="10" clubid="4381" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Mańczak" birthdate="1971-11-04" gender="M" nation="POL" license="501910700407" swrid="4186188" athleteid="4382">
              <RESULTS>
                <RESULT eventid="1076" points="333" reactiontime="+77" swimtime="00:00:31.36" resultid="4383" heatid="5779" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1367" points="206" reactiontime="+83" swimtime="00:03:03.03" resultid="4384" heatid="5898" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="341" reactiontime="+72" swimtime="00:00:28.85" resultid="4385" heatid="5933" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1571" points="272" reactiontime="+76" swimtime="00:01:13.69" resultid="4386" heatid="5967" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2789" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Gruca" birthdate="2000-01-01" gender="F" nation="POL" swrid="4647670" athleteid="2788">
              <RESULTS>
                <RESULT eventid="1093" points="434" reactiontime="+68" swimtime="00:01:22.32" resultid="2790" heatid="5788" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="407" reactiontime="+75" swimtime="00:00:38.51" resultid="2791" heatid="5863" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1316" points="400" reactiontime="+71" swimtime="00:01:16.69" resultid="2792" heatid="5879" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="4517" name="Masters Avia Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" swrid="5439542" athleteid="4526">
              <RESULTS>
                <RESULT eventid="1076" points="354" reactiontime="+81" swimtime="00:00:30.73" resultid="4527" heatid="5777" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1144" points="334" reactiontime="+75" swimtime="00:00:32.02" resultid="4528" heatid="5809" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1333" points="362" reactiontime="+76" swimtime="00:01:09.11" resultid="4529" heatid="5889" lane="4" entrytime="00:01:11.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="393" swimtime="00:00:27.51" resultid="4530" heatid="5934" lane="9" entrytime="00:00:28.30" />
                <RESULT eventid="1537" points="326" reactiontime="+74" swimtime="00:01:10.22" resultid="4531" heatid="5960" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mazur" birthdate="1995-03-13" gender="M" nation="POL" license="104303700009" swrid="4195380" athleteid="4521">
              <RESULTS>
                <RESULT eventid="1076" points="547" reactiontime="+61" swimtime="00:00:26.59" resultid="4522" heatid="5781" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1265" points="607" reactiontime="+66" swimtime="00:00:53.06" resultid="4523" heatid="5857" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="479" reactiontime="+68" swimtime="00:01:02.97" resultid="4524" heatid="5893" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="566" reactiontime="+59" swimtime="00:00:24.37" resultid="4525" heatid="5939" lane="8" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="4518">
              <RESULTS>
                <RESULT eventid="1076" points="248" reactiontime="+77" swimtime="00:00:34.60" resultid="4519" heatid="5777" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1469" points="293" reactiontime="+87" swimtime="00:00:30.35" resultid="4520" heatid="5932" lane="3" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" swrid="4061691" athleteid="4532">
              <RESULTS>
                <RESULT eventid="1076" points="469" swimtime="00:00:27.99" resultid="4533" heatid="5782" lane="2" entrytime="00:00:27.10" />
                <RESULT eventid="1212" points="517" reactiontime="+76" swimtime="00:02:03.80" resultid="4534" heatid="5834" lane="4" entrytime="00:02:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:00:59.83" />
                    <SPLIT distance="150" swimtime="00:01:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="534" reactiontime="+72" swimtime="00:00:55.37" resultid="4535" heatid="5857" lane="6" entrytime="00:00:55.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="507" reactiontime="+69" swimtime="00:00:25.28" resultid="4536" heatid="5937" lane="8" entrytime="00:00:26.30" />
                <RESULT eventid="1571" points="452" reactiontime="+69" swimtime="00:01:02.22" resultid="4537" heatid="5970" lane="2" entrytime="00:01:03.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="462" reactiontime="+55" swimtime="00:01:45.76" resultid="4538" heatid="5914" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.55" />
                    <SPLIT distance="100" swimtime="00:00:54.25" />
                    <SPLIT distance="150" swimtime="00:01:20.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4521" number="1" reactiontime="+55" />
                    <RELAYPOSITION athleteid="4518" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4526" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4532" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="441" reactiontime="+66" swimtime="00:01:58.73" resultid="4539" heatid="5988" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:29.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4526" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="4532" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4521" number="3" reactiontime="+1" />
                    <RELAYPOSITION athleteid="4518" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="4990" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Walkowicz" birthdate="1978-10-04" gender="M" nation="POL" license="512914700048" athleteid="5055">
              <RESULTS>
                <RESULT eventid="1299" points="253" reactiontime="+71" swimtime="00:00:39.91" resultid="5056" heatid="5871" lane="6" entrytime="00:00:36.99" />
                <RESULT eventid="1469" points="222" reactiontime="+70" swimtime="00:00:33.28" resultid="5057" heatid="5931" lane="8" entrytime="00:00:31.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="5035">
              <RESULTS>
                <RESULT eventid="1144" points="146" reactiontime="+70" swimtime="00:00:42.18" resultid="5036" heatid="5803" lane="3" />
                <RESULT eventid="1212" points="210" reactiontime="+96" swimtime="00:02:47.00" resultid="5037" heatid="5831" lane="7" entrytime="00:02:49.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:20.07" />
                    <SPLIT distance="150" swimtime="00:02:04.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="210" swimtime="00:01:15.51" resultid="5038" heatid="5850" lane="7" entrytime="00:01:17.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="146" reactiontime="+69" swimtime="00:03:20.23" resultid="5039" heatid="5905" lane="3" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="139" reactiontime="+68" swimtime="00:01:33.16" resultid="5040" heatid="5956" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="198" reactiontime="+104" swimtime="00:06:04.00" resultid="5041" heatid="5979" lane="6" entrytime="00:06:10.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                    <SPLIT distance="150" swimtime="00:02:13.86" />
                    <SPLIT distance="200" swimtime="00:03:01.46" />
                    <SPLIT distance="250" swimtime="00:03:48.46" />
                    <SPLIT distance="300" swimtime="00:04:35.51" />
                    <SPLIT distance="350" swimtime="00:05:22.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" swrid="5471789" athleteid="5004">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5005" heatid="5780" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="5006" heatid="5819" lane="8" entrytime="00:02:37.00" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="5007" heatid="5871" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="5008" heatid="5907" lane="6" entrytime="00:02:30.50" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5009" heatid="5934" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5010" heatid="5969" lane="3" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" license="512914600004" swrid="5240932" athleteid="5011">
              <RESULTS>
                <RESULT eventid="1093" points="382" reactiontime="+86" swimtime="00:01:25.89" resultid="5012" heatid="5784" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="432" reactiontime="+76" swimtime="00:00:33.86" resultid="5013" heatid="5801" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1282" points="380" reactiontime="+80" swimtime="00:00:39.43" resultid="5014" heatid="5860" lane="2" />
                <RESULT eventid="1316" points="417" reactiontime="+83" swimtime="00:01:15.59" resultid="5015" heatid="5879" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="5016" heatid="5916" lane="5" />
                <RESULT eventid="1520" status="DNS" swimtime="00:00:00.00" resultid="5017" heatid="5954" lane="2" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" license="512914700009" swrid="4992964" athleteid="5023">
              <RESULTS>
                <RESULT eventid="1110" points="339" reactiontime="+80" swimtime="00:01:19.36" resultid="5024" heatid="5794" lane="0" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="338" reactiontime="+75" swimtime="00:02:22.62" resultid="5025" heatid="5833" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="337" swimtime="00:00:36.26" resultid="5026" heatid="5871" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1503" points="287" reactiontime="+80" swimtime="00:03:02.08" resultid="5027" heatid="5948" lane="8" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="310" reactiontime="+77" swimtime="00:05:13.28" resultid="5028" heatid="5981" lane="3" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:55.28" />
                    <SPLIT distance="200" swimtime="00:02:35.37" />
                    <SPLIT distance="250" swimtime="00:03:15.45" />
                    <SPLIT distance="300" swimtime="00:03:55.79" />
                    <SPLIT distance="350" swimtime="00:04:35.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="5029">
              <RESULTS>
                <RESULT eventid="1110" points="397" reactiontime="+78" swimtime="00:01:15.29" resultid="5030" heatid="5792" lane="0" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1299" points="432" reactiontime="+73" swimtime="00:00:33.38" resultid="5031" heatid="5872" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1333" points="356" reactiontime="+77" swimtime="00:01:09.52" resultid="5032" heatid="5891" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="380" reactiontime="+88" swimtime="00:00:27.81" resultid="5033" heatid="5924" lane="5" />
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="5034" heatid="5950" lane="9" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" swrid="5312396" athleteid="5042">
              <RESULTS>
                <RESULT eventid="1144" points="287" reactiontime="+65" swimtime="00:00:33.67" resultid="5043" heatid="5809" lane="1" entrytime="00:00:32.45" entrycourse="SCM" />
                <RESULT eventid="1178" points="338" swimtime="00:02:37.27" resultid="5044" heatid="5818" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="274" swimtime="00:01:15.86" resultid="5045" heatid="5889" lane="2" entrytime="00:01:12.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="315" reactiontime="+73" swimtime="00:02:35.23" resultid="5046" heatid="5907" lane="3" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="150" swimtime="00:01:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="286" reactiontime="+76" swimtime="00:01:13.34" resultid="5047" heatid="5961" lane="1" entrytime="00:01:11.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="309" reactiontime="+85" swimtime="00:05:13.80" resultid="5048" heatid="5980" lane="5" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:52.69" />
                    <SPLIT distance="200" swimtime="00:02:32.79" />
                    <SPLIT distance="250" swimtime="00:03:13.65" />
                    <SPLIT distance="300" swimtime="00:03:53.47" />
                    <SPLIT distance="350" swimtime="00:04:33.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" swrid="5416809" athleteid="4998">
              <RESULTS>
                <RESULT eventid="1076" points="267" reactiontime="+80" swimtime="00:00:33.75" resultid="4999" heatid="5776" lane="0" entrytime="00:00:36.18" entrycourse="SCM" />
                <RESULT eventid="1212" points="284" reactiontime="+91" swimtime="00:02:31.14" resultid="5000" heatid="5827" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:52.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="297" reactiontime="+77" swimtime="00:01:07.30" resultid="5001" heatid="5846" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="258" reactiontime="+77" swimtime="00:00:39.66" resultid="5002" heatid="5865" lane="5" />
                <RESULT eventid="1469" points="286" reactiontime="+82" swimtime="00:00:30.57" resultid="5003" heatid="5930" lane="6" entrytime="00:00:32.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Fluder" birthdate="1986-03-01" gender="M" nation="POL" license="512914700007" swrid="4073249" athleteid="5049">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1212" points="568" reactiontime="+80" swimtime="00:01:59.98" resultid="5050" heatid="5835" lane="3" entrytime="00:02:00.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:00:58.67" />
                    <SPLIT distance="150" swimtime="00:01:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="538" reactiontime="+76" swimtime="00:00:55.25" resultid="5051" heatid="5858" lane="8" entrytime="00:00:54.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="387" reactiontime="+84" swimtime="00:02:28.41" resultid="5052" heatid="5900" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="482" reactiontime="+74" swimtime="00:00:25.70" resultid="5053" heatid="5938" lane="6" entrytime="00:00:25.46" />
                <RESULT eventid="1605" points="535" swimtime="00:04:21.42" resultid="5054" heatid="5984" lane="7" entrytime="00:04:19.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="100" swimtime="00:01:03.83" />
                    <SPLIT distance="150" swimtime="00:01:37.35" />
                    <SPLIT distance="200" swimtime="00:02:11.53" />
                    <SPLIT distance="250" swimtime="00:02:44.95" />
                    <SPLIT distance="300" swimtime="00:03:18.38" />
                    <SPLIT distance="350" swimtime="00:03:51.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Rowiński" birthdate="1990-07-12" gender="M" nation="POL" license="512914700005" swrid="4060623" athleteid="5018">
              <RESULTS>
                <RESULT eventid="1110" points="531" reactiontime="+68" swimtime="00:01:08.32" resultid="5019" heatid="5796" lane="3" entrytime="00:01:04.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="636" swimtime="00:00:29.36" resultid="5020" heatid="5874" lane="2" entrytime="00:00:29.87" entrycourse="SCM" />
                <RESULT eventid="1333" points="458" swimtime="00:01:03.93" resultid="5021" heatid="5893" lane="7" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5022" heatid="5971" lane="1" entrytime="00:00:59.00" />
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="5064" heatid="5820" lane="7" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" swrid="4043251" athleteid="4991">
              <RESULTS>
                <RESULT eventid="1076" points="625" reactiontime="+78" swimtime="00:00:25.43" resultid="4992" heatid="5783" lane="3" entrytime="00:00:25.25" />
                <RESULT eventid="1144" points="566" reactiontime="+65" swimtime="00:00:26.86" resultid="4993" heatid="5811" lane="4" entrytime="00:00:26.26" />
                <RESULT eventid="1265" points="581" reactiontime="+74" swimtime="00:00:53.84" resultid="4994" heatid="5858" lane="2" entrytime="00:00:53.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4995" heatid="5908" lane="3" entrytime="00:02:09.99" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4996" heatid="5940" lane="0" entrytime="00:00:24.24" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4997" heatid="5984" lane="1" entrytime="00:04:19.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Kaczyński" birthdate="1986-01-16" gender="M" nation="POL" license="112914700016" swrid="4060699" athleteid="5058">
              <RESULTS>
                <RESULT eventid="1469" points="507" reactiontime="+71" swimtime="00:00:25.27" resultid="5059" heatid="5940" lane="8" entrytime="00:00:24.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="553" reactiontime="+68" swimtime="00:01:39.63" resultid="5060" heatid="5914" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.97" />
                    <SPLIT distance="100" swimtime="00:00:50.34" />
                    <SPLIT distance="150" swimtime="00:01:15.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5058" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="5018" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="5049" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4991" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1646" points="541" reactiontime="+63" swimtime="00:01:50.93" resultid="5062" heatid="5989" lane="3" entrytime="00:01:54.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="150" swimtime="00:01:25.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4991" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="5029" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="5058" number="3" reactiontime="+8" />
                    <RELAYPOSITION athleteid="5049" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="335" reactiontime="+72" swimtime="00:01:57.74" resultid="5061" heatid="5914" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:00:59.40" />
                    <SPLIT distance="150" swimtime="00:01:29.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4998" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="5023" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="5042" number="3" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5029" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" points="253" reactiontime="+69" swimtime="00:02:22.81" resultid="5063" heatid="5988" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:01:18.65" />
                    <SPLIT distance="150" swimtime="00:01:52.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5035" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5023" number="2" reactiontime="-1" />
                    <RELAYPOSITION athleteid="5042" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4998" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03302" nation="POL" region="02" clubid="5415" name="TMKS Champions">
          <ATHLETES>
            <ATHLETE firstname="Kazimierz" lastname="Piotrowski" birthdate="1952-12-22" gender="M" nation="POL" athleteid="5416">
              <RESULTS>
                <RESULT eventid="1299" points="93" reactiontime="+99" swimtime="00:00:55.73" resultid="5417" heatid="5867" lane="0" entrytime="00:00:55.55" entrycourse="SCM" />
                <RESULT eventid="1469" points="97" reactiontime="+96" swimtime="00:00:43.75" resultid="5418" heatid="5926" lane="8" entrytime="00:00:42.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3014" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Wiesław" lastname="Majcher" birthdate="1950-01-01" gender="M" nation="POL" swrid="5240919" athleteid="3013">
              <RESULTS>
                <RESULT eventid="1110" points="41" reactiontime="+116" swimtime="00:02:40.13" resultid="3015" heatid="5789" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="33" reactiontime="+107" swimtime="00:05:07.50" resultid="3016" heatid="5827" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="100" swimtime="00:02:19.59" />
                    <SPLIT distance="150" swimtime="00:03:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1265" status="DSQ" swimtime="00:00:00.00" resultid="3017" heatid="5847" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="38" swimtime="00:01:14.86" resultid="3018" heatid="5866" lane="7" />
                <RESULT eventid="1469" points="47" reactiontime="+96" swimtime="00:00:55.86" resultid="3019" heatid="5924" lane="2" />
                <RESULT eventid="1503" points="36" reactiontime="+109" swimtime="00:06:00.77" resultid="3020" heatid="5945" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.34" />
                    <SPLIT distance="100" swimtime="00:02:54.52" />
                    <SPLIT distance="150" swimtime="00:04:29.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="5447" name="Swim Masters Zlin">
          <ATHLETES>
            <ATHLETE firstname="Karel" lastname="Steker" birthdate="1981-08-12" gender="M" nation="CZE" athleteid="5448">
              <RESULTS>
                <RESULT eventid="1076" points="323" reactiontime="+79" swimtime="00:00:31.67" resultid="5449" heatid="5778" lane="5" entrytime="00:00:31.32" />
                <RESULT eventid="1144" points="235" reactiontime="+73" swimtime="00:00:35.97" resultid="5450" heatid="5807" lane="3" entrytime="00:00:35.02" />
                <RESULT eventid="1212" points="337" reactiontime="+77" swimtime="00:02:22.77" resultid="5451" heatid="5833" lane="6" entrytime="00:02:20.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="262" reactiontime="+76" swimtime="00:00:39.46" resultid="5452" heatid="5869" lane="2" entrytime="00:00:40.35" />
                <RESULT eventid="1333" points="286" reactiontime="+72" swimtime="00:01:14.79" resultid="5453" heatid="5889" lane="1" entrytime="00:01:13.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="324" reactiontime="+76" swimtime="00:00:29.33" resultid="5454" heatid="5933" lane="3" entrytime="00:00:28.52" />
                <RESULT eventid="1571" points="303" reactiontime="+74" swimtime="00:01:11.11" resultid="5455" heatid="5968" lane="1" entrytime="00:01:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ivo" lastname="Urban" birthdate="1963-04-27" gender="M" nation="CZE" athleteid="5460">
              <RESULTS>
                <RESULT eventid="1076" points="281" swimtime="00:00:33.19" resultid="5461" heatid="5778" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1144" points="222" reactiontime="+83" swimtime="00:00:36.65" resultid="5462" heatid="5805" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1469" points="338" reactiontime="+80" swimtime="00:00:28.92" resultid="5463" heatid="5931" lane="4" entrytime="00:00:30.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michal" lastname="Prilucik" birthdate="1966-09-28" gender="M" nation="CZE" athleteid="5456">
              <RESULTS>
                <RESULT eventid="1144" points="136" reactiontime="+69" swimtime="00:00:43.20" resultid="5457" heatid="5805" lane="2" entrytime="00:00:43.50" />
                <RESULT eventid="1265" points="193" reactiontime="+85" swimtime="00:01:17.73" resultid="5458" heatid="5850" lane="3" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="208" reactiontime="+75" swimtime="00:00:33.99" resultid="5459" heatid="5929" lane="6" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2849" name="Motyl MOSiR Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" license="100908700263" swrid="4791744" athleteid="2850">
              <RESULTS>
                <RESULT eventid="1076" points="470" reactiontime="+71" swimtime="00:00:27.97" resultid="2851" heatid="5782" lane="0" entrytime="00:00:27.79" />
                <RESULT eventid="1178" points="467" reactiontime="+68" swimtime="00:02:21.29" resultid="2852" heatid="5820" lane="8" entrytime="00:02:21.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="450" reactiontime="+83" swimtime="00:00:58.63" resultid="2853" heatid="5857" lane="0" entrytime="00:00:57.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="445" reactiontime="+73" swimtime="00:01:04.54" resultid="2854" heatid="5892" lane="2" entrytime="00:01:03.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="444" reactiontime="+72" swimtime="00:00:26.41" resultid="2855" heatid="5937" lane="6" entrytime="00:00:26.09" />
                <RESULT eventid="1571" points="458" reactiontime="+73" swimtime="00:01:01.98" resultid="2856" heatid="5970" lane="3" entrytime="00:01:01.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" license="100908600388" swrid="4992840" athleteid="2857">
              <RESULTS>
                <RESULT eventid="1093" points="237" reactiontime="+82" swimtime="00:01:40.72" resultid="2858" heatid="5786" lane="4" entrytime="00:01:44.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="228" swimtime="00:03:19.41" resultid="2859" heatid="5813" lane="5" entrytime="00:03:14.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:36.85" />
                    <SPLIT distance="150" swimtime="00:02:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="229" reactiontime="+90" swimtime="00:00:46.67" resultid="2860" heatid="5862" lane="1" entrytime="00:00:48.99" />
                <RESULT eventid="1316" points="249" swimtime="00:01:29.73" resultid="2861" heatid="5878" lane="7" entrytime="00:01:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="271" reactiontime="+79" swimtime="00:00:35.43" resultid="2862" heatid="5918" lane="2" entrytime="00:00:37.99" />
                <RESULT eventid="1486" points="230" reactiontime="+91" swimtime="00:03:39.38" resultid="2863" heatid="5943" lane="5" entrytime="00:03:39.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                    <SPLIT distance="100" swimtime="00:01:47.50" />
                    <SPLIT distance="150" swimtime="00:02:44.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UKSSPARTA" nation="POL" clubid="2808" name="UKS Sparta Grodzisk Mazowiecki">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Głowa" birthdate="1979-10-08" gender="M" nation="POL" athleteid="2828">
              <RESULTS>
                <RESULT eventid="1076" points="379" reactiontime="+76" swimtime="00:00:30.04" resultid="2829" heatid="5778" lane="1" entrytime="00:00:32.05" entrycourse="SCM" />
                <RESULT eventid="1265" points="394" reactiontime="+89" swimtime="00:01:01.25" resultid="2830" heatid="5854" lane="8" entrytime="00:01:03.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="407" swimtime="00:00:27.20" resultid="2831" heatid="5935" lane="7" entrytime="00:00:27.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Zieliński" birthdate="1980-05-18" gender="M" nation="POL" athleteid="2822">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2823" heatid="5772" lane="5" />
                <RESULT eventid="1110" points="345" reactiontime="+85" swimtime="00:01:18.88" resultid="2824" heatid="5794" lane="1" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="373" reactiontime="+92" swimtime="00:00:35.05" resultid="2825" heatid="5865" lane="4" />
                <RESULT eventid="1333" points="313" swimtime="00:01:12.55" resultid="2826" heatid="5889" lane="7" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="335" reactiontime="+86" swimtime="00:02:52.90" resultid="2827" heatid="5949" lane="5" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:21.01" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Plich" birthdate="1978-06-21" gender="M" nation="POL" athleteid="2809">
              <RESULTS>
                <RESULT eventid="1076" points="331" reactiontime="+78" swimtime="00:00:31.43" resultid="2810" heatid="5778" lane="8" entrytime="00:00:32.05" entrycourse="SCM" />
                <RESULT eventid="1144" points="264" reactiontime="+84" swimtime="00:00:34.63" resultid="2811" heatid="5808" lane="4" entrytime="00:00:33.08" entrycourse="SCM" />
                <RESULT eventid="1333" points="284" reactiontime="+78" swimtime="00:01:14.90" resultid="2812" heatid="5888" lane="1" entrytime="00:01:17.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="278" reactiontime="+82" swimtime="00:01:14.00" resultid="2813" heatid="5961" lane="2" entrytime="00:01:10.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Rzewuska" birthdate="1997-05-30" gender="F" nation="POL" swrid="4261695" athleteid="2814">
              <RESULTS>
                <RESULT eventid="1127" points="464" reactiontime="+65" swimtime="00:00:33.05" resultid="2815" heatid="5802" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1384" points="426" reactiontime="+68" swimtime="00:02:38.05" resultid="2816" heatid="5903" lane="3" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="427" reactiontime="+66" swimtime="00:01:12.88" resultid="2817" heatid="5955" lane="3" entrytime="00:01:08.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Milewski" birthdate="1992-03-04" gender="M" nation="POL" swrid="4124793" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1076" points="422" swimtime="00:00:28.99" resultid="2819" heatid="5781" lane="2" entrytime="00:00:28.05" entrycourse="SCM" />
                <RESULT eventid="1265" points="441" reactiontime="+74" swimtime="00:00:59.01" resultid="2820" heatid="5857" lane="5" entrytime="00:00:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="440" reactiontime="+86" swimtime="00:00:26.49" resultid="2821" heatid="5939" lane="0" entrytime="00:00:25.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="417" swimtime="00:01:49.47" resultid="2833" heatid="5914" lane="9" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                    <SPLIT distance="150" swimtime="00:01:21.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2818" number="1" />
                    <RELAYPOSITION athleteid="2828" number="2" />
                    <RELAYPOSITION athleteid="2822" number="3" />
                    <RELAYPOSITION athleteid="2809" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="UKS Sparta Grodzisk Mayowiecki" number="1">
              <RESULTS>
                <RESULT eventid="1646" points="372" reactiontime="+75" swimtime="00:02:05.65" resultid="2832" heatid="5989" lane="1" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:38.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2809" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="2822" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2828" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="2818" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3335" name="MOSiR Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" swrid="4216999" athleteid="3336">
              <RESULTS>
                <RESULT eventid="1076" points="150" reactiontime="+79" swimtime="00:00:40.91" resultid="3337" heatid="5774" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1110" points="102" reactiontime="+85" swimtime="00:01:58.08" resultid="3338" heatid="5790" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="145" reactiontime="+99" swimtime="00:00:48.06" resultid="3339" heatid="5867" lane="6" entrytime="00:00:49.50" />
                <RESULT eventid="1333" points="112" reactiontime="+92" swimtime="00:01:42.08" resultid="3340" heatid="5883" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="164" swimtime="00:00:36.78" resultid="3341" heatid="5928" lane="9" entrytime="00:00:36.50" />
                <RESULT eventid="1571" points="76" reactiontime="+101" swimtime="00:01:52.79" resultid="3342" heatid="5966" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5287" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Lelewski" birthdate="1965-01-01" gender="M" nation="POL" athleteid="5286">
              <RESULTS>
                <RESULT eventid="1503" points="229" swimtime="00:03:16.31" resultid="5288" heatid="5947" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="150" swimtime="00:02:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="251" reactiontime="+85" swimtime="00:05:36.33" resultid="5289" heatid="5980" lane="2" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                    <SPLIT distance="150" swimtime="00:02:02.39" />
                    <SPLIT distance="200" swimtime="00:02:45.45" />
                    <SPLIT distance="250" swimtime="00:03:28.89" />
                    <SPLIT distance="300" swimtime="00:04:11.97" />
                    <SPLIT distance="350" swimtime="00:04:55.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="4600" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Sergiusz" lastname="Olejniczak" birthdate="1978-12-01" gender="M" nation="POL" license="502805700058" athleteid="4682">
              <RESULTS>
                <RESULT eventid="1110" points="359" reactiontime="+74" swimtime="00:01:17.80" resultid="4683" heatid="5795" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="347" reactiontime="+73" swimtime="00:02:35.92" resultid="4684" heatid="5819" lane="0" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="359" reactiontime="+65" swimtime="00:01:09.28" resultid="4685" heatid="5891" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="263" reactiontime="+68" swimtime="00:02:48.78" resultid="4686" heatid="5899" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="353" reactiontime="+76" swimtime="00:02:50.00" resultid="4687" heatid="5949" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:21.23" />
                    <SPLIT distance="150" swimtime="00:02:06.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="331" reactiontime="+69" swimtime="00:05:06.78" resultid="4688" heatid="5982" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:48.68" />
                    <SPLIT distance="200" swimtime="00:02:27.41" />
                    <SPLIT distance="250" swimtime="00:03:06.59" />
                    <SPLIT distance="300" swimtime="00:03:47.06" />
                    <SPLIT distance="350" swimtime="00:04:27.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Szalbierz" birthdate="1968-08-06" gender="M" nation="POL" license="502805700034" swrid="5373990" athleteid="4627">
              <RESULTS>
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1076" reactiontime="+103" status="DSQ" swimtime="00:00:00.00" resultid="4628" heatid="5776" lane="5" entrytime="00:00:34.23" entrycourse="SCM" />
                <RESULT eventid="1333" points="202" reactiontime="+108" swimtime="00:01:23.87" resultid="4629" heatid="5887" lane="8" entrytime="00:01:22.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="265" reactiontime="+101" swimtime="00:00:31.38" resultid="4630" heatid="5931" lane="6" entrytime="00:00:30.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Niedźwiedź" birthdate="1963-07-18" gender="M" nation="POL" license="502805700023" swrid="4754661" athleteid="4722">
              <RESULTS>
                <RESULT eventid="1367" points="77" reactiontime="+84" swimtime="00:04:13.96" resultid="4723" heatid="5897" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.46" />
                    <SPLIT distance="100" swimtime="00:02:00.08" />
                    <SPLIT distance="150" swimtime="00:03:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4724" heatid="5904" lane="4" entrytime="00:04:00.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="4725" heatid="5958" lane="9" entrytime="00:02:00.00" />
                <RESULT eventid="1571" points="83" reactiontime="+111" swimtime="00:01:49.50" resultid="4726" heatid="5965" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="4661">
              <RESULTS>
                <RESULT eventid="1110" points="147" reactiontime="+95" swimtime="00:01:44.70" resultid="4662" heatid="5790" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="206" swimtime="00:00:42.70" resultid="4663" heatid="5868" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="1503" points="117" reactiontime="+104" swimtime="00:04:04.99" resultid="4664" heatid="5946" lane="3" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:51.26" />
                    <SPLIT distance="150" swimtime="00:02:56.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Łatecki" birthdate="1957-05-25" gender="M" nation="POL" license="502805700022" swrid="5464093" athleteid="4693">
              <RESULTS>
                <RESULT eventid="1178" points="40" reactiontime="+105" swimtime="00:05:19.40" resultid="4694" heatid="5816" lane="1" entrytime="00:04:05.00" />
                <RESULT eventid="1401" points="25" reactiontime="+96" swimtime="00:05:59.08" resultid="4695" heatid="5904" lane="5" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.78" />
                    <SPLIT distance="100" swimtime="00:02:53.38" />
                    <SPLIT distance="150" swimtime="00:04:25.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="65" reactiontime="+115" swimtime="00:08:47.68" resultid="4696" heatid="5977" lane="4" entrytime="00:08:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.26" />
                    <SPLIT distance="100" swimtime="00:02:01.67" />
                    <SPLIT distance="150" swimtime="00:03:09.07" />
                    <SPLIT distance="200" swimtime="00:04:17.49" />
                    <SPLIT distance="250" swimtime="00:06:34.34" />
                    <SPLIT distance="300" swimtime="00:07:42.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="4620">
              <RESULTS>
                <RESULT eventid="1076" points="243" reactiontime="+87" swimtime="00:00:34.85" resultid="4621" heatid="5777" lane="1" entrytime="00:00:33.61" entrycourse="SCM" />
                <RESULT eventid="1212" points="234" reactiontime="+88" swimtime="00:02:41.15" resultid="4622" heatid="5831" lane="6" entrytime="00:02:45.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="263" reactiontime="+88" swimtime="00:01:10.13" resultid="4623" heatid="5851" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4624" heatid="5906" lane="8" entrytime="00:03:07.00" />
                <RESULT eventid="1469" points="251" reactiontime="+88" swimtime="00:00:31.92" resultid="4625" heatid="5931" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="4626" heatid="5959" lane="2" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Sztyler" birthdate="1994-11-29" gender="M" nation="POL" license="502805700060" swrid="4227130" athleteid="4658">
              <RESULTS>
                <RESULT eventid="1110" points="556" reactiontime="+61" swimtime="00:01:07.26" resultid="4659" heatid="5796" lane="2" entrytime="00:01:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="573" reactiontime="+61" swimtime="00:00:30.39" resultid="4660" heatid="5874" lane="6" entrytime="00:00:29.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="4639">
              <RESULTS>
                <RESULT eventid="1093" points="254" reactiontime="+66" swimtime="00:01:38.42" resultid="4640" heatid="5787" lane="7" entrytime="00:01:39.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="191" reactiontime="+83" swimtime="00:00:44.40" resultid="4641" heatid="5799" lane="3" entrytime="00:00:44.92" />
                <RESULT eventid="1282" points="256" reactiontime="+71" swimtime="00:00:44.96" resultid="4642" heatid="5862" lane="5" entrytime="00:00:45.47" entrycourse="SCM" />
                <RESULT eventid="1316" points="190" reactiontime="+76" swimtime="00:01:38.14" resultid="4643" heatid="5877" lane="5" entrytime="00:01:39.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="233" reactiontime="+74" swimtime="00:03:38.61" resultid="4644" heatid="5943" lane="6" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.80" />
                    <SPLIT distance="100" swimtime="00:01:47.58" />
                    <SPLIT distance="150" swimtime="00:02:45.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Maciejewski" birthdate="1974-04-11" gender="M" nation="POL" license="502805700028" swrid="5373991" athleteid="4671">
              <RESULTS>
                <RESULT eventid="1110" status="DNS" swimtime="00:00:00.00" resultid="4672" heatid="5791" lane="7" entrytime="00:01:38.00" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="4673" heatid="5851" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="4674" heatid="5868" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4675" heatid="5933" lane="7" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Strójwąs" birthdate="1998-06-29" gender="F" nation="POL" license="502805600061" athleteid="4719">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1451" reactiontime="+60" status="DSQ" swimtime="00:00:00.00" resultid="4721" heatid="5919" lane="4" entrytime="00:00:32.33" />
                <RESULT eventid="1195" points="204" reactiontime="+81" swimtime="00:03:07.55" resultid="5764" heatid="5825" lane="0" entrytime="00:02:31.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:24.05" />
                    <SPLIT distance="150" swimtime="00:02:15.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Jagiełło" birthdate="1979-03-01" gender="M" nation="POL" license="502805700042" swrid="4541616" athleteid="4613">
              <RESULTS>
                <RESULT eventid="1076" points="407" swimtime="00:00:29.34" resultid="4614" heatid="5772" lane="2" />
                <RESULT eventid="1144" points="358" reactiontime="+79" swimtime="00:00:31.28" resultid="4615" heatid="5809" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1299" points="455" reactiontime="+83" swimtime="00:00:32.81" resultid="4616" heatid="5865" lane="3" />
                <RESULT eventid="1333" points="434" reactiontime="+80" swimtime="00:01:05.06" resultid="4617" heatid="5890" lane="3" entrytime="00:01:09.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="451" reactiontime="+76" swimtime="00:00:26.28" resultid="4618" heatid="5935" lane="6" entrytime="00:00:27.02" />
                <RESULT eventid="1537" points="336" reactiontime="+77" swimtime="00:01:09.50" resultid="4619" heatid="5961" lane="7" entrytime="00:01:10.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1984-02-23" gender="F" nation="POL" license="102805600050" athleteid="4704">
              <RESULTS>
                <RESULT eventid="1195" points="245" reactiontime="+85" swimtime="00:02:56.43" resultid="4705" heatid="5823" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="249" reactiontime="+82" swimtime="00:00:45.35" resultid="4706" heatid="5863" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1384" status="DNS" swimtime="00:00:00.00" resultid="4707" heatid="5902" lane="4" entrytime="00:02:55.00" />
                <RESULT eventid="1588" points="259" reactiontime="+83" swimtime="00:06:06.81" resultid="4708" heatid="5973" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:11.39" />
                    <SPLIT distance="200" swimtime="00:02:58.83" />
                    <SPLIT distance="250" swimtime="00:03:46.29" />
                    <SPLIT distance="300" swimtime="00:04:34.22" />
                    <SPLIT distance="350" swimtime="00:05:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1093" points="260" reactiontime="+83" swimtime="00:01:37.68" resultid="5084" heatid="5787" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="263" reactiontime="+88" swimtime="00:03:29.89" resultid="5086" heatid="5944" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:40.77" />
                    <SPLIT distance="150" swimtime="00:02:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gajda" birthdate="1978-02-23" gender="M" nation="POL" license="502805700059" swrid="5272788" athleteid="4676">
              <RESULTS>
                <RESULT eventid="1110" points="225" reactiontime="+86" swimtime="00:01:30.92" resultid="4677" heatid="5792" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="247" reactiontime="+68" swimtime="00:00:35.39" resultid="4678" heatid="5807" lane="2" entrytime="00:00:36.71" entrycourse="SCM" />
                <RESULT eventid="1265" points="241" reactiontime="+83" swimtime="00:01:12.16" resultid="4679" heatid="5851" lane="1" entrytime="00:01:12.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="251" reactiontime="+89" swimtime="00:01:18.09" resultid="4680" heatid="5887" lane="4" entrytime="00:01:19.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="271" reactiontime="+89" swimtime="00:00:31.15" resultid="4681" heatid="5931" lane="5" entrytime="00:00:30.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="4645">
              <RESULTS>
                <RESULT eventid="1110" points="184" reactiontime="+101" swimtime="00:01:37.21" resultid="4646" heatid="5791" lane="3" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="125" reactiontime="+82" swimtime="00:00:44.35" resultid="4647" heatid="5805" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="1299" points="197" swimtime="00:00:43.37" resultid="4648" heatid="5869" lane="9" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1401" points="120" reactiontime="+82" swimtime="00:03:33.81" resultid="4649" heatid="5905" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.12" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="162" reactiontime="+116" swimtime="00:03:40.23" resultid="4650" heatid="5946" lane="5" entrytime="00:03:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.48" />
                    <SPLIT distance="100" swimtime="00:01:47.66" />
                    <SPLIT distance="150" swimtime="00:02:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="120" reactiontime="+91" swimtime="00:01:37.75" resultid="4651" heatid="5958" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="4652">
              <RESULTS>
                <RESULT eventid="1110" points="238" reactiontime="+93" swimtime="00:01:29.22" resultid="4653" heatid="5792" lane="6" entrytime="00:01:29.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="212" reactiontime="+97" swimtime="00:02:46.62" resultid="4654" heatid="5830" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="281" reactiontime="+97" swimtime="00:00:38.55" resultid="4655" heatid="5870" lane="8" entrytime="00:00:38.93" entrycourse="SCM" />
                <RESULT eventid="1503" points="201" swimtime="00:03:25.08" resultid="4656" heatid="5947" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                    <SPLIT distance="150" swimtime="00:02:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="207" reactiontime="+99" swimtime="00:05:58.59" resultid="4657" heatid="5978" lane="4" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:01:49.29" />
                    <SPLIT distance="200" swimtime="00:02:50.19" />
                    <SPLIT distance="250" swimtime="00:03:37.85" />
                    <SPLIT distance="300" swimtime="00:04:25.62" />
                    <SPLIT distance="350" swimtime="00:05:13.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="4665">
              <RESULTS>
                <RESULT eventid="1110" points="172" reactiontime="+101" swimtime="00:01:39.48" resultid="4666" heatid="5791" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="121" reactiontime="+98" swimtime="00:00:44.87" resultid="4667" heatid="5806" lane="6" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1299" points="170" reactiontime="+109" swimtime="00:00:45.56" resultid="4668" heatid="5868" lane="2" entrytime="00:00:44.00" />
                <RESULT eventid="1333" points="149" swimtime="00:01:32.91" resultid="4669" heatid="5885" lane="7" entrytime="00:01:32.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="195" swimtime="00:00:34.76" resultid="4670" heatid="5929" lane="9" entrytime="00:00:34.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="4601">
              <RESULTS>
                <RESULT eventid="1059" points="428" reactiontime="+79" swimtime="00:00:32.35" resultid="4602" heatid="5771" lane="0" entrytime="00:00:32.52" entrycourse="SCM" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas lepszy od Rekordu Polski Kat. F" eventid="1161" points="424" reactiontime="+66" swimtime="00:02:42.15" resultid="4603" heatid="5814" lane="1" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:02:03.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="432" swimtime="00:00:37.78" resultid="4604" heatid="5864" lane="7" entrytime="00:00:38.03" entrycourse="SCM" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1316" points="457" reactiontime="+75" swimtime="00:01:13.36" resultid="4605" heatid="5880" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1554" points="446" reactiontime="+79" swimtime="00:01:11.45" resultid="4606" heatid="5964" lane="3" entrytime="00:01:12.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daria" lastname="Fajkowska" birthdate="1973-03-18" gender="F" nation="POL" license="502805600044" swrid="4992744" athleteid="4689">
              <RESULTS>
                <RESULT eventid="1127" points="408" reactiontime="+80" swimtime="00:00:34.51" resultid="4690" heatid="5802" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1316" points="463" reactiontime="+83" swimtime="00:01:13.01" resultid="4691" heatid="5880" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="390" reactiontime="+73" swimtime="00:01:15.11" resultid="4692" heatid="5955" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Błasiak" birthdate="1955-03-16" gender="M" nation="POL" license="502805700037" swrid="5464088" athleteid="4697">
              <RESULTS>
                <RESULT eventid="1178" points="63" reactiontime="+98" swimtime="00:04:35.17" resultid="4698" heatid="5816" lane="0" entrytime="00:04:24.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.71" />
                    <SPLIT distance="100" swimtime="00:02:19.89" />
                    <SPLIT distance="150" swimtime="00:03:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="87" reactiontime="+89" swimtime="00:03:43.69" resultid="4699" heatid="5828" lane="3" entrytime="00:03:45.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="90" reactiontime="+90" swimtime="00:01:40.27" resultid="4700" heatid="5848" lane="0" entrytime="00:01:42.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="28" reactiontime="+98" swimtime="00:05:55.01" resultid="4701" heatid="5897" lane="0" entrytime="00:05:14.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.06" />
                    <SPLIT distance="100" swimtime="00:02:53.17" />
                    <SPLIT distance="150" swimtime="00:04:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="43" reactiontime="+102" swimtime="00:02:16.95" resultid="4702" heatid="5957" lane="5" entrytime="00:02:09.42" />
                <RESULT eventid="1571" points="25" swimtime="00:02:42.98" resultid="4703" heatid="5965" lane="5" entrytime="00:02:17.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Klusek" birthdate="1975-01-12" gender="F" nation="POL" license="502805600030" swrid="5464092" athleteid="4635">
              <RESULTS>
                <RESULT eventid="1093" points="318" reactiontime="+95" swimtime="00:01:31.28" resultid="4636" heatid="5788" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="243" reactiontime="+99" swimtime="00:03:11.51" resultid="4637" heatid="5895" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:29.06" />
                    <SPLIT distance="150" swimtime="00:02:19.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="268" reactiontime="+98" swimtime="00:01:24.70" resultid="4638" heatid="5964" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="4631">
              <RESULTS>
                <RESULT eventid="1093" points="97" reactiontime="+133" swimtime="00:02:15.46" resultid="4632" heatid="5785" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="86" reactiontime="+125" swimtime="00:01:53.57" resultid="4633" heatid="5841" lane="8" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="91" reactiontime="+121" swimtime="00:01:03.44" resultid="4634" heatid="5861" lane="0" entrytime="00:01:02.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="4607">
              <RESULTS>
                <RESULT eventid="1059" points="309" reactiontime="+83" swimtime="00:00:36.05" resultid="4608" heatid="5770" lane="0" entrytime="00:00:35.04" entrycourse="SCM" />
                <RESULT eventid="1127" points="238" reactiontime="+79" swimtime="00:00:41.28" resultid="4609" heatid="5800" lane="9" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1316" points="277" reactiontime="+92" swimtime="00:01:26.65" resultid="4610" heatid="5879" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="309" reactiontime="+85" swimtime="00:00:33.90" resultid="4611" heatid="5919" lane="6" entrytime="00:00:33.72" entrycourse="SCM" />
                <RESULT eventid="1554" points="205" reactiontime="+95" swimtime="00:01:32.51" resultid="4612" heatid="5964" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-01" gender="F" nation="POL" athleteid="5088">
              <RESULTS>
                <RESULT eventid="1093" points="144" reactiontime="+103" swimtime="00:01:58.71" resultid="5089" heatid="5787" lane="0" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="131" reactiontime="+102" swimtime="00:03:36.92" resultid="5090" heatid="5822" lane="1" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="144" reactiontime="+89" swimtime="00:01:35.81" resultid="5091" heatid="5841" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="146" reactiontime="+101" swimtime="00:00:54.21" resultid="5092" heatid="5863" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1451" points="154" reactiontime="+102" swimtime="00:00:42.72" resultid="5093" heatid="5917" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" swrid="5464087" athleteid="4709">
              <RESULTS>
                <RESULT eventid="1212" points="154" reactiontime="+102" swimtime="00:03:05.38" resultid="4710" heatid="5829" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:26.92" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="127" swimtime="00:01:37.84" resultid="4711" heatid="5885" lane="9" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="50" reactiontime="+103" swimtime="00:00:54.61" resultid="4712" heatid="5928" lane="8" entrytime="00:00:35.80" />
                <RESULT eventid="1605" points="148" reactiontime="+110" swimtime="00:06:41.24" resultid="4713" heatid="5978" lane="2" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:32.92" />
                    <SPLIT distance="150" swimtime="00:02:23.99" />
                    <SPLIT distance="200" swimtime="00:03:16.26" />
                    <SPLIT distance="250" swimtime="00:04:08.26" />
                    <SPLIT distance="300" swimtime="00:04:59.63" />
                    <SPLIT distance="350" swimtime="00:05:50.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Dziarek" birthdate="1959-02-19" gender="M" nation="POL" license="502805700029" swrid="4841500" athleteid="4714">
              <RESULTS>
                <RESULT eventid="1212" points="212" reactiontime="+97" swimtime="00:02:46.55" resultid="4715" heatid="5831" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:03.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="236" swimtime="00:01:12.67" resultid="4716" heatid="5851" lane="9" entrytime="00:01:14.00" />
                <RESULT eventid="1469" points="223" reactiontime="+106" swimtime="00:00:33.20" resultid="4717" heatid="5928" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1605" points="226" reactiontime="+94" swimtime="00:05:48.36" resultid="4718" heatid="5979" lane="3" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:21.61" />
                    <SPLIT distance="150" swimtime="00:02:06.11" />
                    <SPLIT distance="250" swimtime="00:03:36.35" />
                    <SPLIT distance="350" swimtime="00:05:07.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" status="DNF" swimtime="00:00:00.00" resultid="4730" heatid="5913" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4658" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="4682" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="4627" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="4613" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="348" reactiontime="+72" swimtime="00:02:08.51" resultid="4733" heatid="5989" lane="9" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:02.70" />
                    <SPLIT distance="150" swimtime="00:01:38.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4682" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4658" number="2" />
                    <RELAYPOSITION athleteid="4627" number="3" />
                    <RELAYPOSITION athleteid="4676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="219" reactiontime="+95" swimtime="00:02:15.70" resultid="4731" heatid="5912" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:43.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4652" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="4665" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4709" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4620" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="376" swimtime="00:02:08.09" resultid="4729" heatid="5910" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:37.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4601" number="1" />
                    <RELAYPOSITION athleteid="4635" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4607" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4689" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="366" reactiontime="+64" swimtime="00:02:23.01" resultid="4732" heatid="5986" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:48.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4689" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="4635" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4601" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4607" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="268" reactiontime="+78" swimtime="00:02:29.16" resultid="4727" heatid="5837" lane="5" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:01:55.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4607" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4645" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4601" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4620" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="403" reactiontime="+76" swimtime="00:02:10.21" resultid="4728" heatid="5838" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4689" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4658" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4635" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4613" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2763" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-01-01" gender="M" nation="POL" athleteid="2762">
              <RESULTS>
                <RESULT eventid="1076" points="87" reactiontime="+94" swimtime="00:00:48.94" resultid="2764" heatid="5773" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1212" points="101" reactiontime="+105" swimtime="00:03:32.92" resultid="2765" heatid="5828" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:44.29" />
                    <SPLIT distance="150" swimtime="00:02:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="104" reactiontime="+90" swimtime="00:01:35.49" resultid="2766" heatid="5848" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="110" swimtime="00:00:41.96" resultid="2767" heatid="5926" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1605" points="100" reactiontime="+101" swimtime="00:07:36.70" resultid="2768" heatid="5978" lane="0" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                    <SPLIT distance="100" swimtime="00:01:46.57" />
                    <SPLIT distance="150" swimtime="00:02:45.29" />
                    <SPLIT distance="200" swimtime="00:03:43.60" />
                    <SPLIT distance="250" swimtime="00:04:41.94" />
                    <SPLIT distance="300" swimtime="00:05:40.63" />
                    <SPLIT distance="350" swimtime="00:06:40.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5113" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Jawor" birthdate="1976-01-01" gender="M" nation="POL" athleteid="5112">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="5114" heatid="5830" lane="7" entrytime="00:03:00.00" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="5115" heatid="5850" lane="9" entrytime="00:01:19.00" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5116" heatid="5927" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="5117" heatid="5979" lane="1" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2729" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mariusz" lastname="Maciaszek" birthdate="1991-01-01" gender="M" nation="POL" athleteid="2728">
              <RESULTS>
                <RESULT eventid="1076" points="432" reactiontime="+74" swimtime="00:00:28.76" resultid="2730" heatid="5780" lane="1" entrytime="00:00:29.80" />
                <RESULT eventid="1265" points="383" swimtime="00:01:01.84" resultid="2731" heatid="5856" lane="9" entrytime="00:00:59.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="318" reactiontime="+78" swimtime="00:01:12.19" resultid="2732" heatid="5889" lane="3" entrytime="00:01:11.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="439" reactiontime="+76" swimtime="00:00:26.51" resultid="2733" heatid="5937" lane="1" entrytime="00:00:26.26" />
                <RESULT eventid="1571" points="287" reactiontime="+81" swimtime="00:01:12.39" resultid="2734" heatid="5968" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2977" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Edward" lastname="Mężyk" birthdate="1984-01-01" gender="M" nation="POL" swrid="4060389" athleteid="2976">
              <RESULTS>
                <RESULT eventid="1144" points="373" reactiontime="+81" swimtime="00:00:30.85" resultid="2978" heatid="5810" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1265" points="308" swimtime="00:01:06.51" resultid="2979" heatid="5853" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="100111" nation="POL" clubid="2980" name="UKS TRÓJKA Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" swrid="4289072" athleteid="3002">
              <RESULTS>
                <RESULT eventid="1059" points="370" reactiontime="+82" swimtime="00:00:33.94" resultid="3003" heatid="5770" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1195" points="445" reactiontime="+75" swimtime="00:02:24.60" resultid="3004" heatid="5825" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                    <SPLIT distance="150" swimtime="00:01:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="386" reactiontime="+90" swimtime="00:01:08.99" resultid="3005" heatid="5843" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="3006" heatid="5880" lane="6" entrytime="00:01:14.30" />
                <RESULT eventid="1451" points="386" swimtime="00:00:31.49" resultid="3007" heatid="5921" lane="9" entrytime="00:00:30.80" />
                <RESULT eventid="1554" points="391" reactiontime="+84" swimtime="00:01:14.66" resultid="3008" heatid="5964" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" swrid="4602697" athleteid="2988">
              <RESULTS>
                <RESULT eventid="1059" points="554" reactiontime="+77" swimtime="00:00:29.68" resultid="2989" heatid="5771" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1161" points="532" reactiontime="+76" swimtime="00:02:30.38" resultid="2990" heatid="5814" lane="6" entrytime="00:02:35.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="612" reactiontime="+77" swimtime="00:00:59.16" resultid="2991" heatid="5844" lane="5" entrytime="00:00:59.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="576" reactiontime="+76" swimtime="00:01:07.91" resultid="2992" heatid="5881" lane="6" entrytime="00:01:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="625" reactiontime="+74" swimtime="00:00:26.81" resultid="2993" heatid="5922" lane="5" entrytime="00:00:26.74" />
                <RESULT eventid="1554" points="501" reactiontime="+79" swimtime="00:01:08.73" resultid="2994" heatid="5964" lane="5" entrytime="00:01:09.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Chowaniec" birthdate="1995-06-07" gender="M" nation="POL" license="100111700079" swrid="5265087" athleteid="2995">
              <RESULTS>
                <RESULT eventid="1110" points="526" reactiontime="+71" swimtime="00:01:08.52" resultid="2996" heatid="5796" lane="9" entrytime="00:01:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="443" reactiontime="+75" swimtime="00:02:23.79" resultid="2997" heatid="5819" lane="3" entrytime="00:02:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="547" swimtime="00:00:30.87" resultid="2998" heatid="5874" lane="9" entrytime="00:00:31.28" />
                <RESULT eventid="1333" points="466" swimtime="00:01:03.56" resultid="2999" heatid="5892" lane="7" entrytime="00:01:04.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="3000" heatid="5936" lane="3" entrytime="00:00:26.83" />
                <RESULT eventid="1503" points="476" swimtime="00:02:33.85" resultid="3001" heatid="5950" lane="7" entrytime="00:02:39.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:55.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" swrid="4762175" athleteid="2981">
              <RESULTS>
                <RESULT eventid="1076" points="590" reactiontime="+66" swimtime="00:00:25.92" resultid="2982" heatid="5783" lane="7" entrytime="00:00:26.02" />
                <RESULT eventid="1212" points="537" reactiontime="+72" swimtime="00:02:02.20" resultid="2983" heatid="5835" lane="7" entrytime="00:02:02.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="570" reactiontime="+68" swimtime="00:00:54.19" resultid="2984" heatid="5858" lane="1" entrytime="00:00:54.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="483" reactiontime="+68" swimtime="00:01:02.80" resultid="2985" heatid="5892" lane="6" entrytime="00:01:03.45" />
                <RESULT eventid="1469" points="555" reactiontime="+64" swimtime="00:00:24.53" resultid="2986" heatid="5939" lane="4" entrytime="00:00:24.46" />
                <RESULT eventid="1571" points="551" reactiontime="+67" swimtime="00:00:58.27" resultid="2987" heatid="5970" lane="4" entrytime="00:01:00.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5066" name="Litwin Sports">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Drop" birthdate="1966-01-01" gender="F" nation="POL" athleteid="5065">
              <RESULTS>
                <RESULT eventid="1059" points="170" reactiontime="+100" swimtime="00:00:44.00" resultid="5067" heatid="5768" lane="8" entrytime="00:00:55.00" />
                <RESULT eventid="1247" points="189" reactiontime="+95" swimtime="00:01:27.52" resultid="5068" heatid="5841" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="182" reactiontime="+101" swimtime="00:03:14.62" resultid="5069" heatid="5823" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:34.45" />
                    <SPLIT distance="150" swimtime="00:02:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="183" reactiontime="+92" swimtime="00:01:39.47" resultid="5070" heatid="5877" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magda" lastname="Kolasa" birthdate="1991-01-01" gender="F" nation="POL" athleteid="5071">
              <RESULTS>
                <RESULT eventid="1059" points="399" reactiontime="+79" swimtime="00:00:33.10" resultid="5072" heatid="5768" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1247" points="418" reactiontime="+77" swimtime="00:01:07.19" resultid="5073" heatid="5842" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="410" swimtime="00:02:28.61" resultid="5074" heatid="5824" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="387" reactiontime="+75" swimtime="00:01:17.50" resultid="5075" heatid="5878" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Litwin-Żuard" birthdate="1992-01-01" gender="F" nation="POL" athleteid="5079">
              <RESULTS>
                <RESULT eventid="1384" points="443" reactiontime="+75" swimtime="00:02:35.93" resultid="5080" heatid="5903" lane="5" entrytime="00:02:38.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:15.79" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="542" reactiontime="+87" swimtime="00:02:15.39" resultid="5081" heatid="5825" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Krajcarska" birthdate="1994-01-01" gender="F" nation="POL" athleteid="5076">
              <RESULTS>
                <RESULT eventid="1059" points="329" reactiontime="+80" swimtime="00:00:35.30" resultid="5077" heatid="5770" lane="9" entrytime="00:00:36.30" />
                <RESULT eventid="1247" points="292" reactiontime="+78" swimtime="00:01:15.74" resultid="5078" heatid="5842" lane="1" entrytime="00:01:15.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="362" swimtime="00:02:09.68" resultid="5082" heatid="5910" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:41.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5071" number="1" />
                    <RELAYPOSITION athleteid="5065" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="5076" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="5079" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3919" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Kotulski" birthdate="1981-01-01" gender="M" nation="POL" athleteid="3918">
              <RESULTS>
                <RESULT eventid="1265" points="228" reactiontime="+74" swimtime="00:01:13.51" resultid="3920" heatid="5849" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="226" reactiontime="+73" swimtime="00:00:33.07" resultid="3921" heatid="5930" lane="9" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3634" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Królikowski" birthdate="1980-01-01" gender="M" nation="POL" athleteid="3633">
              <RESULTS>
                <RESULT eventid="1537" points="238" reactiontime="+67" swimtime="00:01:17.94" resultid="3635" heatid="5959" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="287" reactiontime="+84" swimtime="00:05:21.68" resultid="3636" heatid="5980" lane="6" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:02:35.48" />
                    <SPLIT distance="250" swimtime="00:03:18.25" />
                    <SPLIT distance="300" swimtime="00:04:00.11" />
                    <SPLIT distance="350" swimtime="00:04:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="14" clubid="4821" name="Uczniowski Klub Sportowy Delfin Legionowo">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Dziadecki" birthdate="1981-05-26" gender="M" nation="POL" license="101414700147" athleteid="4837">
              <RESULTS>
                <RESULT eventid="1110" points="279" swimtime="00:01:24.62" resultid="4838" heatid="5794" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="298" reactiontime="+74" swimtime="00:00:37.77" resultid="4839" heatid="5870" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Strzeszewski" birthdate="1998-08-27" gender="M" nation="POL" license="101414700146" swrid="5461237" athleteid="4822">
              <RESULTS>
                <RESULT eventid="1076" points="533" reactiontime="+62" swimtime="00:00:26.82" resultid="4823" heatid="5782" lane="7" entrytime="00:00:27.30" />
                <RESULT eventid="1212" points="449" reactiontime="+65" swimtime="00:02:09.73" resultid="4824" heatid="5835" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="100" swimtime="00:01:00.90" />
                    <SPLIT distance="150" swimtime="00:01:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="548" reactiontime="+68" swimtime="00:00:54.90" resultid="4825" heatid="5856" lane="5" entrytime="00:00:58.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="541" reactiontime="+62" swimtime="00:00:24.73" resultid="4826" heatid="5937" lane="4" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Perl" birthdate="1996-06-07" gender="M" nation="POL" license="101414700068" swrid="4282344" athleteid="4840">
              <RESULTS>
                <RESULT eventid="1110" points="547" reactiontime="+68" swimtime="00:01:07.64" resultid="4841" heatid="5796" lane="5" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="637" reactiontime="+64" swimtime="00:00:29.34" resultid="4842" heatid="5874" lane="4" entrytime="00:00:28.26" entrycourse="SCM" />
                <RESULT eventid="1333" points="452" reactiontime="+70" swimtime="00:01:04.19" resultid="4843" heatid="5892" lane="4" entrytime="00:01:02.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4844" heatid="5940" lane="4" entrytime="00:00:22.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" license="101414700141" swrid="4992689" athleteid="4845">
              <RESULTS>
                <RESULT eventid="1144" points="219" reactiontime="+81" swimtime="00:00:36.86" resultid="4846" heatid="5806" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1212" points="245" swimtime="00:02:38.65" resultid="4847" heatid="5832" lane="9" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:56.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="210" reactiontime="+88" swimtime="00:02:57.47" resultid="4848" heatid="5906" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="150" swimtime="00:02:10.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="280" swimtime="00:00:30.78" resultid="4849" heatid="5931" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1537" points="208" reactiontime="+89" swimtime="00:01:21.51" resultid="4850" heatid="5959" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Żbikowska" birthdate="1996-01-31" gender="F" nation="POL" license="101414600091" swrid="4605445" athleteid="4832">
              <RESULTS>
                <RESULT eventid="1093" points="427" reactiontime="+71" swimtime="00:01:22.81" resultid="4833" heatid="5788" lane="2" entrytime="00:01:25.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="491" reactiontime="+69" swimtime="00:00:36.19" resultid="4834" heatid="5864" lane="2" entrytime="00:00:37.99" />
                <RESULT eventid="1316" points="418" swimtime="00:01:15.55" resultid="4835" heatid="5880" lane="7" entrytime="00:01:15.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="441" reactiontime="+68" swimtime="00:00:30.12" resultid="4836" heatid="5920" lane="8" entrytime="00:00:31.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Chudorlińska" birthdate="2001-03-13" gender="F" nation="POL" license="101414600039" swrid="4425462" athleteid="4827">
              <RESULTS>
                <RESULT eventid="1282" points="454" reactiontime="+67" swimtime="00:00:37.15" resultid="4829" heatid="5864" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1316" points="412" reactiontime="+65" swimtime="00:01:15.89" resultid="4830" heatid="5880" lane="5" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="439" reactiontime="+66" swimtime="00:00:30.16" resultid="4831" heatid="5921" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1059" points="350" reactiontime="+67" swimtime="00:00:34.57" resultid="5726" heatid="5770" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="5278" name="NoStars">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Medvediev" birthdate="1962-08-09" gender="M" nation="UKR" athleteid="5279">
              <RESULTS>
                <RESULT eventid="1110" points="422" reactiontime="+77" swimtime="00:01:13.73" resultid="5280" heatid="5795" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="350" swimtime="00:02:35.51" resultid="5281" heatid="5819" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="458" reactiontime="+77" swimtime="00:00:32.75" resultid="5282" heatid="5873" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1333" points="357" reactiontime="+72" swimtime="00:01:09.44" resultid="5283" heatid="5891" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="391" reactiontime="+78" swimtime="00:02:44.31" resultid="5284" heatid="5950" lane="0" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.72" />
                    <SPLIT distance="150" swimtime="00:02:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="309" reactiontime="+80" swimtime="00:01:10.60" resultid="5285" heatid="5969" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="4800" name="Towarzystwo Pływackie ,,Masters&apos;&apos; Opole">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" license="100607700003" swrid="4843497" athleteid="4806">
              <RESULTS>
                <RESULT eventid="1076" points="379" reactiontime="+77" swimtime="00:00:30.03" resultid="4807" heatid="5773" lane="8" />
                <RESULT eventid="1144" points="364" reactiontime="+63" swimtime="00:00:31.12" resultid="4808" heatid="5810" lane="8" entrytime="00:00:31.44" entrycourse="SCM" />
                <RESULT eventid="1265" points="378" reactiontime="+88" swimtime="00:01:02.12" resultid="4809" heatid="5845" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4810" heatid="5907" lane="4" entrytime="00:02:28.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Vogel" birthdate="1981-09-20" gender="M" nation="POL" license="100607700016" athleteid="4811">
              <RESULTS>
                <RESULT eventid="1076" points="398" reactiontime="+75" swimtime="00:00:29.56" resultid="4812" heatid="5772" lane="4" />
                <RESULT eventid="1333" points="307" reactiontime="+75" swimtime="00:01:12.99" resultid="4813" heatid="5883" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="283" reactiontime="+75" swimtime="00:01:13.54" resultid="4814" heatid="5957" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Bartnikowska" birthdate="1990-08-21" gender="F" nation="POL" license="100607600002" swrid="5295108" athleteid="4801">
              <RESULTS>
                <RESULT eventid="1059" points="422" reactiontime="+68" swimtime="00:00:32.49" resultid="4802" heatid="5770" lane="6" entrytime="00:00:34.45" entrycourse="SCM" />
                <RESULT eventid="1127" points="479" reactiontime="+68" swimtime="00:00:32.70" resultid="4803" heatid="5802" lane="0" entrytime="00:00:33.09" entrycourse="SCM" />
                <RESULT eventid="1247" points="437" reactiontime="+79" swimtime="00:01:06.21" resultid="4804" heatid="5839" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" status="DNS" swimtime="00:00:00.00" resultid="4805" heatid="5901" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="4580" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-16" gender="M" nation="POL" license="500309700377" swrid="4186249" athleteid="4581">
              <RESULTS>
                <RESULT eventid="1076" points="349" reactiontime="+75" swimtime="00:00:30.88" resultid="4582" heatid="5779" lane="1" entrytime="00:00:30.55" />
                <RESULT eventid="1178" points="332" reactiontime="+81" swimtime="00:02:38.26" resultid="4583" heatid="5818" lane="4" entrytime="00:02:38.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="370" reactiontime="+77" swimtime="00:01:02.59" resultid="4584" heatid="5854" lane="5" entrytime="00:01:02.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="329" swimtime="00:01:11.38" resultid="4585" heatid="5890" lane="9" entrytime="00:01:11.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="364" reactiontime="+77" swimtime="00:00:28.22" resultid="4586" heatid="5934" lane="3" entrytime="00:00:27.95" entrycourse="SCM" />
                <RESULT eventid="1571" points="326" reactiontime="+80" swimtime="00:01:09.36" resultid="4587" heatid="5969" lane="1" entrytime="00:01:09.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Wasilewicz" birthdate="1959-06-15" gender="F" nation="POL" license="500309600230" swrid="4876623" athleteid="4592">
              <RESULTS>
                <RESULT eventid="1195" points="158" swimtime="00:03:24.07" resultid="4593" heatid="5823" lane="0" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="199" swimtime="00:01:25.99" resultid="4594" heatid="5841" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="225" swimtime="00:00:37.66" resultid="4595" heatid="5918" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1520" points="98" reactiontime="+88" swimtime="00:01:58.67" resultid="4596" heatid="5953" lane="0" entrytime="00:01:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Matusik" birthdate="1956-11-05" gender="M" nation="POL" license="500309700229" swrid="4876624" athleteid="4588">
              <RESULTS>
                <RESULT eventid="1110" points="188" reactiontime="+85" swimtime="00:01:36.51" resultid="4589" heatid="5792" lane="7" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="237" swimtime="00:00:40.80" resultid="4590" heatid="5870" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1469" points="188" reactiontime="+76" swimtime="00:00:35.13" resultid="4591" heatid="5929" lane="2" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3202" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sikora" birthdate="1998-01-01" gender="M" nation="POL" swrid="4713953" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1178" points="294" reactiontime="+72" swimtime="00:02:44.87" resultid="3203" heatid="5819" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:02:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="370" reactiontime="+69" swimtime="00:01:02.56" resultid="3204" heatid="5853" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="283" reactiontime="+73" swimtime="00:01:15.00" resultid="3206" heatid="5888" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="381" reactiontime="+68" swimtime="00:00:27.79" resultid="3207" heatid="5936" lane="0" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5358" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Kowalczyk" birthdate="1973-01-01" gender="M" nation="POL" athleteid="5357">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5359" heatid="5778" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="5360" heatid="5849" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5361" heatid="5887" lane="1" entrytime="00:01:22.00" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="5362" heatid="5927" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5363" heatid="5967" lane="0" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2736" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Korzuchowski " birthdate="1999-01-01" gender="M" nation="POL" swrid="4598470" athleteid="2735">
              <RESULTS>
                <RESULT eventid="1144" points="350" reactiontime="+57" swimtime="00:00:31.51" resultid="2737" heatid="5809" lane="7" entrytime="00:00:32.10" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1212" status="DSQ" swimtime="00:00:00.00" resultid="2738" heatid="5833" lane="2" entrytime="00:02:21.30" />
                <RESULT eventid="1265" points="439" reactiontime="+71" swimtime="00:00:59.09" resultid="2739" heatid="5854" lane="1" entrytime="00:01:03.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="310" reactiontime="+56" swimtime="00:02:36.02" resultid="2740" heatid="5908" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:14.95" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="369" reactiontime="+58" swimtime="00:01:07.34" resultid="2741" heatid="5961" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="239" reactiontime="+77" swimtime="00:05:41.86" resultid="2742" heatid="5982" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:01:58.66" />
                    <SPLIT distance="200" swimtime="00:02:42.20" />
                    <SPLIT distance="250" swimtime="00:03:27.14" />
                    <SPLIT distance="300" swimtime="00:04:12.32" />
                    <SPLIT distance="350" swimtime="00:04:57.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3097" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Rybak" birthdate="1996-01-01" gender="M" nation="POL" swrid="4297546" athleteid="3096">
              <RESULTS>
                <RESULT eventid="1076" points="467" reactiontime="+69" swimtime="00:00:28.02" resultid="3098" heatid="5778" lane="4" entrytime="00:00:31.25" />
                <RESULT eventid="1178" points="415" swimtime="00:02:26.93" resultid="3099" heatid="5818" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:10.26" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="505" reactiontime="+75" swimtime="00:00:31.69" resultid="3100" heatid="5873" lane="0" entrytime="00:00:33.50" />
                <RESULT eventid="1333" points="412" reactiontime="+79" swimtime="00:01:06.18" resultid="3101" heatid="5887" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="512" swimtime="00:00:25.20" resultid="3102" heatid="5935" lane="9" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WISKRA" nation="POL" clubid="3494" name="Masters Wisła Kraków">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Korba" birthdate="1969-06-25" gender="M" nation="POL" swrid="5066074" athleteid="3502">
              <RESULTS>
                <RESULT eventid="1110" points="364" reactiontime="+82" swimtime="00:01:17.46" resultid="3503" heatid="5794" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="382" reactiontime="+83" swimtime="00:02:16.93" resultid="3504" heatid="5833" lane="7" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                    <SPLIT distance="150" swimtime="00:01:42.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="396" swimtime="00:01:01.16" resultid="3505" heatid="5854" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="390" reactiontime="+79" swimtime="00:00:34.54" resultid="3506" heatid="5872" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1503" points="320" swimtime="00:02:55.62" resultid="3507" heatid="5949" lane="9" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:24.06" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="369" reactiontime="+90" swimtime="00:04:55.91" resultid="3508" heatid="5982" lane="8" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:46.83" />
                    <SPLIT distance="200" swimtime="00:02:24.80" />
                    <SPLIT distance="250" swimtime="00:03:03.01" />
                    <SPLIT distance="300" swimtime="00:03:41.40" />
                    <SPLIT distance="350" swimtime="00:04:20.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Krokoszyński" birthdate="1930-05-04" gender="M" nation="POL" swrid="4302634" athleteid="3495">
              <RESULTS>
                <RESULT eventid="1110" points="41" reactiontime="+120" swimtime="00:02:39.56" resultid="3496" heatid="5789" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="37" reactiontime="+89" swimtime="00:01:06.38" resultid="3497" heatid="5804" lane="9" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1265" points="44" reactiontime="+119" swimtime="00:02:06.53" resultid="3498" heatid="5845" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="44" swimtime="00:01:11.41" resultid="3499" heatid="5866" lane="2" />
                <RESULT eventid="1469" points="46" swimtime="00:00:55.94" resultid="3500" heatid="5924" lane="7" />
                <RESULT eventid="1537" points="28" reactiontime="+95" swimtime="00:02:38.44" resultid="3501" heatid="5956" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4214" nation="POL" clubid="3343" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Paluszak" birthdate="1967-02-17" gender="M" nation="POL" swrid="5471792" athleteid="3380">
              <RESULTS>
                <RESULT eventid="1076" points="155" reactiontime="+76" swimtime="00:00:40.49" resultid="3381" heatid="5772" lane="6" />
                <RESULT eventid="1212" points="122" reactiontime="+78" swimtime="00:03:20.33" resultid="3382" heatid="5829" lane="0" entrytime="00:03:31.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                    <SPLIT distance="150" swimtime="00:02:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="117" reactiontime="+74" swimtime="00:01:40.49" resultid="3383" heatid="5884" lane="0" entrytime="00:01:45.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="107" reactiontime="+71" swimtime="00:01:40.51" resultid="3384" heatid="5965" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Burdelak" birthdate="1991-07-06" gender="F" nation="POL" swrid="4072596" athleteid="3365">
              <RESULTS>
                <RESULT eventid="1093" points="528" reactiontime="+68" swimtime="00:01:17.14" resultid="3366" heatid="5788" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="546" reactiontime="+66" swimtime="00:00:34.93" resultid="3367" heatid="5864" lane="4" entrytime="00:00:34.80" />
                <RESULT eventid="1316" points="495" swimtime="00:01:11.41" resultid="3368" heatid="5881" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="534" reactiontime="+66" swimtime="00:00:28.25" resultid="3369" heatid="5921" lane="4" entrytime="00:00:28.10" />
                <RESULT eventid="1554" points="399" reactiontime="+69" swimtime="00:01:14.13" resultid="3370" heatid="5964" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szymański" birthdate="1980-10-04" gender="M" nation="POL" swrid="4542528" athleteid="3728">
              <RESULTS>
                <RESULT eventid="1076" points="499" reactiontime="+77" swimtime="00:00:27.41" resultid="3729" heatid="5772" lane="3" />
                <RESULT eventid="1144" points="498" reactiontime="+79" swimtime="00:00:28.02" resultid="3730" heatid="5811" lane="6" entrytime="00:00:28.15" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1333" points="517" reactiontime="+71" swimtime="00:01:01.38" resultid="3731" heatid="5893" lane="8" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="528" reactiontime="+75" swimtime="00:00:24.93" resultid="3732" heatid="5939" lane="5" entrytime="00:00:24.50" />
                <RESULT eventid="1537" points="498" reactiontime="+74" swimtime="00:01:00.97" resultid="3733" heatid="5962" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Szymańska" birthdate="1985-05-31" gender="F" nation="POL" swrid="5312493" athleteid="3723">
              <RESULTS>
                <RESULT eventid="1059" points="156" reactiontime="+96" swimtime="00:00:45.26" resultid="3724" heatid="5767" lane="8" />
                <RESULT eventid="1316" points="198" reactiontime="+87" swimtime="00:01:36.84" resultid="3725" heatid="5877" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3726" heatid="5918" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1588" points="210" reactiontime="+95" swimtime="00:06:33.41" resultid="3727" heatid="5973" lane="5" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:02:18.70" />
                    <SPLIT distance="200" swimtime="00:03:10.07" />
                    <SPLIT distance="250" swimtime="00:04:00.56" />
                    <SPLIT distance="300" swimtime="00:04:52.27" />
                    <SPLIT distance="350" swimtime="00:05:43.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Nawrocka" birthdate="1990-02-15" gender="F" nation="POL" swrid="4806455" athleteid="3350">
              <RESULTS>
                <RESULT eventid="1161" points="384" reactiontime="+86" swimtime="00:02:47.57" resultid="3351" heatid="5814" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                    <SPLIT distance="150" swimtime="00:02:07.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="372" reactiontime="+85" swimtime="00:00:39.71" resultid="3352" heatid="5863" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1316" points="407" reactiontime="+80" swimtime="00:01:16.22" resultid="3353" heatid="5880" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="417" reactiontime="+77" swimtime="00:00:30.68" resultid="3354" heatid="5920" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1588" points="313" reactiontime="+81" swimtime="00:05:44.40" resultid="3355" heatid="5975" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                    <SPLIT distance="200" swimtime="00:02:46.63" />
                    <SPLIT distance="250" swimtime="00:03:31.20" />
                    <SPLIT distance="300" swimtime="00:04:15.74" />
                    <SPLIT distance="350" swimtime="00:05:00.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Nowak" birthdate="1952-12-17" gender="M" nation="POL" swrid="4302652" athleteid="3403">
              <RESULTS>
                <RESULT eventid="1110" points="263" reactiontime="+91" swimtime="00:01:26.29" resultid="3404" heatid="5793" lane="0" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="175" swimtime="00:03:15.69" resultid="3405" heatid="5817" lane="9" entrytime="00:03:26.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:38.54" />
                    <SPLIT distance="150" swimtime="00:02:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="265" swimtime="00:00:39.31" resultid="3406" heatid="5871" lane="9" entrytime="00:00:37.90" />
                <RESULT eventid="1333" points="202" reactiontime="+86" swimtime="00:01:23.96" resultid="3407" heatid="5887" lane="0" entrytime="00:01:23.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="209" reactiontime="+94" swimtime="00:03:22.40" resultid="3408" heatid="5947" lane="8" entrytime="00:03:28.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:38.13" />
                    <SPLIT distance="150" swimtime="00:02:31.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Makomaski" birthdate="1986-05-09" gender="M" nation="POL" swrid="4992665" athleteid="3356">
              <RESULTS>
                <RESULT eventid="1110" points="335" reactiontime="+79" swimtime="00:01:19.64" resultid="3357" heatid="5794" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="383" swimtime="00:00:34.75" resultid="3358" heatid="5872" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1469" points="346" reactiontime="+80" swimtime="00:00:28.70" resultid="3359" heatid="5934" lane="1" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Pfitzner" birthdate="1986-05-24" gender="M" nation="POL" swrid="4992671" athleteid="3397">
              <RESULTS>
                <RESULT eventid="1144" points="381" reactiontime="+84" swimtime="00:00:30.63" resultid="3398" heatid="5810" lane="2" entrytime="00:00:30.80" />
                <RESULT eventid="1212" points="420" swimtime="00:02:12.59" resultid="3399" heatid="5835" lane="9" entrytime="00:02:07.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="150" swimtime="00:01:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="444" reactiontime="+74" swimtime="00:00:58.90" resultid="3400" heatid="5856" lane="3" entrytime="00:00:58.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="3401" heatid="5936" lane="5" entrytime="00:00:26.80" />
                <RESULT eventid="1537" points="356" reactiontime="+79" swimtime="00:01:08.18" resultid="3402" heatid="5961" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" swrid="4302692" athleteid="3371">
              <RESULTS>
                <RESULT eventid="1195" points="68" swimtime="00:04:29.91" resultid="3372" heatid="5822" lane="7" entrytime="00:04:39.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.78" />
                    <SPLIT distance="100" swimtime="00:02:11.86" />
                    <SPLIT distance="150" swimtime="00:03:22.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="58" swimtime="00:02:09.25" resultid="3373" heatid="5840" lane="4" entrytime="00:02:13.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="73" swimtime="00:09:17.46" resultid="3374" heatid="5972" lane="5" entrytime="00:09:38.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.78" />
                    <SPLIT distance="100" swimtime="00:02:14.67" />
                    <SPLIT distance="150" swimtime="00:03:26.80" />
                    <SPLIT distance="200" swimtime="00:04:37.94" />
                    <SPLIT distance="250" swimtime="00:05:48.30" />
                    <SPLIT distance="300" swimtime="00:06:58.40" />
                    <SPLIT distance="350" swimtime="00:08:09.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Sutowski" birthdate="1959-12-03" gender="M" nation="POL" swrid="4992657" athleteid="3360">
              <RESULTS>
                <RESULT eventid="1212" points="150" reactiontime="+100" swimtime="00:03:06.81" resultid="3361" heatid="5829" lane="5" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.48" />
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                    <SPLIT distance="150" swimtime="00:02:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="145" reactiontime="+118" swimtime="00:01:25.41" resultid="3362" heatid="5848" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="132" swimtime="00:00:39.51" resultid="3363" heatid="5927" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="1605" points="154" reactiontime="+109" swimtime="00:06:35.18" resultid="3364" heatid="5978" lane="5" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                    <SPLIT distance="150" swimtime="00:02:22.94" />
                    <SPLIT distance="200" swimtime="00:03:14.64" />
                    <SPLIT distance="250" swimtime="00:04:05.53" />
                    <SPLIT distance="300" swimtime="00:04:56.87" />
                    <SPLIT distance="350" swimtime="00:05:47.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kośla" birthdate="1993-01-05" gender="F" nation="POL" swrid="4086961" athleteid="3344">
              <RESULTS>
                <RESULT eventid="1059" points="430" reactiontime="+75" swimtime="00:00:32.28" resultid="3345" heatid="5771" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1127" points="496" reactiontime="+80" swimtime="00:00:32.32" resultid="3346" heatid="5802" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1384" points="474" reactiontime="+71" swimtime="00:02:32.46" resultid="3347" heatid="5903" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.46" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3348" heatid="5921" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1520" points="531" reactiontime="+67" swimtime="00:01:07.76" resultid="3349" heatid="5955" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" athleteid="3390">
              <RESULTS>
                <RESULT eventid="1076" points="388" reactiontime="+78" swimtime="00:00:29.81" resultid="3391" heatid="5777" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1110" points="409" swimtime="00:01:14.55" resultid="3392" heatid="5795" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="380" reactiontime="+77" swimtime="00:01:02.00" resultid="3393" heatid="5854" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="486" reactiontime="+78" swimtime="00:00:32.11" resultid="3394" heatid="5873" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1469" points="467" reactiontime="+75" swimtime="00:00:25.98" resultid="3395" heatid="5935" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1571" points="260" reactiontime="+79" swimtime="00:01:14.78" resultid="3396" heatid="5968" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" swrid="4183802" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1144" points="355" reactiontime="+72" swimtime="00:00:31.37" resultid="3376" heatid="5809" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1178" points="392" reactiontime="+86" swimtime="00:02:29.69" resultid="3377" heatid="5818" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:55.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="408" reactiontime="+81" swimtime="00:01:00.56" resultid="3378" heatid="5854" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="375" reactiontime="+77" swimtime="00:01:08.32" resultid="3379" heatid="5889" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Sutowski" birthdate="1993-02-18" gender="M" nation="POL" swrid="4073514" athleteid="3385">
              <RESULTS>
                <RESULT eventid="1076" points="291" swimtime="00:00:32.82" resultid="3386" heatid="5777" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1265" points="294" swimtime="00:01:07.52" resultid="3387" heatid="5853" lane="9" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="229" reactiontime="+74" swimtime="00:01:20.50" resultid="3388" heatid="5886" lane="1" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="3389" heatid="5933" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="485" swimtime="00:01:44.09" resultid="3736" heatid="5914" lane="7" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="100" swimtime="00:00:50.58" />
                    <SPLIT distance="150" swimtime="00:01:18.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3728" number="1" />
                    <RELAYPOSITION athleteid="3397" number="2" />
                    <RELAYPOSITION athleteid="3356" number="3" />
                    <RELAYPOSITION athleteid="3390" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="477" reactiontime="+69" swimtime="00:01:55.73" resultid="3738" heatid="5989" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                    <SPLIT distance="150" swimtime="00:01:30.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3728" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3356" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3397" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="3390" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="194" swimtime="00:02:21.09" resultid="3737" heatid="5912" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3403" number="1" />
                    <RELAYPOSITION athleteid="3360" number="2" />
                    <RELAYPOSITION athleteid="3380" number="3" />
                    <RELAYPOSITION athleteid="3385" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1622" points="393" reactiontime="+70" swimtime="00:02:19.71" resultid="3739" heatid="5986" lane="4" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:43.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3344" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3350" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3365" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3723" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1418" points="393" reactiontime="+73" swimtime="00:02:06.24" resultid="3740" heatid="5910" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="100" swimtime="00:00:59.98" />
                    <SPLIT distance="150" swimtime="00:01:37.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3365" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3350" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3723" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="3344" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="517" reactiontime="+75" swimtime="00:01:59.87" resultid="3734" heatid="5838" lane="4" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="150" swimtime="00:01:32.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3728" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3390" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3344" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3365" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="291" reactiontime="+84" swimtime="00:02:25.16" resultid="3735" heatid="5838" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.35" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3723" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="3350" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3397" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3385" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TOOLE" nation="POL" clubid="2864" name="Ukp Torpeda Oleśnica">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-06-29" gender="M" nation="POL" swrid="5416779" athleteid="2865">
              <RESULTS>
                <RESULT eventid="1178" points="98" reactiontime="+117" swimtime="00:03:57.78" resultid="2866" heatid="5816" lane="2" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                    <SPLIT distance="100" swimtime="00:02:01.25" />
                    <SPLIT distance="150" swimtime="00:03:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="112" reactiontime="+104" swimtime="00:03:25.54" resultid="2867" heatid="5829" lane="9" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:42.24" />
                    <SPLIT distance="150" swimtime="00:02:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="107" swimtime="00:01:34.60" resultid="2868" heatid="5848" lane="7" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" status="DNS" swimtime="00:00:00.00" resultid="2869" heatid="5898" lane="9" entrytime="00:03:59.00" />
                <RESULT eventid="1469" points="128" reactiontime="+83" swimtime="00:00:39.98" resultid="2870" heatid="5927" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1605" points="114" reactiontime="+96" swimtime="00:07:16.60" resultid="2871" heatid="5978" lane="1" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                    <SPLIT distance="100" swimtime="00:01:42.97" />
                    <SPLIT distance="150" swimtime="00:02:38.78" />
                    <SPLIT distance="200" swimtime="00:03:34.68" />
                    <SPLIT distance="250" swimtime="00:04:31.41" />
                    <SPLIT distance="300" swimtime="00:05:27.65" />
                    <SPLIT distance="350" swimtime="00:06:23.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3638" name="niezrzeszony" />
        <CLUB type="CLUB" nation="POL" clubid="3225" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Wielechowska" birthdate="1990-01-01" gender="F" nation="POL" athleteid="3224">
              <RESULTS>
                <RESULT eventid="1127" points="270" reactiontime="+73" swimtime="00:00:39.58" resultid="3226" heatid="5801" lane="9" entrytime="00:00:37.70" />
                <RESULT eventid="1195" points="257" reactiontime="+87" swimtime="00:02:53.62" resultid="3227" heatid="5824" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="150" swimtime="00:02:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="284" swimtime="00:00:34.87" resultid="3228" heatid="5919" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1520" points="273" reactiontime="+80" swimtime="00:01:24.58" resultid="3229" heatid="5954" lane="7" entrytime="00:01:20.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00701" nation="POL" region="01" clubid="4567" name="MKS Dziewiątka Dzierżoniów">
          <ATHLETES>
            <ATHLETE firstname="Edyta" lastname="Bejster" birthdate="1981-05-21" gender="F" nation="POL" license="100701600124" swrid="5464069" athleteid="4574">
              <RESULTS>
                <RESULT eventid="1059" points="140" swimtime="00:00:46.88" resultid="4575" heatid="5768" lane="2" entrytime="00:00:45.64" />
                <RESULT eventid="1195" points="138" reactiontime="+85" swimtime="00:03:33.22" resultid="4576" heatid="5823" lane="1" entrytime="00:03:13.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="166" swimtime="00:00:51.87" resultid="4577" heatid="5862" lane="7" entrytime="00:00:48.23" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1316" status="DSQ" swimtime="00:00:00.00" resultid="4578" heatid="5877" lane="7" entrytime="00:01:55.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="163" reactiontime="+86" swimtime="00:00:41.94" resultid="4579" heatid="5918" lane="8" entrytime="00:00:38.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Pisarska" birthdate="1981-11-06" gender="F" nation="POL" license="100701600113" swrid="5464072" athleteid="4568">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1059" points="565" reactiontime="+66" swimtime="00:00:29.49" resultid="4569" heatid="5768" lane="6" entrytime="00:00:45.64" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1127" points="520" reactiontime="+62" swimtime="00:00:31.83" resultid="4570" heatid="5802" lane="5" entrytime="00:00:31.28" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1316" points="542" reactiontime="+66" swimtime="00:01:09.30" resultid="4571" heatid="5881" lane="4" entrytime="00:01:07.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy od Rekordu Polski" eventid="1451" points="572" reactiontime="+65" swimtime="00:00:27.61" resultid="4572" heatid="5922" lane="3" entrytime="00:00:26.93" />
                <RESULT eventid="1520" points="489" reactiontime="+62" swimtime="00:01:09.65" resultid="4573" heatid="5955" lane="6" entrytime="00:01:09.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3217" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Kruczkowski" birthdate="1997-01-01" gender="M" nation="POL" swrid="4225992" athleteid="3216">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3218" heatid="5776" lane="8" entrytime="00:00:35.51" />
                <RESULT eventid="1144" points="286" reactiontime="+67" swimtime="00:00:33.69" resultid="3219" heatid="5809" lane="4" entrytime="00:00:31.81" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3220" heatid="5888" lane="0" entrytime="00:01:19.00" />
                <RESULT eventid="1401" points="298" reactiontime="+72" swimtime="00:02:38.09" resultid="3221" heatid="5907" lane="5" entrytime="00:02:28.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:56.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="310" reactiontime="+71" swimtime="00:01:11.34" resultid="3222" heatid="5960" lane="5" entrytime="00:01:12.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="3223" heatid="5981" lane="5" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3837" name="SMT Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Kowalczyk" birthdate="1976-01-31" gender="F" nation="POL" athleteid="3847">
              <RESULTS>
                <RESULT eventid="1059" points="330" reactiontime="+89" swimtime="00:00:35.28" resultid="3848" heatid="5769" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1195" points="325" reactiontime="+94" swimtime="00:02:40.54" resultid="3849" heatid="5824" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:58.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="328" reactiontime="+97" swimtime="00:01:21.94" resultid="3850" heatid="5879" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="342" reactiontime="+95" swimtime="00:00:32.77" resultid="3851" heatid="5919" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1588" points="301" swimtime="00:05:49.02" resultid="3852" heatid="5975" lane="9" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:05.54" />
                    <SPLIT distance="200" swimtime="00:02:51.02" />
                    <SPLIT distance="250" swimtime="00:03:36.10" />
                    <SPLIT distance="300" swimtime="00:04:21.46" />
                    <SPLIT distance="350" swimtime="00:05:06.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Łubiński" birthdate="1975-07-23" gender="M" nation="POL" athleteid="3863">
              <RESULTS>
                <RESULT eventid="1265" points="136" reactiontime="+98" swimtime="00:01:27.34" resultid="3864" heatid="5848" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="183" reactiontime="+76" swimtime="00:00:44.46" resultid="3865" heatid="5869" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1469" points="164" reactiontime="+87" swimtime="00:00:36.82" resultid="3866" heatid="5927" lane="5" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Bałka" birthdate="1987-11-22" gender="M" nation="POL" swrid="4072794" athleteid="3843">
              <RESULTS>
                <RESULT eventid="1178" points="328" reactiontime="+73" swimtime="00:02:38.89" resultid="3844" heatid="5817" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="350" reactiontime="+74" swimtime="00:02:33.54" resultid="3845" heatid="5898" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="390" reactiontime="+70" swimtime="00:01:05.37" resultid="3846" heatid="5970" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Ryczak" birthdate="1996-04-22" gender="F" nation="POL" swrid="4225999" athleteid="3877">
              <RESULTS>
                <RESULT eventid="1059" points="503" reactiontime="+69" swimtime="00:00:30.65" resultid="3878" heatid="5770" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1127" points="578" reactiontime="+65" swimtime="00:00:30.73" resultid="3879" heatid="5802" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1247" points="508" swimtime="00:01:02.96" resultid="3880" heatid="5844" lane="9" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="546" swimtime="00:00:28.05" resultid="3881" heatid="5922" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1520" points="530" reactiontime="+63" swimtime="00:01:07.80" resultid="3882" heatid="5955" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Rożek" birthdate="1984-05-09" gender="M" nation="POL" athleteid="3870">
              <RESULTS>
                <RESULT eventid="1178" points="168" reactiontime="+92" swimtime="00:03:18.33" resultid="3871" heatid="5816" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:01:36.05" />
                    <SPLIT distance="150" swimtime="00:02:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="208" reactiontime="+82" swimtime="00:02:47.62" resultid="3872" heatid="5830" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="241" reactiontime="+81" swimtime="00:01:12.20" resultid="3873" heatid="5850" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="179" reactiontime="+84" swimtime="00:01:27.33" resultid="3874" heatid="5885" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="270" reactiontime="+80" swimtime="00:00:31.17" resultid="3875" heatid="5929" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1605" points="194" reactiontime="+90" swimtime="00:06:06.17" resultid="3876" heatid="5979" lane="2" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                    <SPLIT distance="150" swimtime="00:02:13.61" />
                    <SPLIT distance="200" swimtime="00:03:00.72" />
                    <SPLIT distance="250" swimtime="00:03:47.69" />
                    <SPLIT distance="300" swimtime="00:04:34.71" />
                    <SPLIT distance="350" swimtime="00:05:21.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Zając" birthdate="1966-06-30" gender="M" nation="POL" athleteid="3893">
              <RESULTS>
                <RESULT eventid="1076" points="255" reactiontime="+96" swimtime="00:00:34.26" resultid="3894" heatid="5776" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1333" points="205" reactiontime="+89" swimtime="00:01:23.47" resultid="3895" heatid="5886" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="271" reactiontime="+89" swimtime="00:00:31.15" resultid="3896" heatid="5931" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Zielińska" birthdate="1980-12-12" gender="F" nation="POL" swrid="5185937" athleteid="3897">
              <RESULTS>
                <RESULT eventid="1127" points="358" reactiontime="+70" swimtime="00:00:36.03" resultid="3898" heatid="5800" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1161" points="377" swimtime="00:02:48.58" resultid="3899" heatid="5814" lane="7" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:17.87" />
                    <SPLIT distance="150" swimtime="00:02:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="376" reactiontime="+72" swimtime="00:01:18.28" resultid="3900" heatid="5879" lane="6" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="355" reactiontime="+94" swimtime="00:02:47.95" resultid="3901" heatid="5903" lane="0" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="363" reactiontime="+72" swimtime="00:01:16.88" resultid="3902" heatid="5954" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="353" swimtime="00:05:30.98" resultid="3903" heatid="5975" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:01:59.84" />
                    <SPLIT distance="200" swimtime="00:02:42.64" />
                    <SPLIT distance="250" swimtime="00:03:25.44" />
                    <SPLIT distance="300" swimtime="00:04:08.93" />
                    <SPLIT distance="350" swimtime="00:04:51.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Krzyżostaniak" birthdate="1993-01-20" gender="F" nation="POL" swrid="4087097" athleteid="3853">
              <RESULTS>
                <RESULT eventid="1127" points="504" reactiontime="+80" swimtime="00:00:32.16" resultid="3854" heatid="5802" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1316" points="435" reactiontime="+82" swimtime="00:01:14.58" resultid="3855" heatid="5879" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="3856" heatid="5921" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1520" points="437" reactiontime="+81" swimtime="00:01:12.33" resultid="3857" heatid="5955" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Sawrymowicz" birthdate="1957-01-01" gender="M" nation="POL" athleteid="3883">
              <RESULTS>
                <RESULT eventid="1333" points="76" swimtime="00:01:55.93" resultid="3884" heatid="5883" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="111" swimtime="00:07:21.04" resultid="3885" heatid="5978" lane="8" entrytime="00:07:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                    <SPLIT distance="100" swimtime="00:01:45.99" />
                    <SPLIT distance="150" swimtime="00:02:41.77" />
                    <SPLIT distance="200" swimtime="00:03:37.39" />
                    <SPLIT distance="250" swimtime="00:04:34.41" />
                    <SPLIT distance="300" swimtime="00:05:32.15" />
                    <SPLIT distance="350" swimtime="00:06:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Adamiak" birthdate="1987-08-03" gender="F" nation="POL" athleteid="3838">
              <RESULTS>
                <RESULT eventid="1093" points="202" reactiontime="+91" swimtime="00:01:46.20" resultid="3839" heatid="5786" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="156" reactiontime="+87" swimtime="00:03:24.87" resultid="3840" heatid="5822" lane="5" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="150" swimtime="00:02:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="197" reactiontime="+89" swimtime="00:00:49.08" resultid="3841" heatid="5862" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="1588" points="186" swimtime="00:06:49.51" resultid="3842" heatid="5973" lane="7" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                    <SPLIT distance="100" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:02:29.75" />
                    <SPLIT distance="200" swimtime="00:03:22.65" />
                    <SPLIT distance="250" swimtime="00:04:15.10" />
                    <SPLIT distance="300" swimtime="00:05:07.43" />
                    <SPLIT distance="350" swimtime="00:05:59.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Kudra" birthdate="1959-11-24" gender="F" nation="POL" athleteid="3858">
              <RESULTS>
                <RESULT eventid="1195" points="62" reactiontime="+138" swimtime="00:04:37.53" resultid="3859" heatid="5822" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                    <SPLIT distance="100" swimtime="00:02:09.46" />
                    <SPLIT distance="150" swimtime="00:03:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="62" swimtime="00:02:06.90" resultid="3860" heatid="5841" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="150" swimtime="00:00:53.68" resultid="3861" heatid="5862" lane="9" entrytime="00:00:55.00" />
                <RESULT eventid="1451" points="93" reactiontime="+139" swimtime="00:00:50.51" resultid="3862" heatid="5917" lane="0" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Stępień-Gielo" birthdate="1961-05-03" gender="F" nation="POL" athleteid="3886">
              <RESULTS>
                <RESULT eventid="1093" points="231" reactiontime="+84" swimtime="00:01:41.62" resultid="3887" heatid="5786" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="149" reactiontime="+78" swimtime="00:00:48.21" resultid="3888" heatid="5799" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1282" points="250" swimtime="00:00:45.33" resultid="3889" heatid="5862" lane="2" entrytime="00:00:47.00" />
                <RESULT eventid="1384" points="132" reactiontime="+73" swimtime="00:03:53.48" resultid="3890" heatid="5902" lane="0" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.87" />
                    <SPLIT distance="100" swimtime="00:01:57.53" />
                    <SPLIT distance="150" swimtime="00:02:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="207" reactiontime="+99" swimtime="00:03:47.25" resultid="3891" heatid="5943" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.38" />
                    <SPLIT distance="100" swimtime="00:01:52.80" />
                    <SPLIT distance="150" swimtime="00:02:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="166" reactiontime="+100" swimtime="00:07:05.48" resultid="3892" heatid="5973" lane="8" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:41.27" />
                    <SPLIT distance="150" swimtime="00:02:36.32" />
                    <SPLIT distance="200" swimtime="00:03:30.96" />
                    <SPLIT distance="250" swimtime="00:04:25.49" />
                    <SPLIT distance="300" swimtime="00:05:19.91" />
                    <SPLIT distance="350" swimtime="00:06:14.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Pawlewicz-Łubińska" birthdate="1972-03-14" gender="F" nation="POL" athleteid="3867">
              <RESULTS>
                <RESULT eventid="1247" points="56" reactiontime="+119" swimtime="00:02:11.07" resultid="3868" heatid="5840" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="62" swimtime="00:00:57.64" resultid="3869" heatid="5917" lane="9" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Zieliński" birthdate="1992-09-02" gender="M" nation="POL" swrid="4072211" athleteid="3904">
              <RESULTS>
                <RESULT eventid="1076" points="570" reactiontime="+75" swimtime="00:00:26.23" resultid="3905" heatid="5780" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1144" points="442" reactiontime="+80" swimtime="00:00:29.15" resultid="3906" heatid="5810" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1265" points="601" reactiontime="+78" swimtime="00:00:53.24" resultid="3907" heatid="5858" lane="9" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="597" reactiontime="+74" swimtime="00:00:23.93" resultid="3908" heatid="5937" lane="5" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="241" reactiontime="+78" swimtime="00:02:11.27" resultid="3916" heatid="5912" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="150" swimtime="00:01:44.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3870" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="3893" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3883" number="3" />
                    <RELAYPOSITION athleteid="3843" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="224" reactiontime="+80" swimtime="00:02:28.74" resultid="3917" heatid="5987" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="150" swimtime="00:01:57.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3843" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="3883" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3893" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3870" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="107" reactiontime="+95" swimtime="00:03:14.81" resultid="3912" heatid="5909" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:32.82" />
                    <SPLIT distance="150" swimtime="00:02:16.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3886" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="3858" number="2" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3838" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="3867" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="115" swimtime="00:03:30.52" resultid="3913" heatid="5985" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.33" />
                    <SPLIT distance="100" swimtime="00:01:43.62" />
                    <SPLIT distance="150" swimtime="00:02:32.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3886" number="1" />
                    <RELAYPOSITION athleteid="3858" number="2" reactiontime="+112" />
                    <RELAYPOSITION athleteid="3838" number="3" reactiontime="+88" />
                    <RELAYPOSITION athleteid="3867" number="4" reactiontime="+92" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1418" points="421" reactiontime="+93" swimtime="00:02:03.35" resultid="3914" heatid="5910" lane="6" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:34.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3847" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="3897" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3853" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3877" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="418" reactiontime="+87" swimtime="00:02:16.86" resultid="3915" heatid="5986" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3853" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3847" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3897" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3877" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="242" reactiontime="+76" swimtime="00:02:34.39" resultid="3909" heatid="5837" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:01:51.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3897" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3847" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3893" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="3883" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="215" reactiontime="+83" swimtime="00:02:40.59" resultid="3910" heatid="5837" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:08.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3886" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3838" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3843" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3870" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1229" points="388" reactiontime="+153" swimtime="00:02:11.91" resultid="3911" heatid="5837" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:01:43.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3853" number="1" reactiontime="+153" />
                    <RELAYPOSITION athleteid="3863" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3904" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3877" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4003" name="niezrzeszony" />
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="4887" name="UKS ,,Trójka&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="4888">
              <RESULTS>
                <RESULT eventid="1178" points="333" reactiontime="+88" swimtime="00:02:38.05" resultid="4889" heatid="5815" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:02:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="370" reactiontime="+82" swimtime="00:02:30.67" resultid="4890" heatid="5896" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="349" reactiontime="+77" swimtime="00:02:50.65" resultid="4891" heatid="5949" lane="4" entrytime="00:02:51.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:06.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4892" heatid="5982" lane="1" entrytime="00:05:06.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" clubid="2885" name="KS Masters Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Gizela" lastname="Wójcik" birthdate="1949-11-16" gender="F" nation="POL" athleteid="2891">
              <RESULTS>
                <RESULT eventid="1093" points="64" swimtime="00:02:35.31" resultid="2892" heatid="5785" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="51" reactiontime="+109" swimtime="00:01:08.86" resultid="2893" heatid="5798" lane="1" />
                <RESULT eventid="1247" points="35" swimtime="00:02:32.91" resultid="2894" heatid="5840" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="59" swimtime="00:01:13.04" resultid="2895" heatid="5860" lane="6" />
                <RESULT eventid="1451" points="34" swimtime="00:01:10.41" resultid="2896" heatid="5916" lane="0" />
                <RESULT eventid="1486" points="60" swimtime="00:05:43.25" resultid="2897" heatid="5942" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.05" />
                    <SPLIT distance="100" swimtime="00:02:42.59" />
                    <SPLIT distance="150" swimtime="00:04:12.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Marchlewski" birthdate="1957-09-11" gender="M" nation="POL" athleteid="2932">
              <RESULTS>
                <RESULT eventid="1110" points="113" reactiontime="+112" swimtime="00:01:54.44" resultid="2933" heatid="5789" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="58" reactiontime="+113" swimtime="00:04:16.11" resultid="2934" heatid="5827" lane="0">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:04:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="69" reactiontime="+105" swimtime="00:01:49.38" resultid="2935" heatid="5846" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="117" reactiontime="+104" swimtime="00:00:51.55" resultid="2936" heatid="5866" lane="6" />
                <RESULT eventid="1469" points="117" reactiontime="+92" swimtime="00:00:41.20" resultid="2937" heatid="5924" lane="3" />
                <RESULT eventid="1503" points="84" reactiontime="+88" swimtime="00:04:33.51" resultid="2938" heatid="5945" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.17" />
                    <SPLIT distance="100" swimtime="00:02:09.70" />
                    <SPLIT distance="150" swimtime="00:03:22.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Kawula" birthdate="1941-10-02" gender="F" nation="POL" athleteid="2886">
              <RESULTS>
                <RESULT eventid="1093" points="10" swimtime="00:04:41.41" resultid="2887" heatid="5784" lane="1" />
                <RESULT eventid="1247" points="15" swimtime="00:03:23.39" resultid="2888" heatid="5840" lane="0" />
                <RESULT eventid="1282" points="9" swimtime="00:02:14.79" resultid="2889" heatid="5860" lane="1" />
                <RESULT eventid="1451" points="17" swimtime="00:01:28.52" resultid="2890" heatid="5916" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zygmunt" lastname="Pawlaczek" birthdate="1949-05-26" gender="M" nation="POL" athleteid="2919">
              <RESULTS>
                <RESULT eventid="1110" points="126" reactiontime="+108" swimtime="00:01:50.15" resultid="2920" heatid="5789" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="101" reactiontime="+97" swimtime="00:03:33.04" resultid="2921" heatid="5826" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:39.43" />
                    <SPLIT distance="150" swimtime="00:02:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="123" reactiontime="+114" swimtime="00:01:30.16" resultid="2922" heatid="5846" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="86" reactiontime="+109" swimtime="00:01:51.36" resultid="2923" heatid="5882" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="144" reactiontime="+107" swimtime="00:00:38.40" resultid="2924" heatid="5924" lane="0" />
                <RESULT eventid="1605" points="97" swimtime="00:07:41.47" resultid="2925" heatid="5977" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:45.27" />
                    <SPLIT distance="200" swimtime="00:03:45.99" />
                    <SPLIT distance="300" swimtime="00:05:44.07" />
                    <SPLIT distance="350" swimtime="00:06:43.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Józefa" lastname="Wołoszczuk" birthdate="1953-01-23" gender="F" nation="POL" athleteid="2905">
              <RESULTS>
                <RESULT eventid="1127" points="34" reactiontime="+94" swimtime="00:01:18.75" resultid="2906" heatid="5797" lane="4" />
                <RESULT eventid="1195" points="40" reactiontime="+111" swimtime="00:05:20.39" resultid="2907" heatid="5821" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.24" />
                    <SPLIT distance="100" swimtime="00:02:35.94" />
                    <SPLIT distance="150" swimtime="00:03:58.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="42" reactiontime="+113" swimtime="00:02:24.00" resultid="2908" heatid="5840" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="26" reactiontime="+113" swimtime="00:03:09.59" resultid="2909" heatid="5876" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="42" reactiontime="+115" swimtime="00:01:05.61" resultid="2910" heatid="5915" lane="3" />
                <RESULT eventid="1520" points="37" reactiontime="+98" swimtime="00:02:43.63" resultid="2911" heatid="5951" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Regina" lastname="Mładszew" birthdate="1952-07-15" gender="F" nation="POL" athleteid="2912">
              <RESULTS>
                <RESULT eventid="1093" points="30" reactiontime="+126" swimtime="00:03:20.03" resultid="2913" heatid="5784" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="30" reactiontime="+188" swimtime="00:01:22.14" resultid="2914" heatid="5798" lane="0" />
                <RESULT eventid="1316" points="29" reactiontime="+129" swimtime="00:03:03.54" resultid="2915" heatid="5876" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="36" reactiontime="+109" swimtime="00:05:59.61" resultid="2916" heatid="5901" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.55" />
                    <SPLIT distance="150" swimtime="00:03:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="34" reactiontime="+112" swimtime="00:01:10.77" resultid="2917" heatid="5916" lane="6" />
                <RESULT eventid="1520" points="34" reactiontime="+149" swimtime="00:02:49.04" resultid="2918" heatid="5952" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pavlo" lastname="Vechirko" birthdate="1968-01-02" gender="M" nation="POL" athleteid="2926">
              <RESULTS>
                <RESULT eventid="1110" points="267" reactiontime="+88" swimtime="00:01:25.92" resultid="2927" heatid="5793" lane="5" entrytime="00:01:23.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="227" reactiontime="+76" swimtime="00:00:36.42" resultid="2928" heatid="5807" lane="7" entrytime="00:00:36.78" entrycourse="SCM" />
                <RESULT eventid="1299" points="278" reactiontime="+85" swimtime="00:00:38.67" resultid="2929" heatid="5870" lane="2" entrytime="00:00:38.30" entrycourse="SCM" />
                <RESULT eventid="1401" points="219" reactiontime="+76" swimtime="00:02:54.99" resultid="2930" heatid="5907" lane="0" entrytime="00:02:44.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:25.57" />
                    <SPLIT distance="150" swimtime="00:02:10.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="2931" heatid="5949" lane="1" entrytime="00:02:57.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janina" lastname="Zając" birthdate="1946-08-16" gender="F" nation="POL" athleteid="2898">
              <RESULTS>
                <RESULT eventid="1093" points="36" reactiontime="+122" swimtime="00:03:08.41" resultid="2899" heatid="5784" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="28" reactiontime="+103" swimtime="00:01:24.11" resultid="2900" heatid="5798" lane="2" />
                <RESULT eventid="1247" points="33" swimtime="00:02:35.19" resultid="2901" heatid="5839" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="34" swimtime="00:06:03.81" resultid="2902" heatid="5901" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.12" />
                    <SPLIT distance="150" swimtime="00:04:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="34" swimtime="00:01:10.42" resultid="2903" heatid="5915" lane="5" />
                <RESULT eventid="1520" points="29" reactiontime="+118" swimtime="00:02:57.72" resultid="2904" heatid="5951" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Jawor" birthdate="1947-04-23" gender="M" nation="POL" swrid="4754745" athleteid="2939">
              <RESULTS>
                <RESULT eventid="1144" points="47" reactiontime="+118" swimtime="00:01:01.48" resultid="2940" heatid="5803" lane="5" />
                <RESULT eventid="1212" points="57" reactiontime="+99" swimtime="00:04:17.17" resultid="2941" heatid="5827" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.95" />
                    <SPLIT distance="100" swimtime="00:03:12.42" />
                    <SPLIT distance="150" swimtime="00:04:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="62" reactiontime="+103" swimtime="00:01:53.32" resultid="2942" heatid="5845" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="50" reactiontime="+111" swimtime="00:04:46.02" resultid="2943" heatid="5904" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.85" />
                    <SPLIT distance="100" swimtime="00:02:19.43" />
                    <SPLIT distance="150" swimtime="00:03:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="77" reactiontime="+90" swimtime="00:00:47.19" resultid="2944" heatid="5923" lane="6" />
                <RESULT eventid="1537" points="44" reactiontime="+124" swimtime="00:02:16.28" resultid="2945" heatid="5957" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3313" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Modzelewski" birthdate="1984-01-01" gender="M" nation="POL" athleteid="3312">
              <RESULTS>
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach." eventid="1144" reactiontime="+76" status="DSQ" swimtime="00:00:00.00" resultid="3314" heatid="5804" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1299" points="222" reactiontime="+71" swimtime="00:00:41.70" resultid="3315" heatid="5868" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="4495" name="KU AZS Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Kister" birthdate="1989-01-01" gender="M" nation="POL" swrid="4992691" athleteid="4123">
              <RESULTS>
                <RESULT eventid="1076" points="395" reactiontime="+77" swimtime="00:00:29.62" resultid="4124" heatid="5779" lane="6" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1110" points="356" reactiontime="+77" swimtime="00:01:18.07" resultid="4125" heatid="5795" lane="9" entrytime="00:01:18.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="385" reactiontime="+78" swimtime="00:00:34.68" resultid="4126" heatid="5872" lane="1" entrytime="00:00:35.50" entrycourse="SCM" />
                <RESULT eventid="1367" points="301" reactiontime="+81" swimtime="00:02:41.34" resultid="4127" heatid="5899" lane="3" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="322" reactiontime="+75" swimtime="00:02:55.31" resultid="4128" heatid="5949" lane="2" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="326" reactiontime="+75" swimtime="00:01:09.38" resultid="4129" heatid="5969" lane="2" entrytime="00:01:08.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" license="508114700069" swrid="4251117" athleteid="4500">
              <RESULTS>
                <RESULT eventid="1265" points="574" reactiontime="+72" swimtime="00:00:54.06" resultid="4501" heatid="5857" lane="2" entrytime="00:00:55.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4502" heatid="5971" lane="9" entrytime="00:00:59.99" />
                <RESULT eventid="1212" points="512" reactiontime="+83" swimtime="00:02:04.14" resultid="5721" heatid="5828" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="100" swimtime="00:00:56.56" />
                    <SPLIT distance="150" swimtime="00:01:28.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-01-01" gender="M" nation="POL" swrid="4086676" athleteid="4130">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4131" heatid="5781" lane="3" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1265" points="549" reactiontime="+69" swimtime="00:00:54.88" resultid="4132" heatid="5858" lane="6" entrytime="00:00:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4133" heatid="5938" lane="0" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="5722" heatid="5810" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5723" heatid="5893" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5724" heatid="5971" lane="0" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Uziak" birthdate="1987-01-01" gender="M" nation="POL" athleteid="4134">
              <RESULTS>
                <RESULT eventid="1265" points="365" swimtime="00:01:02.87" resultid="4135" heatid="5855" lane="9" entrytime="00:01:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="368" reactiontime="+66" swimtime="00:00:28.13" resultid="4136" heatid="5934" lane="4" entrytime="00:00:27.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Godlewski" birthdate="1996-05-26" gender="M" nation="POL" license="108114700059" swrid="4285522" athleteid="4496">
              <RESULTS>
                <RESULT eventid="1110" points="486" reactiontime="+72" swimtime="00:01:10.35" resultid="4497" heatid="5796" lane="0" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="515" reactiontime="+69" swimtime="00:00:31.50" resultid="4498" heatid="5874" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1469" points="461" reactiontime="+71" swimtime="00:00:26.08" resultid="4499" heatid="5932" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="514" reactiontime="+71" swimtime="00:01:42.11" resultid="5725" heatid="5914" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.78" />
                    <SPLIT distance="100" swimtime="00:00:48.90" />
                    <SPLIT distance="150" swimtime="00:01:16.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4130" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4500" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4134" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4496" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01911" nation="POL" region="11" clubid="4735" name="Rybnicki Młodzieżowy Klub Sportowy">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" license="101911600104" swrid="4992966" athleteid="4736">
              <RESULTS>
                <RESULT eventid="1059" points="466" reactiontime="+72" swimtime="00:00:31.44" resultid="4737" heatid="5771" lane="8" entrytime="00:00:31.92" entrycourse="SCM" />
                <RESULT eventid="1127" points="339" reactiontime="+75" swimtime="00:00:36.69" resultid="4738" heatid="5801" lane="8" entrytime="00:00:37.16" entrycourse="SCM" />
                <RESULT eventid="1247" points="458" reactiontime="+72" swimtime="00:01:05.16" resultid="4739" heatid="5843" lane="5" entrytime="00:01:07.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="417" reactiontime="+82" swimtime="00:01:15.59" resultid="4740" heatid="5876" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="506" reactiontime="+69" swimtime="00:00:28.76" resultid="4741" heatid="5921" lane="2" entrytime="00:00:29.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3474" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Budziszewski" birthdate="1997-01-01" gender="M" nation="POL" swrid="4289414" athleteid="3473">
              <RESULTS>
                <RESULT eventid="1076" points="414" reactiontime="+67" swimtime="00:00:29.16" resultid="3475" heatid="5781" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1144" points="292" reactiontime="+64" swimtime="00:00:33.48" resultid="3476" heatid="5809" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1333" points="331" reactiontime="+73" swimtime="00:01:11.18" resultid="3477" heatid="5889" lane="9" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="383" reactiontime="+69" swimtime="00:00:27.74" resultid="3478" heatid="5935" lane="4" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" clubid="3230" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Beata" lastname="Jasko" birthdate="1955-10-10" gender="F" nation="POL" athleteid="3231">
              <RESULTS>
                <RESULT eventid="1093" points="143" reactiontime="+100" swimtime="00:01:59.02" resultid="3232" heatid="5785" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="183" reactiontime="+101" swimtime="00:00:50.28" resultid="3233" heatid="5859" lane="5" />
                <RESULT eventid="1316" points="102" swimtime="00:02:00.59" resultid="3234" heatid="5877" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Halina" lastname="Kaniewska" birthdate="1958-07-20" gender="F" nation="POL" athleteid="3258">
              <RESULTS>
                <RESULT eventid="1059" points="102" reactiontime="+129" swimtime="00:00:52.08" resultid="3259" heatid="5767" lane="1" />
                <RESULT eventid="1127" points="162" reactiontime="+94" swimtime="00:00:46.89" resultid="3260" heatid="5797" lane="5" />
                <RESULT eventid="1316" points="162" reactiontime="+117" swimtime="00:01:43.45" resultid="3261" heatid="5875" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="203" reactiontime="+101" swimtime="00:00:39.01" resultid="3262" heatid="5916" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Chmurski" birthdate="1987-09-23" gender="M" nation="POL" swrid="4060941" athleteid="3263">
              <RESULTS>
                <RESULT eventid="1212" points="462" reactiontime="+71" swimtime="00:02:08.54" resultid="3264" heatid="5835" lane="8" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="150" swimtime="00:01:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="436" reactiontime="+81" swimtime="00:01:04.94" resultid="3265" heatid="5892" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="501" reactiontime="+76" swimtime="00:00:25.37" resultid="3266" heatid="5939" lane="3" entrytime="00:00:24.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefania" lastname="Noetzel" birthdate="1935-08-21" gender="F" nation="POL" swrid="4791734" athleteid="3254">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1093" points="32" swimtime="00:03:14.80" resultid="3255" heatid="5785" lane="2" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1282" points="31" swimtime="00:01:30.48" resultid="3256" heatid="5860" lane="3" entrytime="00:01:23.62" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1486" points="37" swimtime="00:06:42.71" resultid="3257" heatid="5942" lane="7" entrytime="00:06:15.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.75" />
                    <SPLIT distance="100" swimtime="00:03:24.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Woźnicki" birthdate="1972-03-18" gender="M" nation="POL" swrid="4302597" athleteid="3267">
              <RESULTS>
                <RESULT eventid="1110" status="DNS" swimtime="00:00:00.00" resultid="3268" heatid="5790" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="1299" points="180" reactiontime="+87" swimtime="00:00:44.72" resultid="3269" heatid="5868" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Serbin" birthdate="1966-08-10" gender="F" nation="POL" swrid="4302596" athleteid="3243">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy od Rekordu Polski kat. G" eventid="1195" points="408" reactiontime="+74" swimtime="00:02:28.89" resultid="3244" heatid="5825" lane="1" entrytime="00:02:28.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy od Rekordu Polski kat. G" eventid="1247" points="386" reactiontime="+75" swimtime="00:01:08.99" resultid="3245" heatid="5843" lane="6" entrytime="00:01:08.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1588" points="437" reactiontime="+75" swimtime="00:05:08.22" resultid="3246" heatid="5975" lane="6" entrytime="00:05:06.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:52.64" />
                    <SPLIT distance="200" swimtime="00:02:31.71" />
                    <SPLIT distance="250" swimtime="00:03:11.15" />
                    <SPLIT distance="300" swimtime="00:03:50.20" />
                    <SPLIT distance="350" swimtime="00:04:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Grzeszewski" birthdate="1953-09-25" gender="M" nation="POL" swrid="4754656" athleteid="3235">
              <RESULTS>
                <RESULT eventid="1076" points="171" reactiontime="+93" swimtime="00:00:39.13" resultid="3236" heatid="5774" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1299" points="229" swimtime="00:00:41.26" resultid="3237" heatid="5869" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1503" points="165" swimtime="00:03:38.82" resultid="3238" heatid="5945" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                    <SPLIT distance="100" swimtime="00:01:45.74" />
                    <SPLIT distance="150" swimtime="00:02:44.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Kluczyk" birthdate="1987-02-27" gender="M" nation="POL" swrid="4967270" athleteid="3239">
              <RESULTS>
                <RESULT eventid="1178" points="307" reactiontime="+93" swimtime="00:02:42.51" resultid="3240" heatid="5818" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:02:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="219" swimtime="00:02:59.35" resultid="3241" heatid="5899" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:16.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="351" reactiontime="+88" swimtime="00:05:00.67" resultid="3242" heatid="5980" lane="0" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                    <SPLIT distance="200" swimtime="00:02:24.97" />
                    <SPLIT distance="250" swimtime="00:03:03.81" />
                    <SPLIT distance="300" swimtime="00:03:42.27" />
                    <SPLIT distance="350" swimtime="00:04:21.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03508" nation="POL" region="08" clubid="4341" name="Ks &quot;Prestige&quot;">
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Rupa" birthdate="1996-01-11" gender="F" nation="POL" license="103508600006" swrid="4108567" athleteid="4342">
              <RESULTS>
                <RESULT eventid="1059" points="386" reactiontime="+69" swimtime="00:00:33.48" resultid="4343" heatid="5766" lane="4" />
                <RESULT eventid="1127" points="454" reactiontime="+63" swimtime="00:00:33.29" resultid="4344" heatid="5802" lane="9" entrytime="00:00:33.88" entrycourse="SCM" />
                <RESULT eventid="1316" points="429" reactiontime="+54" swimtime="00:01:14.91" resultid="4345" heatid="5876" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="440" reactiontime="+55" swimtime="00:02:36.32" resultid="4346" heatid="5903" lane="6" entrytime="00:02:41.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" status="DNS" swimtime="00:00:00.00" resultid="4347" heatid="5920" lane="0" entrytime="00:00:31.36" />
                <RESULT eventid="1520" status="DNS" swimtime="00:00:00.00" resultid="4348" heatid="5955" lane="0" entrytime="00:01:15.53" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00612" nation="POL" region="12" clubid="4397" name="KS KSZO Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Sejmicki" birthdate="1961-05-04" gender="M" nation="POL" license="500612700426" athleteid="4398">
              <RESULTS>
                <RESULT eventid="1110" points="155" reactiontime="+99" swimtime="00:01:42.92" resultid="4399" heatid="5791" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="205" swimtime="00:00:42.81" resultid="4400" heatid="5868" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1469" points="165" reactiontime="+116" swimtime="00:00:36.72" resultid="4401" heatid="5926" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="1503" points="139" reactiontime="+107" swimtime="00:03:51.88" resultid="4402" heatid="5946" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.47" />
                    <SPLIT distance="100" swimtime="00:01:49.79" />
                    <SPLIT distance="150" swimtime="00:02:51.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Orłowski" birthdate="1960-02-26" gender="M" nation="POL" license="500612700404" athleteid="4403">
              <RESULTS>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1110" reactiontime="+87" status="DSQ" swimtime="00:00:00.00" resultid="4404" heatid="5789" lane="7" />
                <RESULT eventid="1144" points="78" reactiontime="+76" swimtime="00:00:51.85" resultid="4405" heatid="5803" lane="1" />
                <RESULT eventid="1299" points="139" reactiontime="+88" swimtime="00:00:48.66" resultid="4406" heatid="5867" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4407" heatid="5884" lane="2" entrytime="00:01:40.00" />
                <RESULT eventid="1469" points="133" reactiontime="+82" swimtime="00:00:39.41" resultid="4408" heatid="5925" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Żak" birthdate="1959-11-22" gender="M" nation="POL" license="500612700512" athleteid="4409">
              <RESULTS>
                <RESULT eventid="1144" points="129" reactiontime="+98" swimtime="00:00:43.95" resultid="4410" heatid="5805" lane="1" entrytime="00:00:44.00" />
                <RESULT eventid="1333" points="126" reactiontime="+112" swimtime="00:01:38.24" resultid="4411" heatid="5884" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="4412" heatid="5905" lane="9" entrytime="00:04:00.00" />
                <RESULT eventid="1469" points="191" swimtime="00:00:34.96" resultid="4413" heatid="5926" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="4414" heatid="5958" lane="2" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01304" nation="POL" region="04" clubid="4504" name="Landsberg Crew Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" license="501304700001" swrid="4432188" athleteid="2801">
              <RESULTS>
                <RESULT eventid="1178" points="453" reactiontime="+72" swimtime="00:02:22.66" resultid="2802" heatid="5820" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="499" swimtime="00:02:05.26" resultid="2803" heatid="5835" lane="6" entrytime="00:02:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:01.70" />
                    <SPLIT distance="150" swimtime="00:01:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="475" reactiontime="+73" swimtime="00:00:57.59" resultid="2804" heatid="5857" lane="3" entrytime="00:00:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="426" reactiontime="+77" swimtime="00:02:23.85" resultid="2805" heatid="5900" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="432" reactiontime="+75" swimtime="00:02:38.84" resultid="2806" heatid="5950" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="494" reactiontime="+70" swimtime="00:04:28.33" resultid="2807" heatid="5984" lane="2" entrytime="00:04:19.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:36.96" />
                    <SPLIT distance="200" swimtime="00:02:11.13" />
                    <SPLIT distance="250" swimtime="00:02:45.34" />
                    <SPLIT distance="300" swimtime="00:03:19.58" />
                    <SPLIT distance="350" swimtime="00:03:54.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Kaczmarek" birthdate="1992-08-23" gender="F" nation="POL" license="501304600002" athleteid="2794">
              <RESULTS>
                <RESULT eventid="1161" points="508" reactiontime="+73" swimtime="00:02:32.63" resultid="2795" heatid="5814" lane="4" entrytime="00:02:29.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="150" swimtime="00:01:56.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="480" reactiontime="+73" swimtime="00:02:20.98" resultid="2796" heatid="5825" lane="4" entrytime="00:02:14.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="578" reactiontime="+73" swimtime="00:01:00.30" resultid="2797" heatid="5844" lane="1" entrytime="00:01:01.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="573" reactiontime="+76" swimtime="00:01:08.01" resultid="2798" heatid="5881" lane="3" entrytime="00:01:08.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="562" reactiontime="+70" swimtime="00:00:27.78" resultid="2799" heatid="5921" lane="3" entrytime="00:00:28.23" />
                <RESULT eventid="1486" points="465" reactiontime="+79" swimtime="00:02:53.59" resultid="2800" heatid="5944" lane="4" entrytime="00:02:46.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                    <SPLIT distance="150" swimtime="00:02:08.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3514" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Bromberek" birthdate="1957-01-01" gender="M" nation="POL" athleteid="3513">
              <RESULTS>
                <RESULT eventid="1110" points="96" reactiontime="+107" swimtime="00:02:00.63" resultid="3515" heatid="5790" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3516" heatid="5804" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="3517" heatid="5867" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3518" heatid="5883" lane="6" entrytime="00:02:00.00" />
                <RESULT eventid="1469" points="159" reactiontime="+114" swimtime="00:00:37.14" resultid="3519" heatid="5927" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="3520" heatid="5957" lane="6" entrytime="00:02:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="4872" name="UKS ,,Jasień&apos;&apos; Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="4873">
              <RESULTS>
                <RESULT eventid="1093" points="382" swimtime="00:01:25.91" resultid="4874" heatid="5784" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="343" reactiontime="+98" swimtime="00:00:36.57" resultid="4875" heatid="5797" lane="2" />
                <RESULT eventid="1282" points="388" reactiontime="+91" swimtime="00:00:39.13" resultid="4876" heatid="5863" lane="3" entrytime="00:00:40.45" entrycourse="SCM" />
                <RESULT eventid="1316" points="378" swimtime="00:01:18.13" resultid="4877" heatid="5876" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="407" swimtime="00:00:30.92" resultid="4878" heatid="5920" lane="7" entrytime="00:00:31.08" entrycourse="SCM" />
                <RESULT eventid="1520" points="331" swimtime="00:01:19.35" resultid="4879" heatid="5952" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3117" name="JK Team Kraków">
          <ATHLETES>
            <ATHLETE firstname="Agata" lastname="Jasik" birthdate="1984-01-01" gender="F" nation="POL" swrid="5484408" athleteid="3125">
              <RESULTS>
                <RESULT eventid="1195" points="219" reactiontime="+86" swimtime="00:03:02.97" resultid="3126" heatid="5824" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:24.11" />
                    <SPLIT distance="150" swimtime="00:02:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="243" reactiontime="+74" swimtime="00:01:20.47" resultid="3127" heatid="5841" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Zając" birthdate="1984-01-01" gender="M" nation="POL" swrid="5468089" athleteid="3128">
              <RESULTS>
                <RESULT eventid="1076" points="151" reactiontime="+88" swimtime="00:00:40.82" resultid="3129" heatid="5775" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1265" points="169" reactiontime="+81" swimtime="00:01:21.21" resultid="3130" heatid="5849" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="143" reactiontime="+89" swimtime="00:01:34.07" resultid="3131" heatid="5884" lane="4" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szkudlarek" birthdate="1996-04-04" gender="F" nation="POL" swrid="4265739" athleteid="3118">
              <RESULTS>
                <RESULT eventid="1127" points="369" reactiontime="+71" swimtime="00:00:35.66" resultid="3119" heatid="5801" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1195" points="439" swimtime="00:02:25.23" resultid="3120" heatid="5825" lane="2" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="481" reactiontime="+74" swimtime="00:01:04.11" resultid="3121" heatid="5844" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="456" reactiontime="+63" swimtime="00:01:13.38" resultid="3122" heatid="5881" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="470" swimtime="00:00:29.48" resultid="3123" heatid="5922" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1520" points="374" reactiontime="+74" swimtime="00:01:16.18" resultid="3124" heatid="5955" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2778" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Trępała" birthdate="1965-01-01" gender="M" nation="POL" athleteid="2777">
              <RESULTS>
                <RESULT eventid="1076" points="40" reactiontime="+118" swimtime="00:01:03.09" resultid="2779" heatid="5775" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1212" points="54" reactiontime="+109" swimtime="00:04:22.88" resultid="2780" heatid="5829" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.25" />
                    <SPLIT distance="150" swimtime="00:03:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="63" reactiontime="+99" swimtime="00:00:50.64" resultid="2781" heatid="5928" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="2782" heatid="5978" lane="6" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06401" nation="POL" region="01" clubid="4349" name="KS &quot;Swimmers Centrum Ślęza&quot;">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Wolny" birthdate="1960-03-21" gender="M" nation="POL" license="506401700021" swrid="4183808" athleteid="4350">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1144" points="302" reactiontime="+71" swimtime="00:00:33.10" resultid="4351" heatid="5808" lane="3" entrytime="00:00:33.73" entrycourse="SCM" />
                <RESULT eventid="1178" points="341" reactiontime="+78" swimtime="00:02:36.87" resultid="4352" heatid="5815" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:02:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="313" reactiontime="+77" swimtime="00:01:12.56" resultid="4353" heatid="5889" lane="0" entrytime="00:01:13.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="286" reactiontime="+83" swimtime="00:02:40.25" resultid="4354" heatid="5904" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:19.21" />
                    <SPLIT distance="150" swimtime="00:02:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="304" reactiontime="+72" swimtime="00:01:11.81" resultid="4355" heatid="5961" lane="8" entrytime="00:01:11.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5378" name="5styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="5379">
              <RESULTS>
                <RESULT eventid="1212" points="340" reactiontime="+74" swimtime="00:02:22.36" resultid="5380" heatid="5833" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="337" reactiontime="+74" swimtime="00:01:04.55" resultid="5381" heatid="5853" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="330" reactiontime="+77" swimtime="00:00:29.17" resultid="5382" heatid="5933" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1605" points="327" swimtime="00:05:07.85" resultid="5383" heatid="5982" lane="9" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:50.45" />
                    <SPLIT distance="200" swimtime="00:02:29.30" />
                    <SPLIT distance="250" swimtime="00:03:08.54" />
                    <SPLIT distance="300" swimtime="00:03:48.11" />
                    <SPLIT distance="350" swimtime="00:04:28.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" clubid="2747" name="Ks Extreme Team Oborniki">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" swrid="4754624" athleteid="2748">
              <RESULTS>
                <RESULT comment="M7 - Pływak wykonał naprzemienne lub nierównoczesne ruchy nóg." eventid="1076" reactiontime="+84" status="DSQ" swimtime="00:00:00.00" resultid="2749" heatid="5773" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1212" points="106" reactiontime="+88" swimtime="00:03:29.93" resultid="2750" heatid="5829" lane="7" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:36.12" />
                    <SPLIT distance="150" swimtime="00:02:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="126" reactiontime="+90" swimtime="00:01:29.46" resultid="2751" heatid="5848" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="140" reactiontime="+96" swimtime="00:00:38.81" resultid="2752" heatid="5928" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1605" points="87" swimtime="00:07:58.91" resultid="2753" heatid="5978" lane="7" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:52.36" />
                    <SPLIT distance="150" swimtime="00:02:54.63" />
                    <SPLIT distance="200" swimtime="00:03:56.21" />
                    <SPLIT distance="250" swimtime="00:04:58.30" />
                    <SPLIT distance="300" swimtime="00:06:00.34" />
                    <SPLIT distance="350" swimtime="00:07:00.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3309" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Jerzykowski" birthdate="1987-01-01" gender="M" nation="POL" athleteid="3308">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3310" heatid="5774" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1367" points="101" reactiontime="+78" swimtime="00:03:51.97" resultid="3311" heatid="5898" lane="1" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:40.38" />
                    <SPLIT distance="150" swimtime="00:02:39.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3510" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Gawłowicz" birthdate="1987-01-01" gender="M" nation="POL" swrid="4037726" athleteid="3509">
              <RESULTS>
                <RESULT eventid="1076" points="526" reactiontime="+68" swimtime="00:00:26.94" resultid="3511" heatid="5783" lane="0" entrytime="00:00:26.80" />
                <RESULT eventid="1469" points="475" reactiontime="+70" swimtime="00:00:25.82" resultid="3512" heatid="5938" lane="4" entrytime="00:00:25.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3604" name="UKP Marlin">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Ekiert" birthdate="1984-02-18" gender="F" nation="POL" athleteid="3608">
              <RESULTS>
                <RESULT eventid="1451" points="155" reactiontime="+107" swimtime="00:00:42.66" resultid="3609" heatid="5915" lane="4" />
                <RESULT eventid="1520" points="129" reactiontime="+106" swimtime="00:01:48.50" resultid="3610" heatid="5952" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Bauer" birthdate="1963-04-08" gender="M" nation="POL" athleteid="3616">
              <RESULTS>
                <RESULT eventid="1110" status="DNS" swimtime="00:00:00.00" resultid="3617" heatid="5789" lane="2" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="3618" heatid="5826" lane="3" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="3619" heatid="5847" lane="0" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="3620" heatid="5865" lane="6" />
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="3621" heatid="5945" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Markiewicz" birthdate="1994-02-14" gender="F" nation="POL" athleteid="3605">
              <RESULTS>
                <RESULT eventid="1486" points="211" reactiontime="+75" swimtime="00:03:45.79" resultid="3606" heatid="5942" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                    <SPLIT distance="100" swimtime="00:01:49.78" />
                    <SPLIT distance="150" swimtime="00:02:47.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="149" reactiontime="+66" swimtime="00:01:42.78" resultid="3607" heatid="5963" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Kowalczyk" birthdate="1991-01-28" gender="F" nation="POL" athleteid="3622">
              <RESULTS>
                <RESULT eventid="1451" points="146" reactiontime="+95" swimtime="00:00:43.49" resultid="3623" heatid="5916" lane="3" />
                <RESULT eventid="1486" points="113" swimtime="00:04:37.82" resultid="3624" heatid="5942" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.85" />
                    <SPLIT distance="100" swimtime="00:02:07.11" />
                    <SPLIT distance="150" swimtime="00:03:22.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rosiak" birthdate="1973-03-16" gender="M" nation="POL" athleteid="3611">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="3612" heatid="5772" lane="7" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3613" heatid="5803" lane="8" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="3614" heatid="5866" lane="9" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3615" heatid="5883" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5109" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Kuśmider" birthdate="1989-01-01" gender="M" nation="POL" athleteid="5108">
              <RESULTS>
                <RESULT eventid="1469" points="290" reactiontime="+83" swimtime="00:00:30.44" resultid="5110" heatid="5930" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1605" points="327" reactiontime="+93" swimtime="00:05:07.86" resultid="5111" heatid="5980" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                    <SPLIT distance="200" swimtime="00:02:30.96" />
                    <SPLIT distance="250" swimtime="00:03:10.33" />
                    <SPLIT distance="300" swimtime="00:03:50.15" />
                    <SPLIT distance="350" swimtime="00:04:29.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3088" name="Masters Białystok">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Twarowski" birthdate="1965-05-24" gender="M" nation="POL" swrid="5125743" athleteid="3089">
              <RESULTS>
                <RESULT eventid="1144" points="194" reactiontime="+72" swimtime="00:00:38.34" resultid="3090" heatid="5806" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1212" points="184" reactiontime="+95" swimtime="00:02:54.63" resultid="3091" heatid="5830" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:23.51" />
                    <SPLIT distance="150" swimtime="00:02:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="109" reactiontime="+101" swimtime="00:03:46.44" resultid="3092" heatid="5898" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:47.65" />
                    <SPLIT distance="150" swimtime="00:02:48.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="183" reactiontime="+84" swimtime="00:03:06.05" resultid="3093" heatid="5906" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                    <SPLIT distance="150" swimtime="00:02:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="200" reactiontime="+74" swimtime="00:01:22.53" resultid="3094" heatid="5959" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="171" reactiontime="+102" swimtime="00:06:21.90" resultid="3095" heatid="5979" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:30.73" />
                    <SPLIT distance="150" swimtime="00:02:20.40" />
                    <SPLIT distance="200" swimtime="00:03:10.66" />
                    <SPLIT distance="250" swimtime="00:04:00.30" />
                    <SPLIT distance="300" swimtime="00:04:49.47" />
                    <SPLIT distance="350" swimtime="00:05:38.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5265" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Wilkosz" birthdate="1965-01-01" gender="M" nation="POL" athleteid="5264">
              <RESULTS>
                <RESULT eventid="1265" points="171" reactiontime="+84" swimtime="00:01:20.83" resultid="5267" heatid="5849" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="120" reactiontime="+84" swimtime="00:00:44.06" resultid="5426" heatid="5773" lane="6" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11514" nation="POL" region="14" clubid="4777" name="Stowarzyszenie Pływackie Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Fuliński" birthdate="1982-06-03" gender="M" nation="POL" license="111514700186" swrid="4992686" athleteid="4783">
              <RESULTS>
                <RESULT eventid="1265" points="477" reactiontime="+77" swimtime="00:00:57.49" resultid="4784" heatid="5856" lane="0" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="467" reactiontime="+79" swimtime="00:00:25.98" resultid="4785" heatid="5938" lane="8" entrytime="00:00:25.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Karczewski" birthdate="1974-07-07" gender="M" nation="POL" athleteid="3652">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="3653" heatid="5831" lane="9" entrytime="00:02:56.00" entrycourse="LCM" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="3654" heatid="5850" lane="8" entrytime="00:01:18.05" entrycourse="LCM" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="3655" heatid="5929" lane="0" entrytime="00:00:34.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łukasiuk" birthdate="1980-01-02" gender="F" nation="POL" license="511514600187" athleteid="4778">
              <RESULTS>
                <RESULT eventid="1093" points="323" reactiontime="+70" swimtime="00:01:30.86" resultid="4779" heatid="5787" lane="4" entrytime="00:01:32.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" status="DNS" swimtime="00:00:00.00" resultid="4780" heatid="5842" lane="7" entrytime="00:01:15.38" />
                <RESULT eventid="1282" points="355" reactiontime="+62" swimtime="00:00:40.33" resultid="4781" heatid="5863" lane="1" entrytime="00:00:42.60" />
                <RESULT eventid="1451" points="373" reactiontime="+69" swimtime="00:00:31.85" resultid="4782" heatid="5919" lane="5" entrytime="00:00:32.34" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03908" nation="POL" region="08" clubid="4786" name="Stowarzyszenie Sportowe SWIM TRI Rzeszów">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" license="503908700007" athleteid="4794">
              <RESULTS>
                <RESULT eventid="1212" points="433" reactiontime="+74" swimtime="00:02:11.34" resultid="4795" heatid="5834" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="436" reactiontime="+69" swimtime="00:00:59.23" resultid="4796" heatid="5856" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="443" reactiontime="+69" swimtime="00:00:26.44" resultid="4797" heatid="5936" lane="2" entrytime="00:00:26.90" />
                <RESULT eventid="1605" points="416" reactiontime="+72" swimtime="00:04:44.15" resultid="4798" heatid="5983" lane="1" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                    <SPLIT distance="200" swimtime="00:02:19.01" />
                    <SPLIT distance="250" swimtime="00:02:55.53" />
                    <SPLIT distance="300" swimtime="00:03:32.67" />
                    <SPLIT distance="350" swimtime="00:04:08.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-11-15" gender="M" nation="POL" license="503908700008" athleteid="4787">
              <RESULTS>
                <RESULT eventid="1076" points="306" reactiontime="+82" swimtime="00:00:32.25" resultid="4788" heatid="5777" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1144" points="223" reactiontime="+94" swimtime="00:00:36.59" resultid="4789" heatid="5807" lane="8" entrytime="00:00:37.50" />
                <RESULT eventid="1265" points="319" reactiontime="+83" swimtime="00:01:05.72" resultid="4790" heatid="5853" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="242" reactiontime="+80" swimtime="00:01:19.01" resultid="4791" heatid="5887" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="362" reactiontime="+81" swimtime="00:00:28.28" resultid="4792" heatid="5932" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1605" points="310" reactiontime="+82" swimtime="00:05:13.50" resultid="4793" heatid="5981" lane="8" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:51.66" />
                    <SPLIT distance="200" swimtime="00:02:32.23" />
                    <SPLIT distance="250" swimtime="00:03:13.07" />
                    <SPLIT distance="300" swimtime="00:03:53.68" />
                    <SPLIT distance="350" swimtime="00:04:34.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3928" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Bołtuć" birthdate="1983-01-01" gender="F" nation="POL" athleteid="3927">
              <RESULTS>
                <RESULT eventid="1161" points="223" reactiontime="+98" swimtime="00:03:20.75" resultid="3929" heatid="5813" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:37.93" />
                    <SPLIT distance="150" swimtime="00:02:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="283" swimtime="00:02:48.10" resultid="3930" heatid="5823" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:22.93" />
                    <SPLIT distance="150" swimtime="00:02:06.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="209" reactiontime="+89" swimtime="00:01:35.08" resultid="3931" heatid="5875" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="205" reactiontime="+121" swimtime="00:03:21.67" resultid="3932" heatid="5902" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:40.79" />
                    <SPLIT distance="150" swimtime="00:02:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="180" reactiontime="+122" swimtime="00:01:37.10" resultid="3933" heatid="5953" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="294" swimtime="00:05:51.47" resultid="3934" heatid="5974" lane="7" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:09.73" />
                    <SPLIT distance="200" swimtime="00:02:54.57" />
                    <SPLIT distance="250" swimtime="00:03:39.33" />
                    <SPLIT distance="300" swimtime="00:04:24.21" />
                    <SPLIT distance="350" swimtime="00:05:09.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3656" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="Roman" lastname="Zwierzyński" birthdate="1960-05-10" gender="M" nation="POL" athleteid="3704">
              <RESULTS>
                <RESULT eventid="1265" points="69" reactiontime="+123" swimtime="00:01:49.40" resultid="3705" heatid="5847" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="86" swimtime="00:00:57.14" resultid="3706" heatid="5867" lane="9" entrytime="00:00:59.00" />
                <RESULT eventid="1469" points="78" reactiontime="+97" swimtime="00:00:47.04" resultid="3707" heatid="5925" lane="8" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Daroch" birthdate="1956-12-06" gender="M" nation="POL" athleteid="3708">
              <RESULTS>
                <RESULT eventid="1299" points="76" reactiontime="+118" swimtime="00:00:59.49" resultid="3709" heatid="5866" lane="4" entrytime="00:00:59.00" />
                <RESULT eventid="1469" points="73" reactiontime="+113" swimtime="00:00:48.06" resultid="3710" heatid="5925" lane="0" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Michalczuk" birthdate="1970-03-05" gender="M" nation="POL" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1144" points="135" reactiontime="+69" swimtime="00:00:43.24" resultid="3695" heatid="5804" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="213" reactiontime="+87" swimtime="00:02:46.25" resultid="3696" heatid="5831" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="214" reactiontime="+84" swimtime="00:01:15.09" resultid="3697" heatid="5851" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3698" heatid="5884" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1469" points="252" reactiontime="+85" swimtime="00:00:31.91" resultid="3699" heatid="5929" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radosław" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" swrid="4429483" athleteid="3689">
              <RESULTS>
                <RESULT eventid="1110" points="282" reactiontime="+81" swimtime="00:01:24.31" resultid="3690" heatid="5793" lane="1" entrytime="00:01:26.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="3691" heatid="5832" lane="2" entrytime="00:02:38.00" />
                <RESULT eventid="1299" points="267" reactiontime="+86" swimtime="00:00:39.20" resultid="3692" heatid="5870" lane="6" entrytime="00:00:38.04" />
                <RESULT eventid="1503" points="256" reactiontime="+83" swimtime="00:03:09.08" resultid="3693" heatid="5948" lane="1" entrytime="00:03:07.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.38" />
                    <SPLIT distance="150" swimtime="00:02:19.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Bąkowski" birthdate="1984-06-20" gender="M" nation="POL" athleteid="3685">
              <RESULTS>
                <RESULT eventid="1144" points="279" reactiontime="+90" swimtime="00:00:33.97" resultid="3686" heatid="5808" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1333" points="278" reactiontime="+94" swimtime="00:01:15.47" resultid="3687" heatid="5888" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="280" reactiontime="+80" swimtime="00:01:13.85" resultid="3688" heatid="5960" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Burandt" birthdate="1972-12-15" gender="F" nation="POL" swrid="5471721" athleteid="3664">
              <RESULTS>
                <RESULT eventid="1059" points="274" reactiontime="+85" swimtime="00:00:37.53" resultid="3665" heatid="5769" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1195" points="271" reactiontime="+90" swimtime="00:02:50.45" resultid="3666" heatid="5823" lane="3" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="150" swimtime="00:02:07.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="280" reactiontime="+77" swimtime="00:01:16.77" resultid="3667" heatid="5842" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="292" reactiontime="+83" swimtime="00:00:34.54" resultid="3668" heatid="5918" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1588" points="246" swimtime="00:06:13.19" resultid="3669" heatid="5974" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:09.17" />
                    <SPLIT distance="200" swimtime="00:02:56.56" />
                    <SPLIT distance="250" swimtime="00:03:44.22" />
                    <SPLIT distance="300" swimtime="00:04:33.59" />
                    <SPLIT distance="350" swimtime="00:05:23.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Krowicka" birthdate="1960-05-11" gender="F" nation="POL" athleteid="3711">
              <RESULTS>
                <RESULT eventid="1093" points="209" reactiontime="+78" swimtime="00:01:45.08" resultid="3712" heatid="5786" lane="3" entrytime="00:01:48.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="224" reactiontime="+78" swimtime="00:00:47.02" resultid="3713" heatid="5862" lane="3" entrytime="00:00:45.72" />
                <RESULT eventid="1316" points="179" swimtime="00:01:40.23" resultid="3714" heatid="5877" lane="2" entrytime="00:01:40.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="188" swimtime="00:03:54.87" resultid="3715" heatid="5943" lane="7" entrytime="00:03:51.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                    <SPLIT distance="100" swimtime="00:01:51.92" />
                    <SPLIT distance="150" swimtime="00:02:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Chojcan" birthdate="1986-08-04" gender="F" nation="POL" athleteid="3657">
              <RESULTS>
                <RESULT eventid="1059" points="330" reactiontime="+71" swimtime="00:00:35.28" resultid="3658" heatid="5769" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1127" points="317" reactiontime="+66" swimtime="00:00:37.54" resultid="3659" heatid="5800" lane="3" entrytime="00:00:38.15" />
                <RESULT eventid="1350" points="254" reactiontime="+79" swimtime="00:03:08.68" resultid="3660" heatid="5895" lane="6" entrytime="00:03:23.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="150" swimtime="00:02:16.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="318" reactiontime="+74" swimtime="00:02:54.21" resultid="3661" heatid="5902" lane="5" entrytime="00:02:57.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:24.70" />
                    <SPLIT distance="150" swimtime="00:02:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="321" reactiontime="+74" swimtime="00:01:20.15" resultid="3662" heatid="5954" lane="8" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="292" reactiontime="+64" swimtime="00:01:22.27" resultid="3663" heatid="5964" lane="0" entrytime="00:01:23.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Podulka" birthdate="1975-09-29" gender="F" nation="POL" athleteid="3670">
              <RESULTS>
                <RESULT eventid="1059" points="250" reactiontime="+74" swimtime="00:00:38.68" resultid="3671" heatid="5769" lane="9" entrytime="00:00:42.29" />
                <RESULT eventid="1247" points="265" reactiontime="+74" swimtime="00:01:18.14" resultid="3672" heatid="5842" lane="9" entrytime="00:01:19.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="292" reactiontime="+68" swimtime="00:00:34.56" resultid="3673" heatid="5919" lane="8" entrytime="00:00:34.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Wawrzyńczak" birthdate="1990-09-11" gender="F" nation="POL" swrid="4071814" athleteid="3679">
              <RESULTS>
                <RESULT eventid="1059" points="379" swimtime="00:00:33.67" resultid="3680" heatid="5770" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1127" points="360" reactiontime="+74" swimtime="00:00:35.96" resultid="3681" heatid="5801" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1384" points="349" reactiontime="+70" swimtime="00:02:48.84" resultid="3682" heatid="5903" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:19.98" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="355" reactiontime="+72" swimtime="00:01:17.47" resultid="3683" heatid="5954" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="333" swimtime="00:01:18.75" resultid="3684" heatid="5964" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Chudoba" birthdate="1981-03-04" gender="M" nation="POL" athleteid="3700">
              <RESULTS>
                <RESULT eventid="1076" points="428" reactiontime="+78" swimtime="00:00:28.86" resultid="3701" heatid="5780" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1367" points="258" reactiontime="+92" swimtime="00:02:49.82" resultid="3702" heatid="5899" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:07.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="390" reactiontime="+81" swimtime="00:01:05.37" resultid="3703" heatid="5969" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Batóg" birthdate="1972-03-11" gender="F" nation="POL" athleteid="3674">
              <RESULTS>
                <RESULT eventid="1059" points="238" reactiontime="+69" swimtime="00:00:39.31" resultid="3675" heatid="5769" lane="8" entrytime="00:00:40.11" />
                <RESULT eventid="1316" points="279" reactiontime="+81" swimtime="00:01:26.40" resultid="3676" heatid="5878" lane="8" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="313" reactiontime="+78" swimtime="00:00:33.76" resultid="3677" heatid="5919" lane="0" entrytime="00:00:34.42" />
                <RESULT eventid="1554" points="231" reactiontime="+78" swimtime="00:01:28.97" resultid="3678" heatid="5963" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Swim Club Mastars Ślęza" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="285" reactiontime="+89" swimtime="00:02:04.29" resultid="3721" heatid="5912" lane="5" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:00:58.25" />
                    <SPLIT distance="150" swimtime="00:01:31.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3685" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3700" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3694" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="3689" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="307" reactiontime="+86" swimtime="00:02:13.94" resultid="3722" heatid="5988" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                    <SPLIT distance="150" swimtime="00:01:41.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3685" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3689" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3700" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="3694" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Swim Club Mastars Ślęza" number="1">
              <RESULTS>
                <RESULT eventid="1418" points="346" reactiontime="+70" swimtime="00:02:11.65" resultid="3719" heatid="5910" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:37.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3657" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3670" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3679" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3664" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="300" reactiontime="+76" swimtime="00:02:32.80" resultid="3720" heatid="5986" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:25.24" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3657" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3664" number="2" />
                    <RELAYPOSITION athleteid="3679" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3670" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Swim Club Mastars 1" number="1">
              <RESULTS>
                <RESULT eventid="1229" points="318" reactiontime="+85" swimtime="00:02:20.92" resultid="3716" heatid="5838" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="150" swimtime="00:01:49.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3685" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="3664" number="2" />
                    <RELAYPOSITION athleteid="3700" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Swim Club Mastars 2" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa)." eventid="1229" reactiontime="+75" status="DSQ" swimtime="00:00:00.00" resultid="3717" heatid="5837" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3674" number="1" reactiontime="+75" status="DSQ" />
                    <RELAYPOSITION athleteid="3689" number="2" reactiontime="-89" status="DSQ" />
                    <RELAYPOSITION athleteid="3679" number="3" reactiontime="-16" status="DSQ" />
                    <RELAYPOSITION athleteid="3694" number="4" reactiontime="+20" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Swim Club Mastars 3" number="3">
              <RESULTS>
                <RESULT eventid="1229" points="115" reactiontime="+117" swimtime="00:03:17.86" resultid="3718" heatid="5837" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.31" />
                    <SPLIT distance="100" swimtime="00:01:37.66" />
                    <SPLIT distance="150" swimtime="00:02:29.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3708" number="1" reactiontime="+117" />
                    <RELAYPOSITION athleteid="3711" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="3670" number="3" />
                    <RELAYPOSITION athleteid="3704" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3452" name="Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Grażyna" lastname="Heisler" birthdate="1951-01-01" gender="F" nation="POL" swrid="4191114" athleteid="3453">
              <RESULTS>
                <RESULT eventid="1059" points="71" reactiontime="+79" swimtime="00:00:58.65" resultid="3454" heatid="5767" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1127" points="86" reactiontime="+85" swimtime="00:00:57.80" resultid="3455" heatid="5799" lane="9" entrytime="00:01:00.00" />
                <RESULT eventid="1316" points="96" reactiontime="+96" swimtime="00:02:03.04" resultid="3456" heatid="5877" lane="8" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="148" reactiontime="+96" swimtime="00:00:43.26" resultid="3457" heatid="5917" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="1520" points="74" reactiontime="+78" swimtime="00:02:10.72" resultid="3458" heatid="5952" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" swrid="4302086" athleteid="3459">
              <RESULTS>
                <RESULT eventid="1110" points="64" reactiontime="+129" swimtime="00:02:17.94" resultid="3460" heatid="5790" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="42" reactiontime="+95" swimtime="00:01:03.66" resultid="3461" heatid="5804" lane="1" entrytime="00:01:03.00" />
                <RESULT eventid="1299" points="91" reactiontime="+123" swimtime="00:00:55.99" resultid="3462" heatid="5867" lane="8" entrytime="00:00:55.50" />
                <RESULT eventid="1333" points="40" swimtime="00:02:22.93" resultid="3463" heatid="5883" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="48" swimtime="00:00:55.31" resultid="3464" heatid="5925" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1537" points="34" reactiontime="+108" swimtime="00:02:28.90" resultid="3465" heatid="5957" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" clubid="5501" name="Mks Swim Academy Termy Jakuba Oława">
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Mruk" birthdate="1978-09-27" gender="F" nation="POL" license="104501600044" athleteid="5502">
              <RESULTS>
                <RESULT eventid="1059" points="410" reactiontime="+87" swimtime="00:00:32.81" resultid="5503" heatid="5770" lane="3" entrytime="00:00:33.90" />
                <RESULT eventid="1093" points="410" reactiontime="+77" swimtime="00:01:23.88" resultid="5504" heatid="5788" lane="8" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="433" reactiontime="+67" swimtime="00:00:37.73" resultid="5505" heatid="5864" lane="0" entrytime="00:00:38.80" />
                <RESULT eventid="1316" points="415" swimtime="00:01:15.75" resultid="5506" heatid="5880" lane="9" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3626" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Wiesław" lastname="Bar" birthdate="1970-01-01" gender="M" nation="POL" swrid="4992835" athleteid="3625">
              <RESULTS>
                <RESULT eventid="1144" points="259" reactiontime="+70" swimtime="00:00:34.85" resultid="3627" heatid="5807" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1212" points="350" swimtime="00:02:20.98" resultid="3628" heatid="5834" lane="9" entrytime="00:02:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:06.82" />
                    <SPLIT distance="150" swimtime="00:01:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="364" reactiontime="+68" swimtime="00:01:02.91" resultid="3629" heatid="5855" lane="8" entrytime="00:01:01.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="300" reactiontime="+83" swimtime="00:01:13.57" resultid="3630" heatid="5890" lane="0" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="361" reactiontime="+85" swimtime="00:00:28.30" resultid="3631" heatid="5934" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1605" points="338" reactiontime="+78" swimtime="00:05:04.45" resultid="3632" heatid="5982" lane="5" entrytime="00:04:54.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:47.24" />
                    <SPLIT distance="200" swimtime="00:02:26.14" />
                    <SPLIT distance="250" swimtime="00:03:05.22" />
                    <SPLIT distance="300" swimtime="00:03:45.38" />
                    <SPLIT distance="350" swimtime="00:04:25.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01201" nation="POL" region="01" clubid="4597" name="MKS Piast Głogów" />
        <CLUB type="CLUB" nation="POL" clubid="1655" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Grzelczak" birthdate="1985-01-01" gender="M" nation="POL" athleteid="1654">
              <RESULTS>
                <RESULT eventid="1110" points="213" reactiontime="+96" swimtime="00:01:32.65" resultid="1656" heatid="5791" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="126" reactiontime="+95" swimtime="00:03:17.95" resultid="1657" heatid="5830" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                    <SPLIT distance="100" swimtime="00:01:29.98" />
                    <SPLIT distance="150" swimtime="00:02:23.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="226" reactiontime="+92" swimtime="00:00:41.44" resultid="1658" heatid="5869" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1333" points="126" reactiontime="+99" swimtime="00:01:38.26" resultid="1659" heatid="5884" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="190" reactiontime="+93" swimtime="00:03:28.94" resultid="1660" heatid="5946" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:37.61" />
                    <SPLIT distance="150" swimtime="00:02:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="112" reactiontime="+104" swimtime="00:07:19.59" resultid="1661" heatid="5978" lane="3" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:33.91" />
                    <SPLIT distance="150" swimtime="00:02:28.40" />
                    <SPLIT distance="200" swimtime="00:03:27.21" />
                    <SPLIT distance="250" swimtime="00:04:26.43" />
                    <SPLIT distance="300" swimtime="00:05:25.14" />
                    <SPLIT distance="350" swimtime="00:06:24.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00304" nation="POL" region="04" clubid="4815" name="TP Zielona Góra">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Karczewski" birthdate="1974-06-11" gender="M" nation="POL" license="100304700490" swrid="5342868" athleteid="4816">
              <RESULTS>
                <RESULT eventid="1076" points="364" reactiontime="+77" swimtime="00:00:30.45" resultid="4817" heatid="5779" lane="2" entrytime="00:00:30.43" entrycourse="SCM" />
                <RESULT eventid="1265" points="347" swimtime="00:01:03.93" resultid="4818" heatid="5854" lane="9" entrytime="00:01:04.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="321" reactiontime="+77" swimtime="00:00:29.42" resultid="4819" heatid="5933" lane="2" entrytime="00:00:28.92" entrycourse="SCM" />
                <RESULT eventid="1571" points="264" reactiontime="+79" swimtime="00:01:14.44" resultid="4820" heatid="5967" lane="6" entrytime="00:01:16.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIKRA" nation="POL" clubid="5294" name="Stowarzyszenie SIEMACHA Kraków">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska - Latuszek" birthdate="1985-08-01" gender="F" nation="POL" license="503706600141" athleteid="5295">
              <RESULTS>
                <RESULT eventid="1059" points="355" reactiontime="+68" swimtime="00:00:34.41" resultid="5296" heatid="5768" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1127" points="394" reactiontime="+67" swimtime="00:00:34.90" resultid="5297" heatid="5801" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1316" points="408" reactiontime="+60" swimtime="00:01:16.19" resultid="5298" heatid="5880" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="395" reactiontime="+72" swimtime="00:02:42.07" resultid="5299" heatid="5903" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:01:59.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="402" reactiontime="+66" swimtime="00:00:31.06" resultid="5300" heatid="5920" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1520" points="380" swimtime="00:01:15.76" resultid="5301" heatid="5955" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" clubid="5094" name="KS. Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" athleteid="5095">
              <RESULTS>
                <RESULT eventid="1076" points="314" reactiontime="+82" swimtime="00:00:31.98" resultid="5096" heatid="5779" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1144" points="267" reactiontime="+69" swimtime="00:00:34.48" resultid="5097" heatid="5808" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1265" points="290" swimtime="00:01:07.88" resultid="5098" heatid="5854" lane="7" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="250" reactiontime="+84" swimtime="00:02:51.64" resultid="5099" heatid="5899" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="5100" heatid="5960" lane="0" entrytime="00:01:17.00" />
                <RESULT eventid="1571" points="299" reactiontime="+75" swimtime="00:01:11.39" resultid="5101" heatid="5968" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="4744" name="Stowarzyszenie Pływackie MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" athleteid="4752">
              <RESULTS>
                <RESULT eventid="1367" points="124" reactiontime="+101" swimtime="00:03:36.62" resultid="4756" heatid="5896" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.05" />
                    <SPLIT distance="100" swimtime="00:01:47.44" />
                    <SPLIT distance="150" swimtime="00:02:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="176" reactiontime="+97" swimtime="00:00:35.97" resultid="4757" heatid="5927" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pietrzak" birthdate="1988-10-21" gender="M" nation="POL" license="103503700011" athleteid="4771">
              <RESULTS>
                <RESULT eventid="1144" points="258" reactiontime="+74" swimtime="00:00:34.89" resultid="4772" heatid="5807" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1333" points="291" reactiontime="+74" swimtime="00:01:14.32" resultid="4773" heatid="5885" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="344" swimtime="00:00:28.77" resultid="4774" heatid="5932" lane="7" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Ćwikła" birthdate="1975-11-07" gender="M" nation="POL" license="103503700005" swrid="5241236" athleteid="4767">
              <RESULTS>
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="4768" heatid="5809" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4769" heatid="5887" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="4770" heatid="5956" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wójcicki" birthdate="1975-04-28" gender="M" nation="POL" license="103503700001" swrid="5455050" athleteid="4759">
              <RESULTS>
                <RESULT eventid="1110" points="240" reactiontime="+79" swimtime="00:01:28.95" resultid="4760" heatid="5789" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="244" reactiontime="+77" swimtime="00:00:40.40" resultid="4761" heatid="5866" lane="8" />
                <RESULT eventid="1537" points="230" reactiontime="+78" swimtime="00:01:18.83" resultid="4762" heatid="5956" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Wójcicka" birthdate="1975-05-28" gender="F" nation="POL" license="103503600002" athleteid="4763">
              <RESULTS>
                <RESULT eventid="1127" points="279" reactiontime="+77" swimtime="00:00:39.17" resultid="4764" heatid="5797" lane="6" />
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="4765" heatid="5875" lane="4" />
                <RESULT eventid="1520" points="258" reactiontime="+96" swimtime="00:01:26.20" resultid="4766" heatid="5952" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Kawecka" birthdate="1993-09-06" gender="F" nation="POL" license="103503600028" swrid="5118335" athleteid="4745">
              <RESULTS>
                <RESULT eventid="1059" points="251" swimtime="00:00:38.60" resultid="4746" heatid="5767" lane="2" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="4747" heatid="5798" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Dawidek" birthdate="1986-03-13" gender="M" nation="POL" license="103503700029" athleteid="4748">
              <RESULTS>
                <RESULT eventid="1076" points="352" swimtime="00:00:30.79" resultid="4749" heatid="5778" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1333" points="269" reactiontime="+77" swimtime="00:01:16.30" resultid="4750" heatid="5888" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="375" reactiontime="+78" swimtime="00:00:27.94" resultid="4751" heatid="5934" lane="8" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="291" reactiontime="+74" swimtime="00:02:03.38" resultid="4775" heatid="5912" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:35.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4759" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4752" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4771" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="4748" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2843" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Kamiński" birthdate="1965-01-01" gender="M" nation="POL" athleteid="2842">
              <RESULTS>
                <RESULT eventid="1144" points="200" reactiontime="+73" swimtime="00:00:37.96" resultid="2844" heatid="5805" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1212" points="228" reactiontime="+90" swimtime="00:02:42.46" resultid="2845" heatid="5830" lane="4" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:01:59.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="233" reactiontime="+82" swimtime="00:01:13.03" resultid="2846" heatid="5850" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="214" swimtime="00:01:22.30" resultid="2847" heatid="5887" lane="9" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="217" reactiontime="+82" swimtime="00:00:33.53" resultid="2848" heatid="5930" lane="8" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11314" nation="POL" region="14" clubid="3419" name="Fundacja HASTEN">
          <ATHLETES>
            <ATHLETE firstname="Adrianna" lastname="Niewiadomska" birthdate="1999-12-28" gender="F" nation="POL" swrid="4359123" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1247" points="515" reactiontime="+74" swimtime="00:01:02.69" resultid="3433" heatid="5844" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="481" reactiontime="+79" swimtime="00:01:12.12" resultid="3434" heatid="5881" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="575" reactiontime="+67" swimtime="00:00:27.56" resultid="3435" heatid="5922" lane="2" entrytime="00:00:26.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Patrzyk-Grabińska" birthdate="1978-12-13" gender="F" nation="POL" athleteid="3447">
              <RESULTS>
                <RESULT eventid="1059" points="187" reactiontime="+80" swimtime="00:00:42.61" resultid="3448" heatid="5769" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1451" points="234" reactiontime="+82" swimtime="00:00:37.20" resultid="3449" heatid="5918" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Bochyńska-Knapik" birthdate="1990-06-10" gender="F" nation="POL" swrid="4061587" athleteid="3420">
              <RESULTS>
                <RESULT eventid="1127" points="490" reactiontime="+67" swimtime="00:00:32.46" resultid="3421" heatid="5802" lane="6" entrytime="00:00:31.80" />
                <RESULT eventid="1316" points="421" reactiontime="+71" swimtime="00:01:15.39" resultid="3422" heatid="5881" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Napieraj" birthdate="1998-08-13" gender="M" nation="POL" swrid="4282149" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1144" points="536" reactiontime="+63" swimtime="00:00:27.35" resultid="3441" heatid="5811" lane="3" entrytime="00:00:27.20" />
                <RESULT eventid="1178" points="505" reactiontime="+74" swimtime="00:02:17.64" resultid="3442" heatid="5820" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="100" swimtime="00:01:04.18" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="504" reactiontime="+70" swimtime="00:01:01.91" resultid="3443" heatid="5893" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="449" reactiontime="+65" swimtime="00:02:17.85" resultid="3444" heatid="5908" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="531" reactiontime="+69" swimtime="00:00:59.65" resultid="3445" heatid="5962" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="463" reactiontime="+70" swimtime="00:04:34.30" resultid="3446" heatid="5984" lane="0" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:01:00.69" />
                    <SPLIT distance="150" swimtime="00:01:33.11" />
                    <SPLIT distance="200" swimtime="00:02:07.21" />
                    <SPLIT distance="250" swimtime="00:02:42.98" />
                    <SPLIT distance="300" swimtime="00:03:19.91" />
                    <SPLIT distance="350" swimtime="00:03:57.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Pawlaczek" birthdate="1993-01-04" gender="F" nation="POL" swrid="4072670" athleteid="3423">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1059" reactiontime="+55" status="DSQ" swimtime="00:00:00.00" resultid="3424" heatid="5771" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1247" points="629" reactiontime="+77" swimtime="00:00:58.63" resultid="3425" heatid="5844" lane="3" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="619" reactiontime="+72" swimtime="00:00:26.90" resultid="3426" heatid="5922" lane="6" entrytime="00:00:26.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirela" lastname="Olczak" birthdate="1993-02-20" gender="F" nation="POL" swrid="4087182" athleteid="3427">
              <RESULTS>
                <RESULT eventid="1059" points="537" swimtime="00:00:29.98" resultid="3428" heatid="5771" lane="2" entrytime="00:00:29.99" />
                <RESULT eventid="1161" points="500" reactiontime="+64" swimtime="00:02:33.53" resultid="3429" heatid="5814" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="536" swimtime="00:01:09.55" resultid="3430" heatid="5881" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="548" reactiontime="+68" swimtime="00:01:06.73" resultid="3431" heatid="5964" lane="4" entrytime="00:01:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Żarnowska" birthdate="1999-11-11" gender="F" nation="POL" swrid="4359262" athleteid="3436">
              <RESULTS>
                <RESULT eventid="1195" points="399" reactiontime="+71" swimtime="00:02:30.00" resultid="3437" heatid="5825" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="450" reactiontime="+67" swimtime="00:00:29.91" resultid="3438" heatid="5922" lane="0" entrytime="00:00:27.90" />
                <RESULT eventid="1588" points="384" reactiontime="+69" swimtime="00:05:21.73" resultid="3439" heatid="5975" lane="3" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:50.55" />
                    <SPLIT distance="200" swimtime="00:02:31.84" />
                    <SPLIT distance="250" swimtime="00:03:13.72" />
                    <SPLIT distance="300" swimtime="00:03:56.69" />
                    <SPLIT distance="350" swimtime="00:04:40.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="HASTEN Swimming Team" number="1">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1418" points="441" reactiontime="+67" swimtime="00:02:01.49" resultid="3450" heatid="5910" lane="4" entrytime="00:01:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="100" swimtime="00:01:05.04" />
                    <SPLIT distance="150" swimtime="00:01:35.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3427" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3447" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3420" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3423" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="461" reactiontime="+70" swimtime="00:02:12.44" resultid="3451" heatid="5986" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:36.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3420" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="3427" number="2" reactiontime="+7" />
                    <RELAYPOSITION athleteid="3423" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3447" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3317" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Reszka" birthdate="1989-01-01" gender="M" nation="POL" athleteid="3316">
              <RESULTS>
                <RESULT eventid="1144" points="124" reactiontime="+86" swimtime="00:00:44.49" resultid="3318" heatid="5806" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1265" points="132" reactiontime="+80" swimtime="00:01:28.16" resultid="3319" heatid="5848" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5291" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Szot" birthdate="1995-01-01" gender="M" nation="POL" athleteid="5290">
              <RESULTS>
                <RESULT eventid="1110" points="504" reactiontime="+70" swimtime="00:01:09.50" resultid="5292" heatid="5795" lane="5" entrytime="00:01:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="530" reactiontime="+72" swimtime="00:00:31.20" resultid="5293" heatid="5873" lane="4" entrytime="00:00:31.99" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="4387" name="KS JUST SWIM Jelenia Góra">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-06-16" gender="F" nation="POL" license="505201600088" swrid="5435203" athleteid="4394">
              <RESULTS>
                <RESULT eventid="1350" points="170" reactiontime="+98" swimtime="00:03:35.52" resultid="4395" heatid="5895" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:42.13" />
                    <SPLIT distance="150" swimtime="00:02:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="265" reactiontime="+87" swimtime="00:06:03.89" resultid="4396" heatid="5974" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:01:22.19" />
                    <SPLIT distance="150" swimtime="00:02:07.78" />
                    <SPLIT distance="200" swimtime="00:02:54.41" />
                    <SPLIT distance="250" swimtime="00:03:41.31" />
                    <SPLIT distance="300" swimtime="00:04:28.86" />
                    <SPLIT distance="350" swimtime="00:05:16.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="219" reactiontime="+100" swimtime="00:03:22.10" resultid="5757" heatid="5812" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                    <SPLIT distance="100" swimtime="00:01:42.13" />
                    <SPLIT distance="150" swimtime="00:02:36.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-06-05" gender="M" nation="POL" license="505201700087" swrid="5435204" athleteid="4388">
              <RESULTS>
                <RESULT eventid="1076" points="155" reactiontime="+84" swimtime="00:00:40.49" resultid="4389" heatid="5775" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1212" points="157" reactiontime="+88" swimtime="00:03:03.99" resultid="4390" heatid="5830" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:27.97" />
                    <SPLIT distance="150" swimtime="00:02:16.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="106" reactiontime="+93" swimtime="00:03:48.61" resultid="4391" heatid="5898" lane="0" entrytime="00:03:53.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                    <SPLIT distance="100" swimtime="00:01:50.71" />
                    <SPLIT distance="150" swimtime="00:02:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="127" reactiontime="+88" swimtime="00:01:34.93" resultid="4392" heatid="5966" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="146" reactiontime="+91" swimtime="00:06:42.33" resultid="4393" heatid="5979" lane="5" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:30.66" />
                    <SPLIT distance="150" swimtime="00:02:20.66" />
                    <SPLIT distance="200" swimtime="00:03:11.70" />
                    <SPLIT distance="250" swimtime="00:04:03.95" />
                    <SPLIT distance="300" swimtime="00:04:55.86" />
                    <SPLIT distance="350" swimtime="00:05:51.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5370" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Ewelina" lastname="Cuch" birthdate="1979-01-01" gender="F" nation="POL" athleteid="5369">
              <RESULTS>
                <RESULT eventid="1059" points="316" reactiontime="+85" swimtime="00:00:35.79" resultid="5371" heatid="5767" lane="3" />
                <RESULT eventid="1093" points="305" reactiontime="+84" swimtime="00:01:32.56" resultid="5372" heatid="5785" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="306" swimtime="00:00:42.37" resultid="5373" heatid="5860" lane="7" />
                <RESULT eventid="1350" reactiontime="+83" status="DNF" swimtime="00:00:00.00" resultid="5374" heatid="5894" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="290" reactiontime="+67" swimtime="00:03:23.12" resultid="5375" heatid="5942" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                    <SPLIT distance="100" swimtime="00:01:37.60" />
                    <SPLIT distance="150" swimtime="00:02:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="261" reactiontime="+75" swimtime="00:01:25.44" resultid="5376" heatid="5963" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMT" nation="POL" clubid="3021" name="Toruń Multisport Team">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Lietz" birthdate="1952-04-23" gender="M" nation="POL" swrid="4754688" athleteid="3034">
              <RESULTS>
                <RESULT eventid="1212" points="160" reactiontime="+79" swimtime="00:03:02.96" resultid="3035" heatid="5830" lane="0" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                    <SPLIT distance="100" swimtime="00:01:29.57" />
                    <SPLIT distance="150" swimtime="00:02:18.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="198" swimtime="00:01:16.99" resultid="3036" heatid="5850" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="158" reactiontime="+68" swimtime="00:00:46.62" resultid="3037" heatid="5868" lane="0" entrytime="00:00:46.00" />
                <RESULT eventid="1469" points="206" reactiontime="+81" swimtime="00:00:34.11" resultid="3038" heatid="5928" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Gołembiewski" birthdate="1986-10-28" gender="M" nation="POL" athleteid="3039">
              <RESULTS>
                <RESULT eventid="1110" points="484" reactiontime="+82" swimtime="00:01:10.45" resultid="3040" heatid="5795" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="456" reactiontime="+81" swimtime="00:02:09.04" resultid="3041" heatid="5834" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="150" swimtime="00:01:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="496" reactiontime="+80" swimtime="00:00:31.89" resultid="3042" heatid="5873" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1333" points="375" swimtime="00:01:08.31" resultid="3043" heatid="5890" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="402" reactiontime="+87" swimtime="00:02:42.70" resultid="3044" heatid="5950" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="429" swimtime="00:04:41.36" resultid="3045" heatid="5983" lane="7" entrytime="00:04:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="150" swimtime="00:01:41.17" />
                    <SPLIT distance="200" swimtime="00:02:17.31" />
                    <SPLIT distance="250" swimtime="00:02:53.81" />
                    <SPLIT distance="300" swimtime="00:03:30.45" />
                    <SPLIT distance="350" swimtime="00:04:06.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Korolko" birthdate="1940-10-13" gender="M" nation="POL" swrid="4754683" athleteid="3060">
              <RESULTS>
                <RESULT eventid="1144" points="40" reactiontime="+85" swimtime="00:01:04.77" resultid="3061" heatid="5804" lane="8" entrytime="00:01:08.20" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="3062" heatid="5847" lane="4" entrytime="00:01:51.15" />
                <RESULT eventid="1401" points="28" reactiontime="+90" swimtime="00:05:45.20" resultid="3063" heatid="5904" lane="2" entrytime="00:05:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.07" />
                    <SPLIT distance="100" swimtime="00:02:43.59" />
                    <SPLIT distance="150" swimtime="00:04:14.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="85" reactiontime="+109" swimtime="00:00:45.68" resultid="3064" heatid="5925" lane="5" entrytime="00:00:44.61" />
                <RESULT eventid="1537" points="31" reactiontime="+82" swimtime="00:02:33.01" resultid="3065" heatid="5957" lane="3" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Bantkowski" birthdate="1949-08-24" gender="M" nation="POL" swrid="4754679" athleteid="3053">
              <RESULTS>
                <RESULT eventid="1178" points="16" swimtime="00:07:10.38" resultid="3054" heatid="5816" lane="9" entrytime="00:05:20.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.03" />
                    <SPLIT distance="100" swimtime="00:03:42.18" />
                    <SPLIT distance="150" swimtime="00:05:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="3055" heatid="5828" lane="2" entrytime="00:03:58.20" />
                <RESULT eventid="1367" status="DNS" swimtime="00:00:00.00" resultid="3056" heatid="5897" lane="8" entrytime="00:04:45.15" />
                <RESULT eventid="1401" points="11" reactiontime="+104" swimtime="00:07:43.38" resultid="3057" heatid="5904" lane="3" entrytime="00:04:20.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.22" />
                    <SPLIT distance="100" swimtime="00:03:50.24" />
                    <SPLIT distance="150" swimtime="00:05:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="7" reactiontime="+120" swimtime="00:04:05.32" resultid="3058" heatid="5965" lane="6" entrytime="00:03:29.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="3059" heatid="5977" lane="6" entrytime="00:09:31.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Marchewka" birthdate="1981-02-04" gender="M" nation="POL" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1144" points="335" reactiontime="+75" swimtime="00:00:31.97" resultid="3047" heatid="5803" lane="0" />
                <RESULT eventid="1178" points="389" reactiontime="+75" swimtime="00:02:30.14" resultid="3048" heatid="5818" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="424" reactiontime="+78" swimtime="00:01:05.56" resultid="3049" heatid="5882" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="3050" heatid="5907" lane="9" entrytime="00:02:45.00" />
                <RESULT eventid="1469" points="461" swimtime="00:00:26.08" resultid="3051" heatid="5925" lane="9" />
                <RESULT eventid="1537" points="378" reactiontime="+68" swimtime="00:01:06.82" resultid="3052" heatid="5960" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Kordowski" birthdate="1997-10-11" gender="M" nation="POL" athleteid="3022">
              <RESULTS>
                <RESULT eventid="1076" points="408" reactiontime="+74" swimtime="00:00:29.32" resultid="3023" heatid="5779" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1265" points="409" reactiontime="+75" swimtime="00:01:00.52" resultid="3024" heatid="5855" lane="4" entrytime="00:00:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="417" reactiontime="+73" swimtime="00:00:26.97" resultid="3025" heatid="5937" lane="0" entrytime="00:00:26.40" />
                <RESULT eventid="1571" points="302" swimtime="00:01:11.19" resultid="3026" heatid="5968" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucyna" lastname="Serożyńska" birthdate="1955-06-29" gender="F" nation="POL" swrid="5469132" athleteid="3066">
              <RESULTS>
                <RESULT eventid="1195" points="75" reactiontime="+115" swimtime="00:04:20.72" resultid="3067" heatid="5822" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.94" />
                    <SPLIT distance="100" swimtime="00:02:06.53" />
                    <SPLIT distance="150" swimtime="00:03:15.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="107" reactiontime="+118" swimtime="00:01:00.10" resultid="3068" heatid="5861" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1384" points="71" reactiontime="+108" swimtime="00:04:46.33" resultid="3069" heatid="5901" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.62" />
                    <SPLIT distance="100" swimtime="00:02:21.68" />
                    <SPLIT distance="150" swimtime="00:03:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="66" reactiontime="+94" swimtime="00:02:15.52" resultid="3070" heatid="5952" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="83" reactiontime="+124" swimtime="00:08:55.82" resultid="3071" heatid="5973" lane="0" entrytime="00:08:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.69" />
                    <SPLIT distance="150" swimtime="00:03:15.44" />
                    <SPLIT distance="200" swimtime="00:04:24.29" />
                    <SPLIT distance="250" swimtime="00:05:33.86" />
                    <SPLIT distance="300" swimtime="00:06:43.59" />
                    <SPLIT distance="350" swimtime="00:07:52.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Arentewicz" birthdate="1981-03-07" gender="M" nation="POL" swrid="4754686" athleteid="3072">
              <RESULTS>
                <RESULT eventid="1076" points="306" reactiontime="+72" swimtime="00:00:32.25" resultid="3073" heatid="5777" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1212" points="254" reactiontime="+78" swimtime="00:02:36.75" resultid="3074" heatid="5831" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="3075" heatid="5851" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1333" points="237" reactiontime="+79" swimtime="00:01:19.59" resultid="3076" heatid="5886" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="278" reactiontime="+77" swimtime="00:00:30.88" resultid="3077" heatid="5931" lane="1" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Lisiecki" birthdate="1982-01-28" gender="M" nation="POL" swrid="5469119" athleteid="3027">
              <RESULTS>
                <RESULT eventid="1178" points="277" reactiontime="+98" swimtime="00:02:48.10" resultid="3028" heatid="5817" lane="4" entrytime="00:02:58.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="263" reactiontime="+93" swimtime="00:02:34.97" resultid="3029" heatid="5832" lane="6" entrytime="00:02:33.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="242" swimtime="00:01:19.07" resultid="3030" heatid="5888" lane="9" entrytime="00:01:19.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="246" reactiontime="+84" swimtime="00:02:48.42" resultid="3031" heatid="5906" lane="4" entrytime="00:02:46.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:05.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="212" reactiontime="+86" swimtime="00:01:21.04" resultid="3032" heatid="5960" lane="9" entrytime="00:01:18.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="269" swimtime="00:05:28.61" resultid="3033" heatid="5981" lane="7" entrytime="00:05:25.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:01:59.36" />
                    <SPLIT distance="200" swimtime="00:02:41.35" />
                    <SPLIT distance="250" swimtime="00:03:22.81" />
                    <SPLIT distance="300" swimtime="00:04:05.07" />
                    <SPLIT distance="350" swimtime="00:04:47.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" status="DNS" swimtime="00:00:00.00" resultid="3078" heatid="5913" lane="5" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3046" number="1" />
                    <RELAYPOSITION athleteid="3027" number="2" />
                    <RELAYPOSITION athleteid="3072" number="3" />
                    <RELAYPOSITION athleteid="3039" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="3079" heatid="5989" lane="0" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3046" number="1" />
                    <RELAYPOSITION athleteid="3039" number="2" />
                    <RELAYPOSITION athleteid="3072" number="3" />
                    <RELAYPOSITION athleteid="3027" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" clubid="5203" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Jankowiak" birthdate="1981-12-27" gender="M" nation="POL" athleteid="5213">
              <RESULTS>
                <RESULT eventid="1076" points="265" reactiontime="+67" swimtime="00:00:33.85" resultid="5214" heatid="5777" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1265" points="300" reactiontime="+68" swimtime="00:01:07.07" resultid="5215" heatid="5852" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="324" swimtime="00:00:29.35" resultid="5216" heatid="5932" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kaczmarek" birthdate="1983-07-27" gender="M" nation="POL" athleteid="5208">
              <RESULTS>
                <RESULT eventid="1144" points="244" reactiontime="+85" swimtime="00:00:35.54" resultid="5209" heatid="5808" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1265" points="338" reactiontime="+75" swimtime="00:01:04.50" resultid="5210" heatid="5853" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="350" reactiontime="+71" swimtime="00:00:28.58" resultid="5211" heatid="5932" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1537" points="242" reactiontime="+84" swimtime="00:01:17.52" resultid="5212" heatid="5959" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Bernaś" birthdate="1984-02-13" gender="M" nation="POL" athleteid="5204">
              <RESULTS>
                <RESULT eventid="1076" points="324" reactiontime="+69" swimtime="00:00:31.64" resultid="5205" heatid="5779" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1265" points="349" reactiontime="+72" swimtime="00:01:03.79" resultid="5206" heatid="5855" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="364" reactiontime="+73" swimtime="00:00:28.23" resultid="5207" heatid="5936" lane="9" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Niewitecki" birthdate="1959-07-12" gender="M" nation="POL" athleteid="5217">
              <RESULTS>
                <RESULT eventid="1144" points="160" reactiontime="+82" swimtime="00:00:40.90" resultid="5218" heatid="5807" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1333" points="157" reactiontime="+93" swimtime="00:01:31.28" resultid="5219" heatid="5886" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="153" reactiontime="+84" swimtime="00:01:30.32" resultid="5220" heatid="5959" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="311" reactiontime="+94" swimtime="00:02:00.64" resultid="5221" heatid="5913" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5217" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="5208" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="5213" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="5204" number="4" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="281" reactiontime="+81" swimtime="00:02:17.94" resultid="5222" heatid="5988" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5217" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5213" number="2" />
                    <RELAYPOSITION athleteid="5204" number="3" />
                    <RELAYPOSITION athleteid="5208" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" clubid="4013" name="Korona Kraków Masters">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" swrid="5484421" athleteid="4027">
              <RESULTS>
                <RESULT eventid="1110" points="173" reactiontime="+90" swimtime="00:01:39.20" resultid="4028" heatid="5790" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="171" reactiontime="+74" swimtime="00:00:45.41" resultid="4029" heatid="5866" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="1367" points="94" reactiontime="+72" swimtime="00:03:57.35" resultid="4030" heatid="5897" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                    <SPLIT distance="100" swimtime="00:01:46.87" />
                    <SPLIT distance="150" swimtime="00:02:48.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="187" reactiontime="+85" swimtime="00:03:29.97" resultid="4031" heatid="5946" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.42" />
                    <SPLIT distance="100" swimtime="00:01:44.31" />
                    <SPLIT distance="150" swimtime="00:02:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="100" reactiontime="+77" swimtime="00:01:42.80" resultid="4032" heatid="5966" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" swrid="4992907" athleteid="4102">
              <RESULTS>
                <RESULT eventid="1127" points="333" swimtime="00:00:36.93" resultid="4103" heatid="5801" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1316" points="366" reactiontime="+80" swimtime="00:01:18.97" resultid="4104" heatid="5878" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="299" reactiontime="+73" swimtime="00:02:57.78" resultid="4105" heatid="5903" lane="1" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="314" reactiontime="+71" swimtime="00:01:20.70" resultid="4106" heatid="5955" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Łysiak" birthdate="1973-03-30" gender="M" nation="POL" swrid="5468085" athleteid="4021">
              <RESULTS>
                <RESULT eventid="1110" points="311" reactiontime="+77" swimtime="00:01:21.63" resultid="4022" heatid="5793" lane="4" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="280" swimtime="00:02:47.41" resultid="4023" heatid="5818" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:07.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="4024" heatid="5852" lane="7" entrytime="00:01:08.00" />
                <RESULT eventid="1299" points="293" reactiontime="+75" swimtime="00:00:38.00" resultid="4025" heatid="5870" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1503" points="297" reactiontime="+89" swimtime="00:03:00.06" resultid="4026" heatid="5949" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:27.80" />
                    <SPLIT distance="150" swimtime="00:02:14.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Borek" birthdate="1991-01-01" gender="M" nation="POL" swrid="5468079" athleteid="4074">
              <RESULTS>
                <RESULT eventid="1144" points="274" reactiontime="+70" swimtime="00:00:34.19" resultid="4075" heatid="5808" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1299" points="323" swimtime="00:00:36.78" resultid="4076" heatid="5865" lane="7" />
                <RESULT eventid="1333" points="327" reactiontime="+66" swimtime="00:01:11.52" resultid="4077" heatid="5888" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="296" reactiontime="+67" swimtime="00:01:12.44" resultid="4078" heatid="5960" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" swrid="4218717" athleteid="4061">
              <RESULTS>
                <RESULT eventid="1127" points="219" reactiontime="+78" swimtime="00:00:42.42" resultid="4062" heatid="5799" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1195" points="239" swimtime="00:02:57.77" resultid="4063" heatid="5823" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                    <SPLIT distance="100" swimtime="00:01:29.23" />
                    <SPLIT distance="150" swimtime="00:02:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="254" swimtime="00:01:19.29" resultid="4064" heatid="5841" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="214" reactiontime="+95" swimtime="00:01:34.42" resultid="4065" heatid="5877" lane="4" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="172" reactiontime="+85" swimtime="00:01:38.69" resultid="4066" heatid="5953" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="225" reactiontime="+108" swimtime="00:06:24.11" resultid="4067" heatid="5973" lane="6" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                    <SPLIT distance="200" swimtime="00:03:10.61" />
                    <SPLIT distance="250" swimtime="00:04:00.59" />
                    <SPLIT distance="300" swimtime="00:04:51.13" />
                    <SPLIT distance="350" swimtime="00:05:39.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Orlewicz-Musiał" birthdate="1960-05-29" gender="F" nation="POL" swrid="5352178" athleteid="4107">
              <RESULTS>
                <RESULT eventid="1093" points="74" reactiontime="+97" swimtime="00:02:28.19" resultid="4108" heatid="5785" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="74" reactiontime="+107" swimtime="00:04:50.17" resultid="4109" heatid="5812" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.01" />
                    <SPLIT distance="100" swimtime="00:02:16.39" />
                    <SPLIT distance="150" swimtime="00:03:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="80" reactiontime="+100" swimtime="00:01:06.22" resultid="4110" heatid="5859" lane="3" />
                <RESULT eventid="1316" points="77" reactiontime="+89" swimtime="00:02:12.55" resultid="4111" heatid="5876" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="64" swimtime="00:02:17.10" resultid="4112" heatid="5951" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="83" reactiontime="+89" swimtime="00:08:55.95" resultid="4113" heatid="5972" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.45" />
                    <SPLIT distance="100" swimtime="00:02:00.70" />
                    <SPLIT distance="150" swimtime="00:03:08.46" />
                    <SPLIT distance="200" swimtime="00:04:17.09" />
                    <SPLIT distance="250" swimtime="00:05:26.46" />
                    <SPLIT distance="300" swimtime="00:06:37.95" />
                    <SPLIT distance="350" swimtime="00:07:48.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Mleczko" birthdate="1946-10-22" gender="F" nation="POL" swrid="4992813" athleteid="4090">
              <RESULTS>
                <RESULT eventid="1093" points="32" reactiontime="+121" swimtime="00:03:15.03" resultid="4091" heatid="5785" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="17" reactiontime="+83" swimtime="00:01:38.97" resultid="4092" heatid="5798" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="1247" points="26" reactiontime="+120" swimtime="00:02:48.11" resultid="4093" heatid="5840" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="45" reactiontime="+110" swimtime="00:01:19.99" resultid="4094" heatid="5860" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="1451" points="28" reactiontime="+106" swimtime="00:01:14.95" resultid="4095" heatid="5916" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1520" points="16" reactiontime="+71" swimtime="00:03:33.71" resultid="4096" heatid="5952" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" swrid="4992827" athleteid="4054">
              <RESULTS>
                <RESULT eventid="1059" points="221" swimtime="00:00:40.31" resultid="4055" heatid="5769" lane="2" entrytime="00:00:39.00" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1195" points="289" reactiontime="+100" swimtime="00:02:46.90" resultid="4056" heatid="5824" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="287" reactiontime="+91" swimtime="00:01:16.17" resultid="4057" heatid="5842" lane="0" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="201" reactiontime="+91" swimtime="00:03:23.87" resultid="4058" heatid="5895" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:34.11" />
                    <SPLIT distance="150" swimtime="00:02:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="289" swimtime="00:00:34.65" resultid="4059" heatid="5919" lane="1" entrytime="00:00:34.00" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1554" points="216" reactiontime="+90" swimtime="00:01:30.92" resultid="4060" heatid="5963" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska" birthdate="1984-04-20" gender="F" nation="POL" swrid="5468078" athleteid="4097">
              <RESULTS>
                <RESULT eventid="1093" points="94" swimtime="00:02:16.83" resultid="4098" heatid="5785" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="84" reactiontime="+123" swimtime="00:00:58.27" resultid="4099" heatid="5798" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1282" points="94" swimtime="00:01:02.62" resultid="4100" heatid="5860" lane="4" entrytime="00:01:20.00" />
                <RESULT eventid="1486" points="95" swimtime="00:04:54.74" resultid="4101" heatid="5942" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.33" />
                    <SPLIT distance="100" swimtime="00:02:26.21" />
                    <SPLIT distance="150" swimtime="00:03:42.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-03-21" gender="M" nation="POL" swrid="4992712" athleteid="4047">
              <RESULTS>
                <RESULT eventid="1110" points="236" reactiontime="+101" swimtime="00:01:29.44" resultid="4048" heatid="5792" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="246" reactiontime="+89" swimtime="00:02:38.39" resultid="4049" heatid="5832" lane="7" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="293" reactiontime="+85" swimtime="00:01:07.59" resultid="4050" heatid="5852" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="219" reactiontime="+92" swimtime="00:01:21.65" resultid="4051" heatid="5886" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="273" reactiontime="+88" swimtime="00:00:31.04" resultid="4052" heatid="5930" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1503" points="226" reactiontime="+99" swimtime="00:03:17.05" resultid="4053" heatid="5947" lane="3" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                    <SPLIT distance="100" swimtime="00:01:34.05" />
                    <SPLIT distance="150" swimtime="00:02:25.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Jośko" birthdate="1994-07-25" gender="M" nation="POL" swrid="5484409" athleteid="4079">
              <RESULTS>
                <RESULT comment="K15 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu." eventid="1110" reactiontime="+66" status="DSQ" swimtime="00:00:00.00" resultid="4080" heatid="5793" lane="8" entrytime="00:01:26.91" />
                <RESULT eventid="1265" points="344" reactiontime="+67" swimtime="00:01:04.08" resultid="4081" heatid="5852" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="348" reactiontime="+69" swimtime="00:00:35.89" resultid="4082" heatid="5871" lane="3" entrytime="00:00:36.02" />
                <RESULT eventid="1469" points="351" reactiontime="+67" swimtime="00:00:28.57" resultid="4083" heatid="5932" lane="4" entrytime="00:00:29.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mleczko" birthdate="1947-08-26" gender="M" nation="POL" swrid="4992812" athleteid="4033">
              <RESULTS>
                <RESULT eventid="1076" points="94" reactiontime="+121" swimtime="00:00:47.76" resultid="4034" heatid="5774" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1212" points="148" reactiontime="+120" swimtime="00:03:07.71" resultid="4035" heatid="5829" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:31.18" />
                    <SPLIT distance="150" swimtime="00:02:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="173" reactiontime="+133" swimtime="00:01:20.56" resultid="4036" heatid="5850" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="41" reactiontime="+126" swimtime="00:05:13.61" resultid="4037" heatid="5897" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.36" />
                    <SPLIT distance="100" swimtime="00:02:17.26" />
                    <SPLIT distance="150" swimtime="00:03:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="187" reactiontime="+131" swimtime="00:00:35.24" resultid="4038" heatid="5929" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1571" points="60" reactiontime="+128" swimtime="00:02:01.48" resultid="4039" heatid="5966" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" swrid="4992797" athleteid="4014">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1059" points="377" reactiontime="+75" swimtime="00:00:33.73" resultid="4015" heatid="5770" lane="7" entrytime="00:00:34.50" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1127" points="345" reactiontime="+67" swimtime="00:00:36.48" resultid="4016" heatid="5801" lane="0" entrytime="00:00:37.50" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1282" points="421" reactiontime="+75" swimtime="00:00:38.09" resultid="4017" heatid="5864" lane="8" entrytime="00:00:38.70" entrycourse="SCM" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski, Czas Lepszy Od Rekordu Polski" eventid="1316" points="381" reactiontime="+71" swimtime="00:01:17.92" resultid="4018" heatid="5880" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Czas Lepszy od Rekordu Polski" eventid="1451" points="407" reactiontime="+71" swimtime="00:00:30.93" resultid="4019" heatid="5920" lane="1" entrytime="00:00:31.10" />
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1520" points="328" reactiontime="+67" swimtime="00:01:19.52" resultid="4020" heatid="5954" lane="3" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" swrid="4992740" athleteid="4068">
              <RESULTS>
                <RESULT eventid="1076" points="444" reactiontime="+70" swimtime="00:00:28.50" resultid="4069" heatid="5781" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1299" points="395" reactiontime="+70" swimtime="00:00:34.39" resultid="4070" heatid="5872" lane="4" entrytime="00:00:34.33" entrycourse="SCM" />
                <RESULT eventid="1333" points="336" reactiontime="+74" swimtime="00:01:10.85" resultid="4071" heatid="5890" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="441" reactiontime="+72" swimtime="00:00:26.48" resultid="4072" heatid="5935" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4073" heatid="5969" lane="7" entrytime="00:01:09.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Waga" birthdate="1940-07-04" gender="M" nation="POL" swrid="4992823" athleteid="4084">
              <RESULTS>
                <RESULT eventid="1212" points="60" swimtime="00:04:12.66" resultid="4085" heatid="5827" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.27" />
                    <SPLIT distance="100" swimtime="00:02:04.70" />
                    <SPLIT distance="150" swimtime="00:03:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="65" swimtime="00:01:51.48" resultid="4086" heatid="5847" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="40" reactiontime="+105" swimtime="00:01:13.35" resultid="4087" heatid="5866" lane="0" />
                <RESULT eventid="1469" points="74" reactiontime="+107" swimtime="00:00:47.96" resultid="4088" heatid="5923" lane="4" />
                <RESULT eventid="1605" points="66" swimtime="00:08:44.78" resultid="4089" heatid="5977" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.45" />
                    <SPLIT distance="100" swimtime="00:02:05.95" />
                    <SPLIT distance="150" swimtime="00:03:11.95" />
                    <SPLIT distance="200" swimtime="00:04:19.03" />
                    <SPLIT distance="250" swimtime="00:05:27.43" />
                    <SPLIT distance="300" swimtime="00:06:35.82" />
                    <SPLIT distance="350" swimtime="00:07:42.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Piszczek" birthdate="1962-11-10" gender="M" nation="POL" swrid="4992814" athleteid="4040">
              <RESULTS>
                <RESULT eventid="1076" points="331" reactiontime="+86" swimtime="00:00:31.44" resultid="4041" heatid="5778" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1144" points="236" reactiontime="+82" swimtime="00:00:35.93" resultid="4042" heatid="5807" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1299" points="318" reactiontime="+87" swimtime="00:00:36.96" resultid="4043" heatid="5871" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1401" points="243" reactiontime="+168" swimtime="00:02:49.22" resultid="4044" heatid="5906" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:22.89" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="242" reactiontime="+82" swimtime="00:01:17.45" resultid="4045" heatid="5960" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4046" heatid="5968" lane="0" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT comment="O11 - Pływak przeszkadzał innemu zawodnikowi (przez wpłynięcie na tor zajmowany przez innego zawodnika lub w inny sposób)." eventid="1442" reactiontime="+70" status="DSQ" swimtime="00:00:00.00" resultid="4117" heatid="5912" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                    <SPLIT distance="100" swimtime="00:00:57.90" />
                    <SPLIT distance="150" swimtime="00:01:32.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4068" number="1" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="4047" number="2" reactiontime="+61" status="DSQ" />
                    <RELAYPOSITION athleteid="4033" number="3" reactiontime="+47" status="DSQ" />
                    <RELAYPOSITION athleteid="4040" number="4" reactiontime="+21" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="4120" heatid="5988" lane="1" entrytime="00:02:19.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4074" number="1" />
                    <RELAYPOSITION athleteid="4079" number="2" />
                    <RELAYPOSITION athleteid="4021" number="3" />
                    <RELAYPOSITION athleteid="4027" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="291" reactiontime="+67" swimtime="00:02:03.32" resultid="4119" heatid="5913" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:00:59.48" />
                    <SPLIT distance="150" swimtime="00:01:35.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4074" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4021" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4027" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="4079" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1646" points="272" reactiontime="+73" swimtime="00:02:19.44" resultid="4121" heatid="5988" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:01:43.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4040" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4047" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4068" number="3" />
                    <RELAYPOSITION athleteid="4033" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT comment="Czas Lepszy Od Rekordu Polski" eventid="1418" points="354" reactiontime="+78" swimtime="00:02:10.74" resultid="4115" heatid="5910" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:02.59" />
                    <SPLIT distance="150" swimtime="00:01:36.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4014" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="4102" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="4061" number="3" />
                    <RELAYPOSITION athleteid="4054" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1622" points="334" reactiontime="+60" swimtime="00:02:27.53" resultid="4116" heatid="5986" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:15.60" />
                    <SPLIT distance="150" swimtime="00:01:52.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4102" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4014" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4061" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="4054" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1229" points="290" reactiontime="+71" swimtime="00:02:25.22" resultid="4114" heatid="5837" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="150" swimtime="00:01:50.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4102" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4047" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="4040" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4061" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1229" points="289" reactiontime="+95" swimtime="00:02:25.45" resultid="4118" heatid="5838" lane="9" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:01:49.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4054" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="4014" number="2" />
                    <RELAYPOSITION athleteid="4068" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4033" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="4160" name="Stowarzyszenie Pływackie Masters Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Lemańczyk" birthdate="1977-01-01" gender="M" nation="POL" athleteid="5102">
              <RESULTS>
                <RESULT eventid="1110" points="195" reactiontime="+114" swimtime="00:01:35.27" resultid="5103" heatid="5790" lane="3" entrytime="00:01:45.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="173" reactiontime="+82" swimtime="00:02:58.00" resultid="5104" heatid="5829" lane="3" entrytime="00:03:17.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:11.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="167" swimtime="00:01:21.47" resultid="5105" heatid="5849" lane="9" entrytime="00:01:27.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="176" reactiontime="+81" swimtime="00:00:35.97" resultid="5106" heatid="5926" lane="1" entrytime="00:00:42.00" />
                <RESULT eventid="1605" points="164" reactiontime="+98" swimtime="00:06:27.18" resultid="5107" heatid="5976" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:18.00" />
                    <SPLIT distance="200" swimtime="00:03:07.27" />
                    <SPLIT distance="250" swimtime="00:03:57.92" />
                    <SPLIT distance="300" swimtime="00:04:48.34" />
                    <SPLIT distance="350" swimtime="00:05:38.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kieres" birthdate="1984-06-13" gender="M" nation="POL" license="101713700001" swrid="5282844" athleteid="4180">
              <RESULTS>
                <RESULT eventid="1076" points="274" reactiontime="+69" swimtime="00:00:33.45" resultid="4181" heatid="5778" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1110" points="290" reactiontime="+73" swimtime="00:01:23.56" resultid="4182" heatid="5794" lane="5" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="285" swimtime="00:00:38.36" resultid="4183" heatid="5872" lane="9" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1367" points="247" reactiontime="+78" swimtime="00:02:52.34" resultid="4184" heatid="5899" lane="8" entrytime="00:02:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="4185" heatid="5949" lane="0" entrytime="00:02:58.00" entrycourse="SCM" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="4186" heatid="5967" lane="5" entrytime="00:01:15.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-02-10" gender="M" nation="POL" license="101713700005" swrid="4062177" athleteid="4206">
              <RESULTS>
                <RESULT eventid="1076" points="686" reactiontime="+70" swimtime="00:00:24.66" resultid="4207" heatid="5783" lane="5" entrytime="00:00:24.35" entrycourse="SCM" />
                <RESULT eventid="1265" points="643" swimtime="00:00:52.06" resultid="4208" heatid="5858" lane="5" entrytime="00:00:51.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4209" heatid="5940" lane="6" entrytime="00:00:23.34" entrycourse="SCM" />
                <RESULT eventid="1571" points="606" reactiontime="+67" swimtime="00:00:56.45" resultid="4210" heatid="5971" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Łuczak" birthdate="1978-03-18" gender="M" nation="POL" license="501713700016" swrid="5416815" athleteid="4217">
              <RESULTS>
                <RESULT eventid="1110" points="340" reactiontime="+70" swimtime="00:01:19.26" resultid="4218" heatid="5794" lane="8" entrytime="00:01:20.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="376" reactiontime="+70" swimtime="00:00:34.98" resultid="4219" heatid="5872" lane="3" entrytime="00:00:34.82" entrycourse="SCM" />
                <RESULT eventid="1469" points="360" reactiontime="+65" swimtime="00:00:28.32" resultid="4220" heatid="5934" lane="5" entrytime="00:00:27.90" entrycourse="SCM" />
                <RESULT eventid="1503" points="303" reactiontime="+71" swimtime="00:02:58.79" resultid="4221" heatid="5949" lane="8" entrytime="00:02:57.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Gregorowicz" birthdate="1974-10-30" gender="M" nation="POL" license="101713700002" swrid="4992729" athleteid="4168">
              <RESULTS>
                <RESULT eventid="1076" points="483" reactiontime="+70" swimtime="00:00:27.72" resultid="4169" heatid="5772" lane="8" />
                <RESULT eventid="1212" points="476" reactiontime="+68" swimtime="00:02:07.22" resultid="4170" heatid="5835" lane="0" entrytime="00:02:07.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="464" reactiontime="+66" swimtime="00:02:19.76" resultid="4171" heatid="5900" lane="7" entrytime="00:02:20.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:08.09" />
                    <SPLIT distance="150" swimtime="00:01:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="459" reactiontime="+66" swimtime="00:00:26.12" resultid="4172" heatid="5938" lane="5" entrytime="00:00:25.38" entrycourse="SCM" />
                <RESULT eventid="1605" points="490" reactiontime="+71" swimtime="00:04:29.16" resultid="4173" heatid="5983" lane="5" entrytime="00:04:30.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:38.69" />
                    <SPLIT distance="200" swimtime="00:02:12.61" />
                    <SPLIT distance="250" swimtime="00:02:46.90" />
                    <SPLIT distance="300" swimtime="00:03:21.24" />
                    <SPLIT distance="350" swimtime="00:03:55.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Matusiak vel Matuszewski" birthdate="1974-06-25" gender="M" nation="POL" license="501713700004" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1076" points="154" swimtime="00:00:40.50" resultid="4200" heatid="5775" lane="2" entrytime="00:00:38.05" />
                <RESULT eventid="1144" points="151" reactiontime="+78" swimtime="00:00:41.69" resultid="4201" heatid="5806" lane="3" entrytime="00:00:39.92" />
                <RESULT eventid="1265" points="217" reactiontime="+83" swimtime="00:01:14.75" resultid="4202" heatid="5851" lane="2" entrytime="00:01:11.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="138" reactiontime="+90" swimtime="00:03:24.19" resultid="4203" heatid="5906" lane="9" entrytime="00:03:11.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="220" reactiontime="+77" swimtime="00:00:33.37" resultid="4204" heatid="5930" lane="2" entrytime="00:00:32.37" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="4205" heatid="5959" lane="0" entrytime="00:01:29.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Stępień" birthdate="1983-09-29" gender="M" nation="POL" license="501713700010" athleteid="4187">
              <RESULTS>
                <RESULT eventid="1076" points="264" reactiontime="+97" swimtime="00:00:33.88" resultid="4188" heatid="5776" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1212" points="319" reactiontime="+84" swimtime="00:02:25.30" resultid="4189" heatid="5832" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="347" reactiontime="+83" swimtime="00:01:03.94" resultid="4190" heatid="5852" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="311" reactiontime="+77" swimtime="00:00:29.75" resultid="4191" heatid="5933" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1605" points="272" reactiontime="+91" swimtime="00:05:27.44" resultid="4192" heatid="5981" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:55.64" />
                    <SPLIT distance="200" swimtime="00:02:37.87" />
                    <SPLIT distance="250" swimtime="00:03:20.32" />
                    <SPLIT distance="300" swimtime="00:04:03.62" />
                    <SPLIT distance="350" swimtime="00:04:46.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Gozdan" birthdate="1968-08-16" gender="M" nation="POL" license="501713700009" swrid="5230704" athleteid="4193">
              <RESULTS>
                <RESULT eventid="1076" points="146" reactiontime="+87" swimtime="00:00:41.28" resultid="4194" heatid="5775" lane="7" entrytime="00:00:38.93" entrycourse="SCM" />
                <RESULT eventid="1110" points="206" reactiontime="+87" swimtime="00:01:33.59" resultid="4195" heatid="5792" lane="1" entrytime="00:01:32.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="194" reactiontime="+88" swimtime="00:01:17.61" resultid="4196" heatid="5849" lane="4" entrytime="00:01:19.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="229" reactiontime="+89" swimtime="00:00:41.26" resultid="4197" heatid="5868" lane="3" entrytime="00:00:42.60" entrycourse="SCM" />
                <RESULT eventid="1469" points="211" swimtime="00:00:33.82" resultid="4198" heatid="5929" lane="7" entrytime="00:00:33.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Dąbrowski" birthdate="1974-01-14" gender="M" nation="POL" license="501713700022" swrid="5355776" athleteid="4174">
              <RESULTS>
                <RESULT eventid="1076" points="312" reactiontime="+79" swimtime="00:00:32.06" resultid="4175" heatid="5776" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1212" points="334" swimtime="00:02:23.16" resultid="4176" heatid="5833" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="323" reactiontime="+75" swimtime="00:01:05.47" resultid="4177" heatid="5852" lane="6" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="242" reactiontime="+90" swimtime="00:02:49.46" resultid="4178" heatid="5906" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:08.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="312" reactiontime="+80" swimtime="00:05:12.63" resultid="4179" heatid="5981" lane="6" entrytime="00:05:18.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                    <SPLIT distance="200" swimtime="00:02:34.23" />
                    <SPLIT distance="250" swimtime="00:03:14.37" />
                    <SPLIT distance="300" swimtime="00:03:54.44" />
                    <SPLIT distance="350" swimtime="00:04:34.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Koźlikowski" birthdate="1961-09-09" gender="M" nation="POL" license="501713700011" swrid="4992727" athleteid="4211">
              <RESULTS>
                <RESULT eventid="1110" points="236" reactiontime="+94" swimtime="00:01:29.50" resultid="4212" heatid="5791" lane="6" entrytime="00:01:36.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="208" swimtime="00:03:04.78" resultid="4213" heatid="5817" lane="7" entrytime="00:03:06.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:31.07" />
                    <SPLIT distance="150" swimtime="00:02:22.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="200" swimtime="00:01:24.14" resultid="4214" heatid="5886" lane="7" entrytime="00:01:25.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="205" reactiontime="+99" swimtime="00:03:23.50" resultid="4215" heatid="5947" lane="1" entrytime="00:03:22.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                    <SPLIT distance="100" swimtime="00:01:38.32" />
                    <SPLIT distance="150" swimtime="00:02:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="226" reactiontime="+98" swimtime="00:05:48.10" resultid="4216" heatid="5979" lane="4" entrytime="00:05:55.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:04.92" />
                    <SPLIT distance="200" swimtime="00:02:49.93" />
                    <SPLIT distance="250" swimtime="00:03:35.12" />
                    <SPLIT distance="300" swimtime="00:04:20.81" />
                    <SPLIT distance="350" swimtime="00:05:05.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Konopacki" birthdate="1978-04-01" gender="M" nation="POL" license="501713700019" swrid="5282843" athleteid="4222">
              <RESULTS>
                <RESULT eventid="1144" points="319" swimtime="00:00:32.49" resultid="4223" heatid="5803" lane="7" />
                <RESULT eventid="1212" points="423" reactiontime="+69" swimtime="00:02:12.36" resultid="4224" heatid="5834" lane="1" entrytime="00:02:14.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="400" reactiontime="+80" swimtime="00:01:00.99" resultid="4225" heatid="5847" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="292" reactiontime="+71" swimtime="00:02:39.05" resultid="4226" heatid="5907" lane="2" entrytime="00:02:35.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                    <SPLIT distance="150" swimtime="00:01:59.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="308" reactiontime="+54" swimtime="00:01:11.50" resultid="4227" heatid="5961" lane="0" entrytime="00:01:11.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="401" swimtime="00:04:47.82" resultid="4228" heatid="5983" lane="9" entrytime="00:04:48.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:44.51" />
                    <SPLIT distance="200" swimtime="00:02:21.24" />
                    <SPLIT distance="250" swimtime="00:02:58.70" />
                    <SPLIT distance="300" swimtime="00:03:36.04" />
                    <SPLIT distance="350" swimtime="00:04:13.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mieszko" lastname="Palmi-Kukiełko" birthdate="1993-09-15" gender="M" nation="POL" license="101713700006" swrid="4073437" athleteid="4161">
              <RESULTS>
                <RESULT eventid="1076" points="582" reactiontime="+72" swimtime="00:00:26.04" resultid="4162" heatid="5783" lane="8" entrytime="00:00:26.24" />
                <RESULT eventid="1178" points="560" reactiontime="+72" swimtime="00:02:12.95" resultid="4163" heatid="5820" lane="4" entrytime="00:02:09.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="100" swimtime="00:01:04.01" />
                    <SPLIT distance="150" swimtime="00:01:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="549" reactiontime="+74" swimtime="00:01:00.16" resultid="4164" heatid="5893" lane="6" entrytime="00:00:59.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="485" reactiontime="+75" swimtime="00:02:14.40" resultid="4165" heatid="5908" lane="5" entrytime="00:02:07.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="567" reactiontime="+74" swimtime="00:00:57.70" resultid="4166" heatid="5971" lane="6" entrytime="00:00:57.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="526" reactiontime="+73" swimtime="00:04:22.82" resultid="4167" heatid="5984" lane="8" entrytime="00:04:24.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="150" swimtime="00:01:36.34" />
                    <SPLIT distance="200" swimtime="00:02:10.21" />
                    <SPLIT distance="250" swimtime="00:02:43.90" />
                    <SPLIT distance="300" swimtime="00:03:18.33" />
                    <SPLIT distance="350" swimtime="00:03:51.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="527" reactiontime="+70" swimtime="00:01:41.21" resultid="4229" heatid="5914" lane="6" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.42" />
                    <SPLIT distance="100" swimtime="00:00:49.70" />
                    <SPLIT distance="150" swimtime="00:01:16.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4206" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4168" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4222" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="4161" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" points="531" reactiontime="+65" swimtime="00:01:51.67" resultid="4231" heatid="5989" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                    <SPLIT distance="150" swimtime="00:01:25.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4161" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="4217" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="4206" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4168" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1442" points="347" reactiontime="+72" swimtime="00:01:56.40" resultid="4230" heatid="5913" lane="2" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:00:57.02" />
                    <SPLIT distance="150" swimtime="00:01:26.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4174" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4217" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="4187" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4180" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="3325" name="TJ Slovan Karlovy Vary" />
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="4357" name="KS AZS AWF Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Szczutkowski" birthdate="1998-04-11" gender="M" nation="POL" license="100201700161" swrid="4779469" athleteid="4373">
              <RESULTS>
                <RESULT eventid="1110" points="581" reactiontime="+68" swimtime="00:01:06.29" resultid="4374" heatid="5796" lane="6" entrytime="00:01:05.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="638" reactiontime="+67" swimtime="00:00:29.33" resultid="4375" heatid="5866" lane="1" />
                <RESULT eventid="1469" points="597" reactiontime="+64" swimtime="00:00:23.94" resultid="4376" heatid="5940" lane="2" entrytime="00:00:23.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Zawiliński" birthdate="2000-01-01" gender="M" nation="POL" swrid="4910761" athleteid="3637">
              <RESULTS>
                <RESULT eventid="1076" points="498" reactiontime="+70" swimtime="00:00:27.43" resultid="3639" heatid="5781" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1469" points="469" swimtime="00:00:25.94" resultid="3640" heatid="5938" lane="7" entrytime="00:00:25.50" />
                <RESULT eventid="1265" points="489" reactiontime="+69" swimtime="00:00:57.04" resultid="3641" heatid="5856" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Pinkosz" birthdate="1998-04-26" gender="M" nation="POL" license="100201700138" swrid="4368915" athleteid="4365">
              <RESULTS>
                <RESULT eventid="1076" points="522" reactiontime="+58" swimtime="00:00:27.00" resultid="4366" heatid="5783" lane="2" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="1212" points="519" reactiontime="+61" swimtime="00:02:03.63" resultid="4367" heatid="5835" lane="4" entrytime="00:01:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="100" swimtime="00:00:57.79" />
                    <SPLIT distance="150" swimtime="00:01:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="606" reactiontime="+59" swimtime="00:00:53.08" resultid="4368" heatid="5858" lane="4" entrytime="00:00:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="324" reactiontime="+66" swimtime="00:02:37.50" resultid="4369" heatid="5900" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:01:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="482" reactiontime="+59" swimtime="00:01:00.93" resultid="4371" heatid="5971" lane="8" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4372" heatid="5984" lane="5" entrytime="00:04:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" swrid="4236079" athleteid="4358">
              <RESULTS>
                <RESULT eventid="1059" points="549" reactiontime="+72" swimtime="00:00:29.77" resultid="4359" heatid="5771" lane="3" entrytime="00:00:28.87" entrycourse="SCM" />
                <RESULT eventid="1161" points="534" reactiontime="+67" swimtime="00:02:30.16" resultid="4360" heatid="5814" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="553" reactiontime="+71" swimtime="00:01:01.21" resultid="4361" heatid="5844" lane="6" entrytime="00:01:00.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="560" reactiontime="+70" swimtime="00:01:08.55" resultid="4362" heatid="5881" lane="5" entrytime="00:01:08.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="549" reactiontime="+66" swimtime="00:00:27.99" resultid="4363" heatid="5922" lane="1" entrytime="00:00:27.34" entrycourse="SCM" />
                <RESULT eventid="1588" points="522" reactiontime="+67" swimtime="00:04:50.36" resultid="4364" heatid="5975" lane="5" entrytime="00:04:57.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:43.30" />
                    <SPLIT distance="200" swimtime="00:02:20.75" />
                    <SPLIT distance="250" swimtime="00:02:58.35" />
                    <SPLIT distance="300" swimtime="00:03:36.52" />
                    <SPLIT distance="350" swimtime="00:04:14.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jędrzej" lastname="Kuczma" birthdate="1998-05-04" gender="M" nation="POL" license="100201700170" swrid="4418715" athleteid="4377">
              <RESULTS>
                <RESULT eventid="1212" points="559" reactiontime="+69" swimtime="00:02:00.60" resultid="4378" heatid="5827" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="100" swimtime="00:00:57.77" />
                    <SPLIT distance="150" swimtime="00:01:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="515" swimtime="00:00:56.04" resultid="4379" heatid="5846" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="575" reactiontime="+71" swimtime="00:04:15.10" resultid="4380" heatid="5977" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                    <SPLIT distance="100" swimtime="00:00:58.39" />
                    <SPLIT distance="150" swimtime="00:01:30.41" />
                    <SPLIT distance="200" swimtime="00:02:03.33" />
                    <SPLIT distance="250" swimtime="00:02:35.71" />
                    <SPLIT distance="300" swimtime="00:03:09.01" />
                    <SPLIT distance="350" swimtime="00:03:42.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="4242" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="4262">
              <RESULTS>
                <RESULT eventid="1110" points="174" swimtime="00:01:38.97" resultid="4263" heatid="5791" lane="2" entrytime="00:01:37.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="87" swimtime="00:03:43.46" resultid="4264" heatid="5829" lane="2" entrytime="00:03:26.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:44.45" />
                    <SPLIT distance="150" swimtime="00:02:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="204" reactiontime="+76" swimtime="00:00:42.85" resultid="4265" heatid="5868" lane="5" entrytime="00:00:42.03" entrycourse="SCM" />
                <RESULT eventid="1333" points="97" swimtime="00:01:47.11" resultid="4266" heatid="5884" lane="7" entrytime="00:01:43.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="158" reactiontime="+73" swimtime="00:00:37.22" resultid="4267" heatid="5927" lane="1" entrytime="00:00:38.51" entrycourse="SCM" />
                <RESULT eventid="1537" points="50" reactiontime="+79" swimtime="00:02:10.47" resultid="4268" heatid="5957" lane="4" entrytime="00:02:04.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Safrończyk" birthdate="1988-05-30" gender="M" nation="POL" license="510414700001" swrid="4072743" athleteid="4269">
              <RESULTS>
                <RESULT eventid="1110" status="DNS" swimtime="00:00:00.00" resultid="4270" heatid="5796" lane="4" entrytime="00:01:01.76" entrycourse="SCM" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="4271" heatid="5874" lane="5" entrytime="00:00:28.53" entrycourse="SCM" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4272" heatid="5893" lane="5" entrytime="00:00:57.50" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4273" heatid="5940" lane="5" entrytime="00:00:23.20" />
                <RESULT eventid="1503" status="DNS" swimtime="00:00:00.00" resultid="4274" heatid="5950" lane="5" entrytime="00:02:24.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="510414600003" swrid="5240601" athleteid="4255">
              <RESULTS>
                <RESULT eventid="1093" points="411" reactiontime="+73" swimtime="00:01:23.84" resultid="4256" heatid="5788" lane="1" entrytime="00:01:26.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="317" reactiontime="+79" swimtime="00:02:41.79" resultid="4257" heatid="5822" lane="4" entrytime="00:03:26.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="406" reactiontime="+76" swimtime="00:00:38.54" resultid="4258" heatid="5864" lane="1" entrytime="00:00:38.18" entrycourse="SCM" />
                <RESULT eventid="1316" points="314" reactiontime="+68" swimtime="00:01:23.09" resultid="4259" heatid="5879" lane="8" entrytime="00:01:24.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="383" reactiontime="+85" swimtime="00:03:05.27" resultid="4260" heatid="5944" lane="3" entrytime="00:03:05.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:01:29.52" />
                    <SPLIT distance="150" swimtime="00:02:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="330" reactiontime="+83" swimtime="00:05:38.29" resultid="4261" heatid="5974" lane="5" entrytime="00:05:49.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                    <SPLIT distance="200" swimtime="00:02:49.61" />
                    <SPLIT distance="250" swimtime="00:03:31.98" />
                    <SPLIT distance="300" swimtime="00:04:15.01" />
                    <SPLIT distance="350" swimtime="00:04:57.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" athleteid="3133">
              <RESULTS>
                <RESULT eventid="1144" points="97" reactiontime="+81" swimtime="00:00:48.22" resultid="3134" heatid="5805" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="1212" points="87" reactiontime="+85" swimtime="00:03:44.21" resultid="3135" heatid="5827" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="100" swimtime="00:01:43.53" />
                    <SPLIT distance="150" swimtime="00:02:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="97" reactiontime="+90" swimtime="00:01:37.76" resultid="3136" heatid="5846" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="87" reactiontime="+98" swimtime="00:03:57.94" resultid="3137" heatid="5904" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.53" />
                    <SPLIT distance="100" swimtime="00:01:56.64" />
                    <SPLIT distance="150" swimtime="00:02:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="127" reactiontime="+82" swimtime="00:00:40.07" resultid="3138" heatid="5926" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1537" points="85" reactiontime="+89" swimtime="00:01:49.84" resultid="3139" heatid="5957" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="4243">
              <RESULTS>
                <RESULT eventid="1076" points="142" swimtime="00:00:41.62" resultid="4244" heatid="5774" lane="2" entrytime="00:00:41.85" />
                <RESULT eventid="1367" points="107" reactiontime="+102" swimtime="00:03:47.90" resultid="4245" heatid="5897" lane="6" entrytime="00:04:00.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:39.16" />
                    <SPLIT distance="150" swimtime="00:02:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="192" reactiontime="+114" swimtime="00:03:27.95" resultid="4246" heatid="5945" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="126" swimtime="00:01:35.30" resultid="4247" heatid="5965" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Matusiewicz" birthdate="1998-04-12" gender="M" nation="POL" license="110414700069" swrid="5058424" athleteid="4248">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="4249" heatid="5773" lane="4" entrytime="00:00:47.72" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="4250" heatid="5829" lane="1" entrytime="00:03:28.88" />
                <RESULT eventid="1265" status="DNS" swimtime="00:00:00.00" resultid="4251" heatid="5848" lane="2" entrytime="00:01:32.12" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="4252" heatid="5884" lane="9" entrytime="00:01:45.75" />
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4253" heatid="5926" lane="6" entrytime="00:00:40.30" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4254" heatid="5976" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Domeracki" birthdate="1982-02-27" gender="M" nation="POL" license="510414700038" athleteid="4275">
              <RESULTS>
                <RESULT eventid="1212" points="262" reactiontime="+99" swimtime="00:02:35.13" resultid="4276" heatid="5832" lane="3" entrytime="00:02:32.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="237" swimtime="00:01:12.54" resultid="4277" heatid="5852" lane="9" entrytime="00:01:09.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" status="DNS" swimtime="00:00:00.00" resultid="4278" heatid="5930" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="1605" status="DNS" swimtime="00:00:00.00" resultid="4279" heatid="5981" lane="4" entrytime="00:05:11.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1442" points="147" reactiontime="+86" swimtime="00:02:34.95" resultid="4280" heatid="5911" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:01.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3133" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="4262" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4243" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4275" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1646" status="DNS" swimtime="00:00:00.00" resultid="4281" heatid="5987" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3133" number="1" />
                    <RELAYPOSITION athleteid="4262" number="2" />
                    <RELAYPOSITION athleteid="4243" number="3" />
                    <RELAYPOSITION athleteid="4275" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="4545" name="MKS ,,Astoria&apos;&apos; Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Ciężki" birthdate="1994-09-30" gender="M" nation="POL" license="102202700137" swrid="4289450" athleteid="4560">
              <RESULTS>
                <RESULT eventid="1212" points="534" reactiontime="+80" swimtime="00:02:02.43" resultid="4561" heatid="5826" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="100" swimtime="00:00:57.08" />
                    <SPLIT distance="150" swimtime="00:01:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="512" reactiontime="+78" swimtime="00:00:56.15" resultid="4562" heatid="5857" lane="8" entrytime="00:00:56.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="518" reactiontime="+73" swimtime="00:00:25.09" resultid="4563" heatid="5923" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Krasicki" birthdate="1995-02-17" gender="M" nation="POL" license="102202700140" swrid="4169744" athleteid="4564">
              <RESULTS>
                <RESULT eventid="1265" points="522" swimtime="00:00:55.80" resultid="4565" heatid="5847" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="508" reactiontime="+75" swimtime="00:00:25.26" resultid="4566" heatid="5923" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wawrzyniec" lastname="Manczak" birthdate="1948-06-03" gender="M" nation="POL" license="102202700108" swrid="4186189" athleteid="4551">
              <RESULTS>
                <RESULT eventid="1144" points="127" reactiontime="+87" swimtime="00:00:44.20" resultid="4552" heatid="5803" lane="6" />
                <RESULT eventid="1265" points="111" reactiontime="+95" swimtime="00:01:33.45" resultid="4553" heatid="5846" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="159" swimtime="00:00:37.15" resultid="4554" heatid="5924" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="4546">
              <RESULTS>
                <RESULT eventid="1144" points="88" reactiontime="+84" swimtime="00:00:49.92" resultid="4547" heatid="5804" lane="6" entrytime="00:00:53.36" entrycourse="SCM" />
                <RESULT eventid="1299" points="156" reactiontime="+75" swimtime="00:00:46.85" resultid="4548" heatid="5867" lane="5" entrytime="00:00:48.74" entrycourse="SCM" />
                <RESULT eventid="1469" points="140" swimtime="00:00:38.78" resultid="4549" heatid="5927" lane="7" entrytime="00:00:38.04" entrycourse="SCM" />
                <RESULT eventid="1537" points="64" reactiontime="+91" swimtime="00:02:00.73" resultid="4550" heatid="5958" lane="0" entrytime="00:01:55.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Bakuniak" birthdate="1996-03-25" gender="F" nation="POL" license="102202600136" swrid="4169734" athleteid="4555">
              <RESULTS>
                <RESULT eventid="1195" points="524" reactiontime="+57" swimtime="00:02:16.97" resultid="4556" heatid="5822" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="476" reactiontime="+65" swimtime="00:01:04.32" resultid="4557" heatid="5843" lane="4" entrytime="00:01:04.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1384" points="475" reactiontime="+74" swimtime="00:02:32.35" resultid="4558" heatid="5901" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="150" swimtime="00:01:52.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1588" points="565" reactiontime="+66" swimtime="00:04:42.90" resultid="4559" heatid="5975" lane="4" entrytime="00:04:44.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="150" swimtime="00:01:42.11" />
                    <SPLIT distance="200" swimtime="00:02:18.14" />
                    <SPLIT distance="250" swimtime="00:02:53.98" />
                    <SPLIT distance="300" swimtime="00:03:30.83" />
                    <SPLIT distance="350" swimtime="00:04:08.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3923" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Bogusiak" birthdate="1982-01-01" gender="M" nation="POL" athleteid="3922">
              <RESULTS>
                <RESULT eventid="1265" points="198" reactiontime="+92" swimtime="00:01:17.04" resultid="3924" heatid="5849" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="177" reactiontime="+90" swimtime="00:00:35.88" resultid="3925" heatid="5928" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1605" points="147" reactiontime="+96" swimtime="00:06:41.57" resultid="3926" heatid="5979" lane="8" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:30.11" />
                    <SPLIT distance="200" swimtime="00:03:12.26" />
                    <SPLIT distance="250" swimtime="00:04:05.31" />
                    <SPLIT distance="300" swimtime="00:04:58.29" />
                    <SPLIT distance="350" swimtime="00:05:50.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="4851" name="UKP Unia Oświęcim">
          <ATHLETES>
            <ATHLETE firstname="Jolanta" lastname="Płatek" birthdate="1971-09-10" gender="F" nation="POL" license="501006600380" swrid="4992931" athleteid="4864">
              <RESULTS>
                <RESULT eventid="1127" points="302" reactiontime="+80" swimtime="00:00:38.15" resultid="4865" heatid="5800" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1384" points="257" reactiontime="+80" swimtime="00:03:06.93" resultid="4866" heatid="5902" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:19.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1520" points="265" reactiontime="+83" swimtime="00:01:25.42" resultid="4867" heatid="5953" lane="5" entrytime="00:01:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Lipniarska-Skubis" birthdate="1952-07-01" gender="F" nation="POL" license="501006600377" athleteid="4852">
              <RESULTS>
                <RESULT eventid="1093" points="86" swimtime="00:02:21.02" resultid="4853" heatid="5786" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="90" swimtime="00:01:03.71" resultid="4854" heatid="5861" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="1451" points="71" swimtime="00:00:55.25" resultid="4855" heatid="5917" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1486" points="90" swimtime="00:04:59.40" resultid="4856" heatid="5942" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.71" />
                    <SPLIT distance="100" swimtime="00:02:22.71" />
                    <SPLIT distance="150" swimtime="00:03:41.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ilona" lastname="Szkudlarz" birthdate="1966-05-03" gender="F" nation="POL" license="501006600383" swrid="4992932" athleteid="4857">
              <RESULTS>
                <RESULT eventid="1093" points="229" reactiontime="+82" swimtime="00:01:41.91" resultid="4858" heatid="5787" lane="8" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="193" reactiontime="+73" swimtime="00:00:44.26" resultid="4859" heatid="5799" lane="6" entrytime="00:00:45.50" />
                <RESULT eventid="1247" points="237" reactiontime="+84" swimtime="00:01:21.18" resultid="4860" heatid="5841" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="222" reactiontime="+88" swimtime="00:00:47.15" resultid="4861" heatid="5862" lane="6" entrytime="00:00:46.50" />
                <RESULT eventid="1451" points="274" reactiontime="+80" swimtime="00:00:35.29" resultid="4862" heatid="5918" lane="3" entrytime="00:00:36.50" />
                <RESULT eventid="1520" points="186" reactiontime="+81" swimtime="00:01:36.00" resultid="4863" heatid="5953" lane="1" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Dorywalski" birthdate="1961-03-16" gender="M" nation="POL" license="501006700378" swrid="4992929" athleteid="4868">
              <RESULTS>
                <RESULT eventid="1144" points="187" reactiontime="+70" swimtime="00:00:38.84" resultid="4869" heatid="5806" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1401" points="191" reactiontime="+72" swimtime="00:03:03.37" resultid="4870" heatid="5906" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                    <SPLIT distance="100" swimtime="00:01:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="199" reactiontime="+78" swimtime="00:01:22.74" resultid="4871" heatid="5959" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5365" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Klimaszyk" birthdate="1995-01-01" gender="M" nation="POL" athleteid="5364">
              <RESULTS>
                <RESULT eventid="1076" points="395" reactiontime="+64" swimtime="00:00:29.64" resultid="5366" heatid="5782" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1212" points="387" reactiontime="+65" swimtime="00:02:16.28" resultid="5367" heatid="5826" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:01:01.21" />
                    <SPLIT distance="150" swimtime="00:01:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="425" reactiontime="+65" swimtime="00:00:26.81" resultid="5368" heatid="5938" lane="3" entrytime="00:00:25.43" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" clubid="2769" name="AZS AWF Katowice">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Ślężyński" birthdate="1931-04-27" gender="M" nation="POL" license="100611700315" swrid="4992723" athleteid="2770">
              <RESULTS>
                <RESULT eventid="1110" points="26" reactiontime="+134" swimtime="00:03:05.63" resultid="2771" heatid="5789" lane="4" entrytime="00:02:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="19" reactiontime="+89" swimtime="00:06:08.90" resultid="2772" heatid="5828" lane="9" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.04" />
                    <SPLIT distance="100" swimtime="00:03:01.83" />
                    <SPLIT distance="150" swimtime="00:04:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="15" swimtime="00:02:59.59" resultid="2773" heatid="5847" lane="2" entrytime="00:02:29.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="29" reactiontime="+94" swimtime="00:01:22.10" resultid="2774" heatid="5866" lane="3" entrytime="00:01:08.57" />
                <RESULT eventid="1503" points="24" reactiontime="+94" swimtime="00:06:51.70" resultid="2775" heatid="5945" lane="4" entrytime="00:05:23.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.21" />
                    <SPLIT distance="100" swimtime="00:03:22.20" />
                    <SPLIT distance="150" swimtime="00:05:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej a przed sygnałem startu." eventid="1605" status="DSQ" swimtime="00:00:00.00" resultid="2776" heatid="5977" lane="2" entrytime="00:10:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:39.74" />
                    <SPLIT distance="100" swimtime="00:03:33.13" />
                    <SPLIT distance="150" swimtime="00:05:21.10" />
                    <SPLIT distance="200" swimtime="00:07:03.33" />
                    <SPLIT distance="250" swimtime="00:08:48.50" />
                    <SPLIT distance="300" swimtime="00:10:28.91" />
                    <SPLIT distance="350" swimtime="00:12:13.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5728" name="Rydułtowy">
          <ATHLETES>
            <ATHLETE firstname="Rudolf" lastname="Bugla" birthdate="1940-01-01" gender="M" nation="POL" athleteid="5735">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="5736" heatid="5772" lane="0" />
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="5737" heatid="5815" lane="3" />
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="5738" heatid="5882" lane="4" />
                <RESULT eventid="1401" status="DNS" swimtime="00:00:00.00" resultid="5739" heatid="5904" lane="7" />
                <RESULT eventid="1537" status="DNS" swimtime="00:00:00.00" resultid="5740" heatid="5957" lane="1" />
                <RESULT eventid="1571" status="DNS" swimtime="00:00:00.00" resultid="5741" heatid="5965" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-01-01" gender="M" nation="POL" athleteid="5727">
              <RESULTS>
                <RESULT eventid="1076" points="176" reactiontime="+72" swimtime="00:00:38.75" resultid="5729" heatid="5774" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1144" points="141" reactiontime="+90" swimtime="00:00:42.64" resultid="5730" heatid="5806" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1367" points="86" reactiontime="+84" swimtime="00:04:05.12" resultid="5731" heatid="5897" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:56.97" />
                    <SPLIT distance="150" swimtime="00:03:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="123" reactiontime="+103" swimtime="00:03:32.12" resultid="5732" heatid="5905" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.88" />
                    <SPLIT distance="100" swimtime="00:01:46.25" />
                    <SPLIT distance="150" swimtime="00:02:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1537" points="139" reactiontime="+95" swimtime="00:01:33.28" resultid="5733" heatid="5958" lane="3" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="89" swimtime="00:01:46.98" resultid="5734" heatid="5966" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Władysław" lastname="Szurek" birthdate="1940-01-01" gender="M" nation="POL" athleteid="5742">
              <RESULTS>
                <RESULT eventid="1144" points="8" reactiontime="+79" swimtime="00:01:48.66" resultid="5743" heatid="5803" lane="4" />
                <RESULT eventid="1212" points="17" swimtime="00:06:24.35" resultid="5744" heatid="5827" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.49" />
                    <SPLIT distance="100" swimtime="00:03:01.37" />
                    <SPLIT distance="150" swimtime="00:04:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="15" swimtime="00:03:01.74" resultid="5745" heatid="5846" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="8" reactiontime="+94" swimtime="00:08:47.45" resultid="5746" heatid="5904" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:50.62" />
                    <SPLIT distance="100" swimtime="00:04:07.28" />
                    <SPLIT distance="150" swimtime="00:06:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="17" reactiontime="+81" swimtime="00:01:18.01" resultid="5747" heatid="5924" lane="8" />
                <RESULT eventid="1537" points="7" reactiontime="+89" swimtime="00:04:04.52" resultid="5748" heatid="5957" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:51.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Irczyk" birthdate="1951-01-01" gender="M" nation="POL" athleteid="5749">
              <RESULTS>
                <RESULT eventid="1178" points="63" reactiontime="+132" swimtime="00:04:34.70" resultid="5750" heatid="5816" lane="8" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.91" />
                    <SPLIT distance="100" swimtime="00:02:30.30" />
                    <SPLIT distance="150" swimtime="00:03:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="79" reactiontime="+124" swimtime="00:03:50.88" resultid="5751" heatid="5828" lane="8" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.09" />
                    <SPLIT distance="100" swimtime="00:01:56.86" />
                    <SPLIT distance="150" swimtime="00:02:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="52" reactiontime="+127" swimtime="00:02:11.51" resultid="5752" heatid="5883" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1367" points="45" reactiontime="+106" swimtime="00:05:04.29" resultid="5753" heatid="5897" lane="7" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.48" />
                    <SPLIT distance="100" swimtime="00:02:28.98" />
                    <SPLIT distance="150" swimtime="00:03:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="93" reactiontime="+118" swimtime="00:04:24.98" resultid="5754" heatid="5946" lane="9" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.33" />
                    <SPLIT distance="100" swimtime="00:02:07.74" />
                    <SPLIT distance="150" swimtime="00:03:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="97" swimtime="00:07:41.37" resultid="5755" heatid="5978" lane="9" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.30" />
                    <SPLIT distance="100" swimtime="00:01:53.61" />
                    <SPLIT distance="150" swimtime="00:02:53.85" />
                    <SPLIT distance="200" swimtime="00:03:54.20" />
                    <SPLIT distance="250" swimtime="00:04:53.86" />
                    <SPLIT distance="300" swimtime="00:05:50.29" />
                    <SPLIT distance="350" swimtime="00:06:47.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5200" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Dańkowski" birthdate="2000-01-01" gender="M" nation="POL" athleteid="5199">
              <RESULTS>
                <RESULT eventid="1469" points="468" reactiontime="+66" swimtime="00:00:25.95" resultid="5201" heatid="5938" lane="9" entrytime="00:00:26.00" />
                <RESULT eventid="1605" points="446" reactiontime="+65" swimtime="00:04:37.76" resultid="5202" heatid="5983" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:06.37" />
                    <SPLIT distance="150" swimtime="00:01:41.44" />
                    <SPLIT distance="200" swimtime="00:02:16.75" />
                    <SPLIT distance="250" swimtime="00:02:51.81" />
                    <SPLIT distance="300" swimtime="00:03:27.31" />
                    <SPLIT distance="350" swimtime="00:04:03.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3480" name="niezrzeszony">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Rusinowicz" birthdate="1944-01-01" gender="M" nation="POL" athleteid="3479">
              <RESULTS>
                <RESULT eventid="1110" points="69" reactiontime="+124" swimtime="00:02:14.61" resultid="3481" heatid="5790" lane="0" entrytime="00:02:12.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="59" reactiontime="+133" swimtime="00:04:14.63" resultid="3482" heatid="5828" lane="1" entrytime="00:04:15.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.15" />
                    <SPLIT distance="100" swimtime="00:02:02.85" />
                    <SPLIT distance="150" swimtime="00:03:09.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="64" reactiontime="+117" swimtime="00:01:52.14" resultid="3483" heatid="5847" lane="5" entrytime="00:01:51.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1401" points="48" reactiontime="+74" swimtime="00:04:48.99" resultid="3484" heatid="5904" lane="6" entrytime="00:04:45.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.68" />
                    <SPLIT distance="100" swimtime="00:02:18.19" />
                    <SPLIT distance="150" swimtime="00:03:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="60" reactiontime="+121" swimtime="00:05:06.03" resultid="3485" heatid="5946" lane="0" entrytime="00:04:49.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.35" />
                    <SPLIT distance="100" swimtime="00:02:24.45" />
                    <SPLIT distance="150" swimtime="00:03:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="62" reactiontime="+154" swimtime="00:08:54.54" resultid="3486" heatid="5977" lane="3" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                    <SPLIT distance="100" swimtime="00:02:06.00" />
                    <SPLIT distance="150" swimtime="00:03:14.34" />
                    <SPLIT distance="200" swimtime="00:04:22.59" />
                    <SPLIT distance="250" swimtime="00:05:30.65" />
                    <SPLIT distance="300" swimtime="00:06:39.55" />
                    <SPLIT distance="350" swimtime="00:07:48.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Harenda" birthdate="1968-01-01" gender="M" nation="POL" athleteid="3487">
              <RESULTS>
                <RESULT eventid="1076" points="219" reactiontime="+83" swimtime="00:00:36.06" resultid="3488" heatid="5776" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1212" points="241" reactiontime="+90" swimtime="00:02:39.66" resultid="3489" heatid="5832" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:01:57.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="280" reactiontime="+87" swimtime="00:01:08.67" resultid="3490" heatid="5852" lane="3" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="3491" heatid="5888" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="1537" points="181" reactiontime="+88" swimtime="00:01:25.29" resultid="3492" heatid="5959" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1605" points="211" swimtime="00:05:56.24" resultid="3493" heatid="5980" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:02:02.26" />
                    <SPLIT distance="200" swimtime="00:02:48.57" />
                    <SPLIT distance="250" swimtime="00:03:35.11" />
                    <SPLIT distance="300" swimtime="00:04:22.29" />
                    <SPLIT distance="350" swimtime="00:05:10.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3647" name="niezrzeszona">
          <ATHLETES>
            <ATHLETE firstname="Angelika" lastname="Wróbel" birthdate="1997-01-01" gender="F" nation="POL" swrid="4373387" athleteid="3646">
              <RESULTS>
                <RESULT eventid="1195" points="537" reactiontime="+90" swimtime="00:02:15.83" resultid="3648" heatid="5825" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:40.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="581" swimtime="00:01:00.21" resultid="3649" heatid="5844" lane="7" entrytime="00:01:00.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="563" reactiontime="+82" swimtime="00:00:27.76" resultid="3650" heatid="5922" lane="8" entrytime="00:00:27.58" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="5268" name="Artamonov Team">
          <ATHLETES>
            <ATHLETE firstname="Borys" lastname="Kushch" birthdate="1989-06-15" gender="M" nation="UKR" athleteid="3108">
              <RESULTS>
                <RESULT eventid="1265" points="307" swimtime="00:01:06.59" resultid="3109" heatid="5853" lane="7" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="359" reactiontime="+76" swimtime="00:00:28.35" resultid="3110" heatid="5933" lane="6" entrytime="00:00:28.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artem" lastname="Panchenko" birthdate="1992-12-24" gender="M" nation="UKR" athleteid="3111">
              <RESULTS>
                <RESULT eventid="1110" points="537" reactiontime="+74" swimtime="00:01:08.06" resultid="3112" heatid="5796" lane="8" entrytime="00:01:08.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="555" reactiontime="+72" swimtime="00:00:30.72" resultid="3113" heatid="5874" lane="8" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1333" points="413" reactiontime="+73" swimtime="00:01:06.17" resultid="3114" heatid="5892" lane="0" entrytime="00:01:06.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1503" points="475" reactiontime="+77" swimtime="00:02:33.94" resultid="3115" heatid="5950" lane="8" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1571" points="382" reactiontime="+73" swimtime="00:01:05.82" resultid="3116" heatid="5969" lane="6" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05806" nation="POL" region="06" clubid="4234" name="IKS Druga Strona Sportu">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" license="505806600021" swrid="5484417" athleteid="4235">
              <RESULTS>
                <RESULT eventid="1059" points="39" swimtime="00:01:11.68" resultid="4236" heatid="5766" lane="5" />
                <RESULT eventid="1127" points="76" reactiontime="+64" swimtime="00:01:00.21" resultid="4237" heatid="5798" lane="4" entrytime="00:01:02.95" entrycourse="SCM" />
                <RESULT eventid="1247" points="76" swimtime="00:01:58.23" resultid="4238" heatid="5840" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="71" reactiontime="+124" swimtime="00:02:16.01" resultid="4239" heatid="5876" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1451" points="90" reactiontime="+116" swimtime="00:00:51.03" resultid="4240" heatid="5917" lane="1" entrytime="00:00:53.24" entrycourse="SCM" />
                <RESULT eventid="1520" points="73" reactiontime="+121" swimtime="00:02:11.28" resultid="4241" heatid="5951" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
